library ieee;
use ieee.std_logic_1164.all;

entity VN2CN_wire is
  port (
      VN_data_out : in std_logic_vector(12287 downto 0);
      VN_sign_out : in std_logic_vector(12287 downto 0);
      CN_data_in : out std_logic_vector(12287 downto 0);
      CN_sign_in : out std_logic_vector(12287 downto 0)
    
  ) ;
end VN2CN_wire ;

architecture arch of VN2CN_wire is
signal CN0_data_in : std_logic_vector(31 downto 0);
signal CN0_sign_in : std_logic_vector(31 downto 0);
signal CN1_data_in : std_logic_vector(31 downto 0);
signal CN1_sign_in : std_logic_vector(31 downto 0);
signal CN2_data_in : std_logic_vector(31 downto 0);
signal CN2_sign_in : std_logic_vector(31 downto 0);
signal CN3_data_in : std_logic_vector(31 downto 0);
signal CN3_sign_in : std_logic_vector(31 downto 0);
signal CN4_data_in : std_logic_vector(31 downto 0);
signal CN4_sign_in : std_logic_vector(31 downto 0);
signal CN5_data_in : std_logic_vector(31 downto 0);
signal CN5_sign_in : std_logic_vector(31 downto 0);
signal CN6_data_in : std_logic_vector(31 downto 0);
signal CN6_sign_in : std_logic_vector(31 downto 0);
signal CN7_data_in : std_logic_vector(31 downto 0);
signal CN7_sign_in : std_logic_vector(31 downto 0);
signal CN8_data_in : std_logic_vector(31 downto 0);
signal CN8_sign_in : std_logic_vector(31 downto 0);
signal CN9_data_in : std_logic_vector(31 downto 0);
signal CN9_sign_in : std_logic_vector(31 downto 0);
signal CN10_data_in : std_logic_vector(31 downto 0);
signal CN10_sign_in : std_logic_vector(31 downto 0);
signal CN11_data_in : std_logic_vector(31 downto 0);
signal CN11_sign_in : std_logic_vector(31 downto 0);
signal CN12_data_in : std_logic_vector(31 downto 0);
signal CN12_sign_in : std_logic_vector(31 downto 0);
signal CN13_data_in : std_logic_vector(31 downto 0);
signal CN13_sign_in : std_logic_vector(31 downto 0);
signal CN14_data_in : std_logic_vector(31 downto 0);
signal CN14_sign_in : std_logic_vector(31 downto 0);
signal CN15_data_in : std_logic_vector(31 downto 0);
signal CN15_sign_in : std_logic_vector(31 downto 0);
signal CN16_data_in : std_logic_vector(31 downto 0);
signal CN16_sign_in : std_logic_vector(31 downto 0);
signal CN17_data_in : std_logic_vector(31 downto 0);
signal CN17_sign_in : std_logic_vector(31 downto 0);
signal CN18_data_in : std_logic_vector(31 downto 0);
signal CN18_sign_in : std_logic_vector(31 downto 0);
signal CN19_data_in : std_logic_vector(31 downto 0);
signal CN19_sign_in : std_logic_vector(31 downto 0);
signal CN20_data_in : std_logic_vector(31 downto 0);
signal CN20_sign_in : std_logic_vector(31 downto 0);
signal CN21_data_in : std_logic_vector(31 downto 0);
signal CN21_sign_in : std_logic_vector(31 downto 0);
signal CN22_data_in : std_logic_vector(31 downto 0);
signal CN22_sign_in : std_logic_vector(31 downto 0);
signal CN23_data_in : std_logic_vector(31 downto 0);
signal CN23_sign_in : std_logic_vector(31 downto 0);
signal CN24_data_in : std_logic_vector(31 downto 0);
signal CN24_sign_in : std_logic_vector(31 downto 0);
signal CN25_data_in : std_logic_vector(31 downto 0);
signal CN25_sign_in : std_logic_vector(31 downto 0);
signal CN26_data_in : std_logic_vector(31 downto 0);
signal CN26_sign_in : std_logic_vector(31 downto 0);
signal CN27_data_in : std_logic_vector(31 downto 0);
signal CN27_sign_in : std_logic_vector(31 downto 0);
signal CN28_data_in : std_logic_vector(31 downto 0);
signal CN28_sign_in : std_logic_vector(31 downto 0);
signal CN29_data_in : std_logic_vector(31 downto 0);
signal CN29_sign_in : std_logic_vector(31 downto 0);
signal CN30_data_in : std_logic_vector(31 downto 0);
signal CN30_sign_in : std_logic_vector(31 downto 0);
signal CN31_data_in : std_logic_vector(31 downto 0);
signal CN31_sign_in : std_logic_vector(31 downto 0);
signal CN32_data_in : std_logic_vector(31 downto 0);
signal CN32_sign_in : std_logic_vector(31 downto 0);
signal CN33_data_in : std_logic_vector(31 downto 0);
signal CN33_sign_in : std_logic_vector(31 downto 0);
signal CN34_data_in : std_logic_vector(31 downto 0);
signal CN34_sign_in : std_logic_vector(31 downto 0);
signal CN35_data_in : std_logic_vector(31 downto 0);
signal CN35_sign_in : std_logic_vector(31 downto 0);
signal CN36_data_in : std_logic_vector(31 downto 0);
signal CN36_sign_in : std_logic_vector(31 downto 0);
signal CN37_data_in : std_logic_vector(31 downto 0);
signal CN37_sign_in : std_logic_vector(31 downto 0);
signal CN38_data_in : std_logic_vector(31 downto 0);
signal CN38_sign_in : std_logic_vector(31 downto 0);
signal CN39_data_in : std_logic_vector(31 downto 0);
signal CN39_sign_in : std_logic_vector(31 downto 0);
signal CN40_data_in : std_logic_vector(31 downto 0);
signal CN40_sign_in : std_logic_vector(31 downto 0);
signal CN41_data_in : std_logic_vector(31 downto 0);
signal CN41_sign_in : std_logic_vector(31 downto 0);
signal CN42_data_in : std_logic_vector(31 downto 0);
signal CN42_sign_in : std_logic_vector(31 downto 0);
signal CN43_data_in : std_logic_vector(31 downto 0);
signal CN43_sign_in : std_logic_vector(31 downto 0);
signal CN44_data_in : std_logic_vector(31 downto 0);
signal CN44_sign_in : std_logic_vector(31 downto 0);
signal CN45_data_in : std_logic_vector(31 downto 0);
signal CN45_sign_in : std_logic_vector(31 downto 0);
signal CN46_data_in : std_logic_vector(31 downto 0);
signal CN46_sign_in : std_logic_vector(31 downto 0);
signal CN47_data_in : std_logic_vector(31 downto 0);
signal CN47_sign_in : std_logic_vector(31 downto 0);
signal CN48_data_in : std_logic_vector(31 downto 0);
signal CN48_sign_in : std_logic_vector(31 downto 0);
signal CN49_data_in : std_logic_vector(31 downto 0);
signal CN49_sign_in : std_logic_vector(31 downto 0);
signal CN50_data_in : std_logic_vector(31 downto 0);
signal CN50_sign_in : std_logic_vector(31 downto 0);
signal CN51_data_in : std_logic_vector(31 downto 0);
signal CN51_sign_in : std_logic_vector(31 downto 0);
signal CN52_data_in : std_logic_vector(31 downto 0);
signal CN52_sign_in : std_logic_vector(31 downto 0);
signal CN53_data_in : std_logic_vector(31 downto 0);
signal CN53_sign_in : std_logic_vector(31 downto 0);
signal CN54_data_in : std_logic_vector(31 downto 0);
signal CN54_sign_in : std_logic_vector(31 downto 0);
signal CN55_data_in : std_logic_vector(31 downto 0);
signal CN55_sign_in : std_logic_vector(31 downto 0);
signal CN56_data_in : std_logic_vector(31 downto 0);
signal CN56_sign_in : std_logic_vector(31 downto 0);
signal CN57_data_in : std_logic_vector(31 downto 0);
signal CN57_sign_in : std_logic_vector(31 downto 0);
signal CN58_data_in : std_logic_vector(31 downto 0);
signal CN58_sign_in : std_logic_vector(31 downto 0);
signal CN59_data_in : std_logic_vector(31 downto 0);
signal CN59_sign_in : std_logic_vector(31 downto 0);
signal CN60_data_in : std_logic_vector(31 downto 0);
signal CN60_sign_in : std_logic_vector(31 downto 0);
signal CN61_data_in : std_logic_vector(31 downto 0);
signal CN61_sign_in : std_logic_vector(31 downto 0);
signal CN62_data_in : std_logic_vector(31 downto 0);
signal CN62_sign_in : std_logic_vector(31 downto 0);
signal CN63_data_in : std_logic_vector(31 downto 0);
signal CN63_sign_in : std_logic_vector(31 downto 0);
signal CN64_data_in : std_logic_vector(31 downto 0);
signal CN64_sign_in : std_logic_vector(31 downto 0);
signal CN65_data_in : std_logic_vector(31 downto 0);
signal CN65_sign_in : std_logic_vector(31 downto 0);
signal CN66_data_in : std_logic_vector(31 downto 0);
signal CN66_sign_in : std_logic_vector(31 downto 0);
signal CN67_data_in : std_logic_vector(31 downto 0);
signal CN67_sign_in : std_logic_vector(31 downto 0);
signal CN68_data_in : std_logic_vector(31 downto 0);
signal CN68_sign_in : std_logic_vector(31 downto 0);
signal CN69_data_in : std_logic_vector(31 downto 0);
signal CN69_sign_in : std_logic_vector(31 downto 0);
signal CN70_data_in : std_logic_vector(31 downto 0);
signal CN70_sign_in : std_logic_vector(31 downto 0);
signal CN71_data_in : std_logic_vector(31 downto 0);
signal CN71_sign_in : std_logic_vector(31 downto 0);
signal CN72_data_in : std_logic_vector(31 downto 0);
signal CN72_sign_in : std_logic_vector(31 downto 0);
signal CN73_data_in : std_logic_vector(31 downto 0);
signal CN73_sign_in : std_logic_vector(31 downto 0);
signal CN74_data_in : std_logic_vector(31 downto 0);
signal CN74_sign_in : std_logic_vector(31 downto 0);
signal CN75_data_in : std_logic_vector(31 downto 0);
signal CN75_sign_in : std_logic_vector(31 downto 0);
signal CN76_data_in : std_logic_vector(31 downto 0);
signal CN76_sign_in : std_logic_vector(31 downto 0);
signal CN77_data_in : std_logic_vector(31 downto 0);
signal CN77_sign_in : std_logic_vector(31 downto 0);
signal CN78_data_in : std_logic_vector(31 downto 0);
signal CN78_sign_in : std_logic_vector(31 downto 0);
signal CN79_data_in : std_logic_vector(31 downto 0);
signal CN79_sign_in : std_logic_vector(31 downto 0);
signal CN80_data_in : std_logic_vector(31 downto 0);
signal CN80_sign_in : std_logic_vector(31 downto 0);
signal CN81_data_in : std_logic_vector(31 downto 0);
signal CN81_sign_in : std_logic_vector(31 downto 0);
signal CN82_data_in : std_logic_vector(31 downto 0);
signal CN82_sign_in : std_logic_vector(31 downto 0);
signal CN83_data_in : std_logic_vector(31 downto 0);
signal CN83_sign_in : std_logic_vector(31 downto 0);
signal CN84_data_in : std_logic_vector(31 downto 0);
signal CN84_sign_in : std_logic_vector(31 downto 0);
signal CN85_data_in : std_logic_vector(31 downto 0);
signal CN85_sign_in : std_logic_vector(31 downto 0);
signal CN86_data_in : std_logic_vector(31 downto 0);
signal CN86_sign_in : std_logic_vector(31 downto 0);
signal CN87_data_in : std_logic_vector(31 downto 0);
signal CN87_sign_in : std_logic_vector(31 downto 0);
signal CN88_data_in : std_logic_vector(31 downto 0);
signal CN88_sign_in : std_logic_vector(31 downto 0);
signal CN89_data_in : std_logic_vector(31 downto 0);
signal CN89_sign_in : std_logic_vector(31 downto 0);
signal CN90_data_in : std_logic_vector(31 downto 0);
signal CN90_sign_in : std_logic_vector(31 downto 0);
signal CN91_data_in : std_logic_vector(31 downto 0);
signal CN91_sign_in : std_logic_vector(31 downto 0);
signal CN92_data_in : std_logic_vector(31 downto 0);
signal CN92_sign_in : std_logic_vector(31 downto 0);
signal CN93_data_in : std_logic_vector(31 downto 0);
signal CN93_sign_in : std_logic_vector(31 downto 0);
signal CN94_data_in : std_logic_vector(31 downto 0);
signal CN94_sign_in : std_logic_vector(31 downto 0);
signal CN95_data_in : std_logic_vector(31 downto 0);
signal CN95_sign_in : std_logic_vector(31 downto 0);
signal CN96_data_in : std_logic_vector(31 downto 0);
signal CN96_sign_in : std_logic_vector(31 downto 0);
signal CN97_data_in : std_logic_vector(31 downto 0);
signal CN97_sign_in : std_logic_vector(31 downto 0);
signal CN98_data_in : std_logic_vector(31 downto 0);
signal CN98_sign_in : std_logic_vector(31 downto 0);
signal CN99_data_in : std_logic_vector(31 downto 0);
signal CN99_sign_in : std_logic_vector(31 downto 0);
signal CN100_data_in : std_logic_vector(31 downto 0);
signal CN100_sign_in : std_logic_vector(31 downto 0);
signal CN101_data_in : std_logic_vector(31 downto 0);
signal CN101_sign_in : std_logic_vector(31 downto 0);
signal CN102_data_in : std_logic_vector(31 downto 0);
signal CN102_sign_in : std_logic_vector(31 downto 0);
signal CN103_data_in : std_logic_vector(31 downto 0);
signal CN103_sign_in : std_logic_vector(31 downto 0);
signal CN104_data_in : std_logic_vector(31 downto 0);
signal CN104_sign_in : std_logic_vector(31 downto 0);
signal CN105_data_in : std_logic_vector(31 downto 0);
signal CN105_sign_in : std_logic_vector(31 downto 0);
signal CN106_data_in : std_logic_vector(31 downto 0);
signal CN106_sign_in : std_logic_vector(31 downto 0);
signal CN107_data_in : std_logic_vector(31 downto 0);
signal CN107_sign_in : std_logic_vector(31 downto 0);
signal CN108_data_in : std_logic_vector(31 downto 0);
signal CN108_sign_in : std_logic_vector(31 downto 0);
signal CN109_data_in : std_logic_vector(31 downto 0);
signal CN109_sign_in : std_logic_vector(31 downto 0);
signal CN110_data_in : std_logic_vector(31 downto 0);
signal CN110_sign_in : std_logic_vector(31 downto 0);
signal CN111_data_in : std_logic_vector(31 downto 0);
signal CN111_sign_in : std_logic_vector(31 downto 0);
signal CN112_data_in : std_logic_vector(31 downto 0);
signal CN112_sign_in : std_logic_vector(31 downto 0);
signal CN113_data_in : std_logic_vector(31 downto 0);
signal CN113_sign_in : std_logic_vector(31 downto 0);
signal CN114_data_in : std_logic_vector(31 downto 0);
signal CN114_sign_in : std_logic_vector(31 downto 0);
signal CN115_data_in : std_logic_vector(31 downto 0);
signal CN115_sign_in : std_logic_vector(31 downto 0);
signal CN116_data_in : std_logic_vector(31 downto 0);
signal CN116_sign_in : std_logic_vector(31 downto 0);
signal CN117_data_in : std_logic_vector(31 downto 0);
signal CN117_sign_in : std_logic_vector(31 downto 0);
signal CN118_data_in : std_logic_vector(31 downto 0);
signal CN118_sign_in : std_logic_vector(31 downto 0);
signal CN119_data_in : std_logic_vector(31 downto 0);
signal CN119_sign_in : std_logic_vector(31 downto 0);
signal CN120_data_in : std_logic_vector(31 downto 0);
signal CN120_sign_in : std_logic_vector(31 downto 0);
signal CN121_data_in : std_logic_vector(31 downto 0);
signal CN121_sign_in : std_logic_vector(31 downto 0);
signal CN122_data_in : std_logic_vector(31 downto 0);
signal CN122_sign_in : std_logic_vector(31 downto 0);
signal CN123_data_in : std_logic_vector(31 downto 0);
signal CN123_sign_in : std_logic_vector(31 downto 0);
signal CN124_data_in : std_logic_vector(31 downto 0);
signal CN124_sign_in : std_logic_vector(31 downto 0);
signal CN125_data_in : std_logic_vector(31 downto 0);
signal CN125_sign_in : std_logic_vector(31 downto 0);
signal CN126_data_in : std_logic_vector(31 downto 0);
signal CN126_sign_in : std_logic_vector(31 downto 0);
signal CN127_data_in : std_logic_vector(31 downto 0);
signal CN127_sign_in : std_logic_vector(31 downto 0);
signal CN128_data_in : std_logic_vector(31 downto 0);
signal CN128_sign_in : std_logic_vector(31 downto 0);
signal CN129_data_in : std_logic_vector(31 downto 0);
signal CN129_sign_in : std_logic_vector(31 downto 0);
signal CN130_data_in : std_logic_vector(31 downto 0);
signal CN130_sign_in : std_logic_vector(31 downto 0);
signal CN131_data_in : std_logic_vector(31 downto 0);
signal CN131_sign_in : std_logic_vector(31 downto 0);
signal CN132_data_in : std_logic_vector(31 downto 0);
signal CN132_sign_in : std_logic_vector(31 downto 0);
signal CN133_data_in : std_logic_vector(31 downto 0);
signal CN133_sign_in : std_logic_vector(31 downto 0);
signal CN134_data_in : std_logic_vector(31 downto 0);
signal CN134_sign_in : std_logic_vector(31 downto 0);
signal CN135_data_in : std_logic_vector(31 downto 0);
signal CN135_sign_in : std_logic_vector(31 downto 0);
signal CN136_data_in : std_logic_vector(31 downto 0);
signal CN136_sign_in : std_logic_vector(31 downto 0);
signal CN137_data_in : std_logic_vector(31 downto 0);
signal CN137_sign_in : std_logic_vector(31 downto 0);
signal CN138_data_in : std_logic_vector(31 downto 0);
signal CN138_sign_in : std_logic_vector(31 downto 0);
signal CN139_data_in : std_logic_vector(31 downto 0);
signal CN139_sign_in : std_logic_vector(31 downto 0);
signal CN140_data_in : std_logic_vector(31 downto 0);
signal CN140_sign_in : std_logic_vector(31 downto 0);
signal CN141_data_in : std_logic_vector(31 downto 0);
signal CN141_sign_in : std_logic_vector(31 downto 0);
signal CN142_data_in : std_logic_vector(31 downto 0);
signal CN142_sign_in : std_logic_vector(31 downto 0);
signal CN143_data_in : std_logic_vector(31 downto 0);
signal CN143_sign_in : std_logic_vector(31 downto 0);
signal CN144_data_in : std_logic_vector(31 downto 0);
signal CN144_sign_in : std_logic_vector(31 downto 0);
signal CN145_data_in : std_logic_vector(31 downto 0);
signal CN145_sign_in : std_logic_vector(31 downto 0);
signal CN146_data_in : std_logic_vector(31 downto 0);
signal CN146_sign_in : std_logic_vector(31 downto 0);
signal CN147_data_in : std_logic_vector(31 downto 0);
signal CN147_sign_in : std_logic_vector(31 downto 0);
signal CN148_data_in : std_logic_vector(31 downto 0);
signal CN148_sign_in : std_logic_vector(31 downto 0);
signal CN149_data_in : std_logic_vector(31 downto 0);
signal CN149_sign_in : std_logic_vector(31 downto 0);
signal CN150_data_in : std_logic_vector(31 downto 0);
signal CN150_sign_in : std_logic_vector(31 downto 0);
signal CN151_data_in : std_logic_vector(31 downto 0);
signal CN151_sign_in : std_logic_vector(31 downto 0);
signal CN152_data_in : std_logic_vector(31 downto 0);
signal CN152_sign_in : std_logic_vector(31 downto 0);
signal CN153_data_in : std_logic_vector(31 downto 0);
signal CN153_sign_in : std_logic_vector(31 downto 0);
signal CN154_data_in : std_logic_vector(31 downto 0);
signal CN154_sign_in : std_logic_vector(31 downto 0);
signal CN155_data_in : std_logic_vector(31 downto 0);
signal CN155_sign_in : std_logic_vector(31 downto 0);
signal CN156_data_in : std_logic_vector(31 downto 0);
signal CN156_sign_in : std_logic_vector(31 downto 0);
signal CN157_data_in : std_logic_vector(31 downto 0);
signal CN157_sign_in : std_logic_vector(31 downto 0);
signal CN158_data_in : std_logic_vector(31 downto 0);
signal CN158_sign_in : std_logic_vector(31 downto 0);
signal CN159_data_in : std_logic_vector(31 downto 0);
signal CN159_sign_in : std_logic_vector(31 downto 0);
signal CN160_data_in : std_logic_vector(31 downto 0);
signal CN160_sign_in : std_logic_vector(31 downto 0);
signal CN161_data_in : std_logic_vector(31 downto 0);
signal CN161_sign_in : std_logic_vector(31 downto 0);
signal CN162_data_in : std_logic_vector(31 downto 0);
signal CN162_sign_in : std_logic_vector(31 downto 0);
signal CN163_data_in : std_logic_vector(31 downto 0);
signal CN163_sign_in : std_logic_vector(31 downto 0);
signal CN164_data_in : std_logic_vector(31 downto 0);
signal CN164_sign_in : std_logic_vector(31 downto 0);
signal CN165_data_in : std_logic_vector(31 downto 0);
signal CN165_sign_in : std_logic_vector(31 downto 0);
signal CN166_data_in : std_logic_vector(31 downto 0);
signal CN166_sign_in : std_logic_vector(31 downto 0);
signal CN167_data_in : std_logic_vector(31 downto 0);
signal CN167_sign_in : std_logic_vector(31 downto 0);
signal CN168_data_in : std_logic_vector(31 downto 0);
signal CN168_sign_in : std_logic_vector(31 downto 0);
signal CN169_data_in : std_logic_vector(31 downto 0);
signal CN169_sign_in : std_logic_vector(31 downto 0);
signal CN170_data_in : std_logic_vector(31 downto 0);
signal CN170_sign_in : std_logic_vector(31 downto 0);
signal CN171_data_in : std_logic_vector(31 downto 0);
signal CN171_sign_in : std_logic_vector(31 downto 0);
signal CN172_data_in : std_logic_vector(31 downto 0);
signal CN172_sign_in : std_logic_vector(31 downto 0);
signal CN173_data_in : std_logic_vector(31 downto 0);
signal CN173_sign_in : std_logic_vector(31 downto 0);
signal CN174_data_in : std_logic_vector(31 downto 0);
signal CN174_sign_in : std_logic_vector(31 downto 0);
signal CN175_data_in : std_logic_vector(31 downto 0);
signal CN175_sign_in : std_logic_vector(31 downto 0);
signal CN176_data_in : std_logic_vector(31 downto 0);
signal CN176_sign_in : std_logic_vector(31 downto 0);
signal CN177_data_in : std_logic_vector(31 downto 0);
signal CN177_sign_in : std_logic_vector(31 downto 0);
signal CN178_data_in : std_logic_vector(31 downto 0);
signal CN178_sign_in : std_logic_vector(31 downto 0);
signal CN179_data_in : std_logic_vector(31 downto 0);
signal CN179_sign_in : std_logic_vector(31 downto 0);
signal CN180_data_in : std_logic_vector(31 downto 0);
signal CN180_sign_in : std_logic_vector(31 downto 0);
signal CN181_data_in : std_logic_vector(31 downto 0);
signal CN181_sign_in : std_logic_vector(31 downto 0);
signal CN182_data_in : std_logic_vector(31 downto 0);
signal CN182_sign_in : std_logic_vector(31 downto 0);
signal CN183_data_in : std_logic_vector(31 downto 0);
signal CN183_sign_in : std_logic_vector(31 downto 0);
signal CN184_data_in : std_logic_vector(31 downto 0);
signal CN184_sign_in : std_logic_vector(31 downto 0);
signal CN185_data_in : std_logic_vector(31 downto 0);
signal CN185_sign_in : std_logic_vector(31 downto 0);
signal CN186_data_in : std_logic_vector(31 downto 0);
signal CN186_sign_in : std_logic_vector(31 downto 0);
signal CN187_data_in : std_logic_vector(31 downto 0);
signal CN187_sign_in : std_logic_vector(31 downto 0);
signal CN188_data_in : std_logic_vector(31 downto 0);
signal CN188_sign_in : std_logic_vector(31 downto 0);
signal CN189_data_in : std_logic_vector(31 downto 0);
signal CN189_sign_in : std_logic_vector(31 downto 0);
signal CN190_data_in : std_logic_vector(31 downto 0);
signal CN190_sign_in : std_logic_vector(31 downto 0);
signal CN191_data_in : std_logic_vector(31 downto 0);
signal CN191_sign_in : std_logic_vector(31 downto 0);
signal CN192_data_in : std_logic_vector(31 downto 0);
signal CN192_sign_in : std_logic_vector(31 downto 0);
signal CN193_data_in : std_logic_vector(31 downto 0);
signal CN193_sign_in : std_logic_vector(31 downto 0);
signal CN194_data_in : std_logic_vector(31 downto 0);
signal CN194_sign_in : std_logic_vector(31 downto 0);
signal CN195_data_in : std_logic_vector(31 downto 0);
signal CN195_sign_in : std_logic_vector(31 downto 0);
signal CN196_data_in : std_logic_vector(31 downto 0);
signal CN196_sign_in : std_logic_vector(31 downto 0);
signal CN197_data_in : std_logic_vector(31 downto 0);
signal CN197_sign_in : std_logic_vector(31 downto 0);
signal CN198_data_in : std_logic_vector(31 downto 0);
signal CN198_sign_in : std_logic_vector(31 downto 0);
signal CN199_data_in : std_logic_vector(31 downto 0);
signal CN199_sign_in : std_logic_vector(31 downto 0);
signal CN200_data_in : std_logic_vector(31 downto 0);
signal CN200_sign_in : std_logic_vector(31 downto 0);
signal CN201_data_in : std_logic_vector(31 downto 0);
signal CN201_sign_in : std_logic_vector(31 downto 0);
signal CN202_data_in : std_logic_vector(31 downto 0);
signal CN202_sign_in : std_logic_vector(31 downto 0);
signal CN203_data_in : std_logic_vector(31 downto 0);
signal CN203_sign_in : std_logic_vector(31 downto 0);
signal CN204_data_in : std_logic_vector(31 downto 0);
signal CN204_sign_in : std_logic_vector(31 downto 0);
signal CN205_data_in : std_logic_vector(31 downto 0);
signal CN205_sign_in : std_logic_vector(31 downto 0);
signal CN206_data_in : std_logic_vector(31 downto 0);
signal CN206_sign_in : std_logic_vector(31 downto 0);
signal CN207_data_in : std_logic_vector(31 downto 0);
signal CN207_sign_in : std_logic_vector(31 downto 0);
signal CN208_data_in : std_logic_vector(31 downto 0);
signal CN208_sign_in : std_logic_vector(31 downto 0);
signal CN209_data_in : std_logic_vector(31 downto 0);
signal CN209_sign_in : std_logic_vector(31 downto 0);
signal CN210_data_in : std_logic_vector(31 downto 0);
signal CN210_sign_in : std_logic_vector(31 downto 0);
signal CN211_data_in : std_logic_vector(31 downto 0);
signal CN211_sign_in : std_logic_vector(31 downto 0);
signal CN212_data_in : std_logic_vector(31 downto 0);
signal CN212_sign_in : std_logic_vector(31 downto 0);
signal CN213_data_in : std_logic_vector(31 downto 0);
signal CN213_sign_in : std_logic_vector(31 downto 0);
signal CN214_data_in : std_logic_vector(31 downto 0);
signal CN214_sign_in : std_logic_vector(31 downto 0);
signal CN215_data_in : std_logic_vector(31 downto 0);
signal CN215_sign_in : std_logic_vector(31 downto 0);
signal CN216_data_in : std_logic_vector(31 downto 0);
signal CN216_sign_in : std_logic_vector(31 downto 0);
signal CN217_data_in : std_logic_vector(31 downto 0);
signal CN217_sign_in : std_logic_vector(31 downto 0);
signal CN218_data_in : std_logic_vector(31 downto 0);
signal CN218_sign_in : std_logic_vector(31 downto 0);
signal CN219_data_in : std_logic_vector(31 downto 0);
signal CN219_sign_in : std_logic_vector(31 downto 0);
signal CN220_data_in : std_logic_vector(31 downto 0);
signal CN220_sign_in : std_logic_vector(31 downto 0);
signal CN221_data_in : std_logic_vector(31 downto 0);
signal CN221_sign_in : std_logic_vector(31 downto 0);
signal CN222_data_in : std_logic_vector(31 downto 0);
signal CN222_sign_in : std_logic_vector(31 downto 0);
signal CN223_data_in : std_logic_vector(31 downto 0);
signal CN223_sign_in : std_logic_vector(31 downto 0);
signal CN224_data_in : std_logic_vector(31 downto 0);
signal CN224_sign_in : std_logic_vector(31 downto 0);
signal CN225_data_in : std_logic_vector(31 downto 0);
signal CN225_sign_in : std_logic_vector(31 downto 0);
signal CN226_data_in : std_logic_vector(31 downto 0);
signal CN226_sign_in : std_logic_vector(31 downto 0);
signal CN227_data_in : std_logic_vector(31 downto 0);
signal CN227_sign_in : std_logic_vector(31 downto 0);
signal CN228_data_in : std_logic_vector(31 downto 0);
signal CN228_sign_in : std_logic_vector(31 downto 0);
signal CN229_data_in : std_logic_vector(31 downto 0);
signal CN229_sign_in : std_logic_vector(31 downto 0);
signal CN230_data_in : std_logic_vector(31 downto 0);
signal CN230_sign_in : std_logic_vector(31 downto 0);
signal CN231_data_in : std_logic_vector(31 downto 0);
signal CN231_sign_in : std_logic_vector(31 downto 0);
signal CN232_data_in : std_logic_vector(31 downto 0);
signal CN232_sign_in : std_logic_vector(31 downto 0);
signal CN233_data_in : std_logic_vector(31 downto 0);
signal CN233_sign_in : std_logic_vector(31 downto 0);
signal CN234_data_in : std_logic_vector(31 downto 0);
signal CN234_sign_in : std_logic_vector(31 downto 0);
signal CN235_data_in : std_logic_vector(31 downto 0);
signal CN235_sign_in : std_logic_vector(31 downto 0);
signal CN236_data_in : std_logic_vector(31 downto 0);
signal CN236_sign_in : std_logic_vector(31 downto 0);
signal CN237_data_in : std_logic_vector(31 downto 0);
signal CN237_sign_in : std_logic_vector(31 downto 0);
signal CN238_data_in : std_logic_vector(31 downto 0);
signal CN238_sign_in : std_logic_vector(31 downto 0);
signal CN239_data_in : std_logic_vector(31 downto 0);
signal CN239_sign_in : std_logic_vector(31 downto 0);
signal CN240_data_in : std_logic_vector(31 downto 0);
signal CN240_sign_in : std_logic_vector(31 downto 0);
signal CN241_data_in : std_logic_vector(31 downto 0);
signal CN241_sign_in : std_logic_vector(31 downto 0);
signal CN242_data_in : std_logic_vector(31 downto 0);
signal CN242_sign_in : std_logic_vector(31 downto 0);
signal CN243_data_in : std_logic_vector(31 downto 0);
signal CN243_sign_in : std_logic_vector(31 downto 0);
signal CN244_data_in : std_logic_vector(31 downto 0);
signal CN244_sign_in : std_logic_vector(31 downto 0);
signal CN245_data_in : std_logic_vector(31 downto 0);
signal CN245_sign_in : std_logic_vector(31 downto 0);
signal CN246_data_in : std_logic_vector(31 downto 0);
signal CN246_sign_in : std_logic_vector(31 downto 0);
signal CN247_data_in : std_logic_vector(31 downto 0);
signal CN247_sign_in : std_logic_vector(31 downto 0);
signal CN248_data_in : std_logic_vector(31 downto 0);
signal CN248_sign_in : std_logic_vector(31 downto 0);
signal CN249_data_in : std_logic_vector(31 downto 0);
signal CN249_sign_in : std_logic_vector(31 downto 0);
signal CN250_data_in : std_logic_vector(31 downto 0);
signal CN250_sign_in : std_logic_vector(31 downto 0);
signal CN251_data_in : std_logic_vector(31 downto 0);
signal CN251_sign_in : std_logic_vector(31 downto 0);
signal CN252_data_in : std_logic_vector(31 downto 0);
signal CN252_sign_in : std_logic_vector(31 downto 0);
signal CN253_data_in : std_logic_vector(31 downto 0);
signal CN253_sign_in : std_logic_vector(31 downto 0);
signal CN254_data_in : std_logic_vector(31 downto 0);
signal CN254_sign_in : std_logic_vector(31 downto 0);
signal CN255_data_in : std_logic_vector(31 downto 0);
signal CN255_sign_in : std_logic_vector(31 downto 0);
signal CN256_data_in : std_logic_vector(31 downto 0);
signal CN256_sign_in : std_logic_vector(31 downto 0);
signal CN257_data_in : std_logic_vector(31 downto 0);
signal CN257_sign_in : std_logic_vector(31 downto 0);
signal CN258_data_in : std_logic_vector(31 downto 0);
signal CN258_sign_in : std_logic_vector(31 downto 0);
signal CN259_data_in : std_logic_vector(31 downto 0);
signal CN259_sign_in : std_logic_vector(31 downto 0);
signal CN260_data_in : std_logic_vector(31 downto 0);
signal CN260_sign_in : std_logic_vector(31 downto 0);
signal CN261_data_in : std_logic_vector(31 downto 0);
signal CN261_sign_in : std_logic_vector(31 downto 0);
signal CN262_data_in : std_logic_vector(31 downto 0);
signal CN262_sign_in : std_logic_vector(31 downto 0);
signal CN263_data_in : std_logic_vector(31 downto 0);
signal CN263_sign_in : std_logic_vector(31 downto 0);
signal CN264_data_in : std_logic_vector(31 downto 0);
signal CN264_sign_in : std_logic_vector(31 downto 0);
signal CN265_data_in : std_logic_vector(31 downto 0);
signal CN265_sign_in : std_logic_vector(31 downto 0);
signal CN266_data_in : std_logic_vector(31 downto 0);
signal CN266_sign_in : std_logic_vector(31 downto 0);
signal CN267_data_in : std_logic_vector(31 downto 0);
signal CN267_sign_in : std_logic_vector(31 downto 0);
signal CN268_data_in : std_logic_vector(31 downto 0);
signal CN268_sign_in : std_logic_vector(31 downto 0);
signal CN269_data_in : std_logic_vector(31 downto 0);
signal CN269_sign_in : std_logic_vector(31 downto 0);
signal CN270_data_in : std_logic_vector(31 downto 0);
signal CN270_sign_in : std_logic_vector(31 downto 0);
signal CN271_data_in : std_logic_vector(31 downto 0);
signal CN271_sign_in : std_logic_vector(31 downto 0);
signal CN272_data_in : std_logic_vector(31 downto 0);
signal CN272_sign_in : std_logic_vector(31 downto 0);
signal CN273_data_in : std_logic_vector(31 downto 0);
signal CN273_sign_in : std_logic_vector(31 downto 0);
signal CN274_data_in : std_logic_vector(31 downto 0);
signal CN274_sign_in : std_logic_vector(31 downto 0);
signal CN275_data_in : std_logic_vector(31 downto 0);
signal CN275_sign_in : std_logic_vector(31 downto 0);
signal CN276_data_in : std_logic_vector(31 downto 0);
signal CN276_sign_in : std_logic_vector(31 downto 0);
signal CN277_data_in : std_logic_vector(31 downto 0);
signal CN277_sign_in : std_logic_vector(31 downto 0);
signal CN278_data_in : std_logic_vector(31 downto 0);
signal CN278_sign_in : std_logic_vector(31 downto 0);
signal CN279_data_in : std_logic_vector(31 downto 0);
signal CN279_sign_in : std_logic_vector(31 downto 0);
signal CN280_data_in : std_logic_vector(31 downto 0);
signal CN280_sign_in : std_logic_vector(31 downto 0);
signal CN281_data_in : std_logic_vector(31 downto 0);
signal CN281_sign_in : std_logic_vector(31 downto 0);
signal CN282_data_in : std_logic_vector(31 downto 0);
signal CN282_sign_in : std_logic_vector(31 downto 0);
signal CN283_data_in : std_logic_vector(31 downto 0);
signal CN283_sign_in : std_logic_vector(31 downto 0);
signal CN284_data_in : std_logic_vector(31 downto 0);
signal CN284_sign_in : std_logic_vector(31 downto 0);
signal CN285_data_in : std_logic_vector(31 downto 0);
signal CN285_sign_in : std_logic_vector(31 downto 0);
signal CN286_data_in : std_logic_vector(31 downto 0);
signal CN286_sign_in : std_logic_vector(31 downto 0);
signal CN287_data_in : std_logic_vector(31 downto 0);
signal CN287_sign_in : std_logic_vector(31 downto 0);
signal CN288_data_in : std_logic_vector(31 downto 0);
signal CN288_sign_in : std_logic_vector(31 downto 0);
signal CN289_data_in : std_logic_vector(31 downto 0);
signal CN289_sign_in : std_logic_vector(31 downto 0);
signal CN290_data_in : std_logic_vector(31 downto 0);
signal CN290_sign_in : std_logic_vector(31 downto 0);
signal CN291_data_in : std_logic_vector(31 downto 0);
signal CN291_sign_in : std_logic_vector(31 downto 0);
signal CN292_data_in : std_logic_vector(31 downto 0);
signal CN292_sign_in : std_logic_vector(31 downto 0);
signal CN293_data_in : std_logic_vector(31 downto 0);
signal CN293_sign_in : std_logic_vector(31 downto 0);
signal CN294_data_in : std_logic_vector(31 downto 0);
signal CN294_sign_in : std_logic_vector(31 downto 0);
signal CN295_data_in : std_logic_vector(31 downto 0);
signal CN295_sign_in : std_logic_vector(31 downto 0);
signal CN296_data_in : std_logic_vector(31 downto 0);
signal CN296_sign_in : std_logic_vector(31 downto 0);
signal CN297_data_in : std_logic_vector(31 downto 0);
signal CN297_sign_in : std_logic_vector(31 downto 0);
signal CN298_data_in : std_logic_vector(31 downto 0);
signal CN298_sign_in : std_logic_vector(31 downto 0);
signal CN299_data_in : std_logic_vector(31 downto 0);
signal CN299_sign_in : std_logic_vector(31 downto 0);
signal CN300_data_in : std_logic_vector(31 downto 0);
signal CN300_sign_in : std_logic_vector(31 downto 0);
signal CN301_data_in : std_logic_vector(31 downto 0);
signal CN301_sign_in : std_logic_vector(31 downto 0);
signal CN302_data_in : std_logic_vector(31 downto 0);
signal CN302_sign_in : std_logic_vector(31 downto 0);
signal CN303_data_in : std_logic_vector(31 downto 0);
signal CN303_sign_in : std_logic_vector(31 downto 0);
signal CN304_data_in : std_logic_vector(31 downto 0);
signal CN304_sign_in : std_logic_vector(31 downto 0);
signal CN305_data_in : std_logic_vector(31 downto 0);
signal CN305_sign_in : std_logic_vector(31 downto 0);
signal CN306_data_in : std_logic_vector(31 downto 0);
signal CN306_sign_in : std_logic_vector(31 downto 0);
signal CN307_data_in : std_logic_vector(31 downto 0);
signal CN307_sign_in : std_logic_vector(31 downto 0);
signal CN308_data_in : std_logic_vector(31 downto 0);
signal CN308_sign_in : std_logic_vector(31 downto 0);
signal CN309_data_in : std_logic_vector(31 downto 0);
signal CN309_sign_in : std_logic_vector(31 downto 0);
signal CN310_data_in : std_logic_vector(31 downto 0);
signal CN310_sign_in : std_logic_vector(31 downto 0);
signal CN311_data_in : std_logic_vector(31 downto 0);
signal CN311_sign_in : std_logic_vector(31 downto 0);
signal CN312_data_in : std_logic_vector(31 downto 0);
signal CN312_sign_in : std_logic_vector(31 downto 0);
signal CN313_data_in : std_logic_vector(31 downto 0);
signal CN313_sign_in : std_logic_vector(31 downto 0);
signal CN314_data_in : std_logic_vector(31 downto 0);
signal CN314_sign_in : std_logic_vector(31 downto 0);
signal CN315_data_in : std_logic_vector(31 downto 0);
signal CN315_sign_in : std_logic_vector(31 downto 0);
signal CN316_data_in : std_logic_vector(31 downto 0);
signal CN316_sign_in : std_logic_vector(31 downto 0);
signal CN317_data_in : std_logic_vector(31 downto 0);
signal CN317_sign_in : std_logic_vector(31 downto 0);
signal CN318_data_in : std_logic_vector(31 downto 0);
signal CN318_sign_in : std_logic_vector(31 downto 0);
signal CN319_data_in : std_logic_vector(31 downto 0);
signal CN319_sign_in : std_logic_vector(31 downto 0);
signal CN320_data_in : std_logic_vector(31 downto 0);
signal CN320_sign_in : std_logic_vector(31 downto 0);
signal CN321_data_in : std_logic_vector(31 downto 0);
signal CN321_sign_in : std_logic_vector(31 downto 0);
signal CN322_data_in : std_logic_vector(31 downto 0);
signal CN322_sign_in : std_logic_vector(31 downto 0);
signal CN323_data_in : std_logic_vector(31 downto 0);
signal CN323_sign_in : std_logic_vector(31 downto 0);
signal CN324_data_in : std_logic_vector(31 downto 0);
signal CN324_sign_in : std_logic_vector(31 downto 0);
signal CN325_data_in : std_logic_vector(31 downto 0);
signal CN325_sign_in : std_logic_vector(31 downto 0);
signal CN326_data_in : std_logic_vector(31 downto 0);
signal CN326_sign_in : std_logic_vector(31 downto 0);
signal CN327_data_in : std_logic_vector(31 downto 0);
signal CN327_sign_in : std_logic_vector(31 downto 0);
signal CN328_data_in : std_logic_vector(31 downto 0);
signal CN328_sign_in : std_logic_vector(31 downto 0);
signal CN329_data_in : std_logic_vector(31 downto 0);
signal CN329_sign_in : std_logic_vector(31 downto 0);
signal CN330_data_in : std_logic_vector(31 downto 0);
signal CN330_sign_in : std_logic_vector(31 downto 0);
signal CN331_data_in : std_logic_vector(31 downto 0);
signal CN331_sign_in : std_logic_vector(31 downto 0);
signal CN332_data_in : std_logic_vector(31 downto 0);
signal CN332_sign_in : std_logic_vector(31 downto 0);
signal CN333_data_in : std_logic_vector(31 downto 0);
signal CN333_sign_in : std_logic_vector(31 downto 0);
signal CN334_data_in : std_logic_vector(31 downto 0);
signal CN334_sign_in : std_logic_vector(31 downto 0);
signal CN335_data_in : std_logic_vector(31 downto 0);
signal CN335_sign_in : std_logic_vector(31 downto 0);
signal CN336_data_in : std_logic_vector(31 downto 0);
signal CN336_sign_in : std_logic_vector(31 downto 0);
signal CN337_data_in : std_logic_vector(31 downto 0);
signal CN337_sign_in : std_logic_vector(31 downto 0);
signal CN338_data_in : std_logic_vector(31 downto 0);
signal CN338_sign_in : std_logic_vector(31 downto 0);
signal CN339_data_in : std_logic_vector(31 downto 0);
signal CN339_sign_in : std_logic_vector(31 downto 0);
signal CN340_data_in : std_logic_vector(31 downto 0);
signal CN340_sign_in : std_logic_vector(31 downto 0);
signal CN341_data_in : std_logic_vector(31 downto 0);
signal CN341_sign_in : std_logic_vector(31 downto 0);
signal CN342_data_in : std_logic_vector(31 downto 0);
signal CN342_sign_in : std_logic_vector(31 downto 0);
signal CN343_data_in : std_logic_vector(31 downto 0);
signal CN343_sign_in : std_logic_vector(31 downto 0);
signal CN344_data_in : std_logic_vector(31 downto 0);
signal CN344_sign_in : std_logic_vector(31 downto 0);
signal CN345_data_in : std_logic_vector(31 downto 0);
signal CN345_sign_in : std_logic_vector(31 downto 0);
signal CN346_data_in : std_logic_vector(31 downto 0);
signal CN346_sign_in : std_logic_vector(31 downto 0);
signal CN347_data_in : std_logic_vector(31 downto 0);
signal CN347_sign_in : std_logic_vector(31 downto 0);
signal CN348_data_in : std_logic_vector(31 downto 0);
signal CN348_sign_in : std_logic_vector(31 downto 0);
signal CN349_data_in : std_logic_vector(31 downto 0);
signal CN349_sign_in : std_logic_vector(31 downto 0);
signal CN350_data_in : std_logic_vector(31 downto 0);
signal CN350_sign_in : std_logic_vector(31 downto 0);
signal CN351_data_in : std_logic_vector(31 downto 0);
signal CN351_sign_in : std_logic_vector(31 downto 0);
signal CN352_data_in : std_logic_vector(31 downto 0);
signal CN352_sign_in : std_logic_vector(31 downto 0);
signal CN353_data_in : std_logic_vector(31 downto 0);
signal CN353_sign_in : std_logic_vector(31 downto 0);
signal CN354_data_in : std_logic_vector(31 downto 0);
signal CN354_sign_in : std_logic_vector(31 downto 0);
signal CN355_data_in : std_logic_vector(31 downto 0);
signal CN355_sign_in : std_logic_vector(31 downto 0);
signal CN356_data_in : std_logic_vector(31 downto 0);
signal CN356_sign_in : std_logic_vector(31 downto 0);
signal CN357_data_in : std_logic_vector(31 downto 0);
signal CN357_sign_in : std_logic_vector(31 downto 0);
signal CN358_data_in : std_logic_vector(31 downto 0);
signal CN358_sign_in : std_logic_vector(31 downto 0);
signal CN359_data_in : std_logic_vector(31 downto 0);
signal CN359_sign_in : std_logic_vector(31 downto 0);
signal CN360_data_in : std_logic_vector(31 downto 0);
signal CN360_sign_in : std_logic_vector(31 downto 0);
signal CN361_data_in : std_logic_vector(31 downto 0);
signal CN361_sign_in : std_logic_vector(31 downto 0);
signal CN362_data_in : std_logic_vector(31 downto 0);
signal CN362_sign_in : std_logic_vector(31 downto 0);
signal CN363_data_in : std_logic_vector(31 downto 0);
signal CN363_sign_in : std_logic_vector(31 downto 0);
signal CN364_data_in : std_logic_vector(31 downto 0);
signal CN364_sign_in : std_logic_vector(31 downto 0);
signal CN365_data_in : std_logic_vector(31 downto 0);
signal CN365_sign_in : std_logic_vector(31 downto 0);
signal CN366_data_in : std_logic_vector(31 downto 0);
signal CN366_sign_in : std_logic_vector(31 downto 0);
signal CN367_data_in : std_logic_vector(31 downto 0);
signal CN367_sign_in : std_logic_vector(31 downto 0);
signal CN368_data_in : std_logic_vector(31 downto 0);
signal CN368_sign_in : std_logic_vector(31 downto 0);
signal CN369_data_in : std_logic_vector(31 downto 0);
signal CN369_sign_in : std_logic_vector(31 downto 0);
signal CN370_data_in : std_logic_vector(31 downto 0);
signal CN370_sign_in : std_logic_vector(31 downto 0);
signal CN371_data_in : std_logic_vector(31 downto 0);
signal CN371_sign_in : std_logic_vector(31 downto 0);
signal CN372_data_in : std_logic_vector(31 downto 0);
signal CN372_sign_in : std_logic_vector(31 downto 0);
signal CN373_data_in : std_logic_vector(31 downto 0);
signal CN373_sign_in : std_logic_vector(31 downto 0);
signal CN374_data_in : std_logic_vector(31 downto 0);
signal CN374_sign_in : std_logic_vector(31 downto 0);
signal CN375_data_in : std_logic_vector(31 downto 0);
signal CN375_sign_in : std_logic_vector(31 downto 0);
signal CN376_data_in : std_logic_vector(31 downto 0);
signal CN376_sign_in : std_logic_vector(31 downto 0);
signal CN377_data_in : std_logic_vector(31 downto 0);
signal CN377_sign_in : std_logic_vector(31 downto 0);
signal CN378_data_in : std_logic_vector(31 downto 0);
signal CN378_sign_in : std_logic_vector(31 downto 0);
signal CN379_data_in : std_logic_vector(31 downto 0);
signal CN379_sign_in : std_logic_vector(31 downto 0);
signal CN380_data_in : std_logic_vector(31 downto 0);
signal CN380_sign_in : std_logic_vector(31 downto 0);
signal CN381_data_in : std_logic_vector(31 downto 0);
signal CN381_sign_in : std_logic_vector(31 downto 0);
signal CN382_data_in : std_logic_vector(31 downto 0);
signal CN382_sign_in : std_logic_vector(31 downto 0);
signal CN383_data_in : std_logic_vector(31 downto 0);
signal CN383_sign_in : std_logic_vector(31 downto 0);
signal VN0_data_out : std_logic_vector(5 downto 0);
signal VN0_sign_out : std_logic_vector(5 downto 0);
signal VN1_data_out : std_logic_vector(5 downto 0);
signal VN1_sign_out : std_logic_vector(5 downto 0);
signal VN2_data_out : std_logic_vector(5 downto 0);
signal VN2_sign_out : std_logic_vector(5 downto 0);
signal VN3_data_out : std_logic_vector(5 downto 0);
signal VN3_sign_out : std_logic_vector(5 downto 0);
signal VN4_data_out : std_logic_vector(5 downto 0);
signal VN4_sign_out : std_logic_vector(5 downto 0);
signal VN5_data_out : std_logic_vector(5 downto 0);
signal VN5_sign_out : std_logic_vector(5 downto 0);
signal VN6_data_out : std_logic_vector(5 downto 0);
signal VN6_sign_out : std_logic_vector(5 downto 0);
signal VN7_data_out : std_logic_vector(5 downto 0);
signal VN7_sign_out : std_logic_vector(5 downto 0);
signal VN8_data_out : std_logic_vector(5 downto 0);
signal VN8_sign_out : std_logic_vector(5 downto 0);
signal VN9_data_out : std_logic_vector(5 downto 0);
signal VN9_sign_out : std_logic_vector(5 downto 0);
signal VN10_data_out : std_logic_vector(5 downto 0);
signal VN10_sign_out : std_logic_vector(5 downto 0);
signal VN11_data_out : std_logic_vector(5 downto 0);
signal VN11_sign_out : std_logic_vector(5 downto 0);
signal VN12_data_out : std_logic_vector(5 downto 0);
signal VN12_sign_out : std_logic_vector(5 downto 0);
signal VN13_data_out : std_logic_vector(5 downto 0);
signal VN13_sign_out : std_logic_vector(5 downto 0);
signal VN14_data_out : std_logic_vector(5 downto 0);
signal VN14_sign_out : std_logic_vector(5 downto 0);
signal VN15_data_out : std_logic_vector(5 downto 0);
signal VN15_sign_out : std_logic_vector(5 downto 0);
signal VN16_data_out : std_logic_vector(5 downto 0);
signal VN16_sign_out : std_logic_vector(5 downto 0);
signal VN17_data_out : std_logic_vector(5 downto 0);
signal VN17_sign_out : std_logic_vector(5 downto 0);
signal VN18_data_out : std_logic_vector(5 downto 0);
signal VN18_sign_out : std_logic_vector(5 downto 0);
signal VN19_data_out : std_logic_vector(5 downto 0);
signal VN19_sign_out : std_logic_vector(5 downto 0);
signal VN20_data_out : std_logic_vector(5 downto 0);
signal VN20_sign_out : std_logic_vector(5 downto 0);
signal VN21_data_out : std_logic_vector(5 downto 0);
signal VN21_sign_out : std_logic_vector(5 downto 0);
signal VN22_data_out : std_logic_vector(5 downto 0);
signal VN22_sign_out : std_logic_vector(5 downto 0);
signal VN23_data_out : std_logic_vector(5 downto 0);
signal VN23_sign_out : std_logic_vector(5 downto 0);
signal VN24_data_out : std_logic_vector(5 downto 0);
signal VN24_sign_out : std_logic_vector(5 downto 0);
signal VN25_data_out : std_logic_vector(5 downto 0);
signal VN25_sign_out : std_logic_vector(5 downto 0);
signal VN26_data_out : std_logic_vector(5 downto 0);
signal VN26_sign_out : std_logic_vector(5 downto 0);
signal VN27_data_out : std_logic_vector(5 downto 0);
signal VN27_sign_out : std_logic_vector(5 downto 0);
signal VN28_data_out : std_logic_vector(5 downto 0);
signal VN28_sign_out : std_logic_vector(5 downto 0);
signal VN29_data_out : std_logic_vector(5 downto 0);
signal VN29_sign_out : std_logic_vector(5 downto 0);
signal VN30_data_out : std_logic_vector(5 downto 0);
signal VN30_sign_out : std_logic_vector(5 downto 0);
signal VN31_data_out : std_logic_vector(5 downto 0);
signal VN31_sign_out : std_logic_vector(5 downto 0);
signal VN32_data_out : std_logic_vector(5 downto 0);
signal VN32_sign_out : std_logic_vector(5 downto 0);
signal VN33_data_out : std_logic_vector(5 downto 0);
signal VN33_sign_out : std_logic_vector(5 downto 0);
signal VN34_data_out : std_logic_vector(5 downto 0);
signal VN34_sign_out : std_logic_vector(5 downto 0);
signal VN35_data_out : std_logic_vector(5 downto 0);
signal VN35_sign_out : std_logic_vector(5 downto 0);
signal VN36_data_out : std_logic_vector(5 downto 0);
signal VN36_sign_out : std_logic_vector(5 downto 0);
signal VN37_data_out : std_logic_vector(5 downto 0);
signal VN37_sign_out : std_logic_vector(5 downto 0);
signal VN38_data_out : std_logic_vector(5 downto 0);
signal VN38_sign_out : std_logic_vector(5 downto 0);
signal VN39_data_out : std_logic_vector(5 downto 0);
signal VN39_sign_out : std_logic_vector(5 downto 0);
signal VN40_data_out : std_logic_vector(5 downto 0);
signal VN40_sign_out : std_logic_vector(5 downto 0);
signal VN41_data_out : std_logic_vector(5 downto 0);
signal VN41_sign_out : std_logic_vector(5 downto 0);
signal VN42_data_out : std_logic_vector(5 downto 0);
signal VN42_sign_out : std_logic_vector(5 downto 0);
signal VN43_data_out : std_logic_vector(5 downto 0);
signal VN43_sign_out : std_logic_vector(5 downto 0);
signal VN44_data_out : std_logic_vector(5 downto 0);
signal VN44_sign_out : std_logic_vector(5 downto 0);
signal VN45_data_out : std_logic_vector(5 downto 0);
signal VN45_sign_out : std_logic_vector(5 downto 0);
signal VN46_data_out : std_logic_vector(5 downto 0);
signal VN46_sign_out : std_logic_vector(5 downto 0);
signal VN47_data_out : std_logic_vector(5 downto 0);
signal VN47_sign_out : std_logic_vector(5 downto 0);
signal VN48_data_out : std_logic_vector(5 downto 0);
signal VN48_sign_out : std_logic_vector(5 downto 0);
signal VN49_data_out : std_logic_vector(5 downto 0);
signal VN49_sign_out : std_logic_vector(5 downto 0);
signal VN50_data_out : std_logic_vector(5 downto 0);
signal VN50_sign_out : std_logic_vector(5 downto 0);
signal VN51_data_out : std_logic_vector(5 downto 0);
signal VN51_sign_out : std_logic_vector(5 downto 0);
signal VN52_data_out : std_logic_vector(5 downto 0);
signal VN52_sign_out : std_logic_vector(5 downto 0);
signal VN53_data_out : std_logic_vector(5 downto 0);
signal VN53_sign_out : std_logic_vector(5 downto 0);
signal VN54_data_out : std_logic_vector(5 downto 0);
signal VN54_sign_out : std_logic_vector(5 downto 0);
signal VN55_data_out : std_logic_vector(5 downto 0);
signal VN55_sign_out : std_logic_vector(5 downto 0);
signal VN56_data_out : std_logic_vector(5 downto 0);
signal VN56_sign_out : std_logic_vector(5 downto 0);
signal VN57_data_out : std_logic_vector(5 downto 0);
signal VN57_sign_out : std_logic_vector(5 downto 0);
signal VN58_data_out : std_logic_vector(5 downto 0);
signal VN58_sign_out : std_logic_vector(5 downto 0);
signal VN59_data_out : std_logic_vector(5 downto 0);
signal VN59_sign_out : std_logic_vector(5 downto 0);
signal VN60_data_out : std_logic_vector(5 downto 0);
signal VN60_sign_out : std_logic_vector(5 downto 0);
signal VN61_data_out : std_logic_vector(5 downto 0);
signal VN61_sign_out : std_logic_vector(5 downto 0);
signal VN62_data_out : std_logic_vector(5 downto 0);
signal VN62_sign_out : std_logic_vector(5 downto 0);
signal VN63_data_out : std_logic_vector(5 downto 0);
signal VN63_sign_out : std_logic_vector(5 downto 0);
signal VN64_data_out : std_logic_vector(5 downto 0);
signal VN64_sign_out : std_logic_vector(5 downto 0);
signal VN65_data_out : std_logic_vector(5 downto 0);
signal VN65_sign_out : std_logic_vector(5 downto 0);
signal VN66_data_out : std_logic_vector(5 downto 0);
signal VN66_sign_out : std_logic_vector(5 downto 0);
signal VN67_data_out : std_logic_vector(5 downto 0);
signal VN67_sign_out : std_logic_vector(5 downto 0);
signal VN68_data_out : std_logic_vector(5 downto 0);
signal VN68_sign_out : std_logic_vector(5 downto 0);
signal VN69_data_out : std_logic_vector(5 downto 0);
signal VN69_sign_out : std_logic_vector(5 downto 0);
signal VN70_data_out : std_logic_vector(5 downto 0);
signal VN70_sign_out : std_logic_vector(5 downto 0);
signal VN71_data_out : std_logic_vector(5 downto 0);
signal VN71_sign_out : std_logic_vector(5 downto 0);
signal VN72_data_out : std_logic_vector(5 downto 0);
signal VN72_sign_out : std_logic_vector(5 downto 0);
signal VN73_data_out : std_logic_vector(5 downto 0);
signal VN73_sign_out : std_logic_vector(5 downto 0);
signal VN74_data_out : std_logic_vector(5 downto 0);
signal VN74_sign_out : std_logic_vector(5 downto 0);
signal VN75_data_out : std_logic_vector(5 downto 0);
signal VN75_sign_out : std_logic_vector(5 downto 0);
signal VN76_data_out : std_logic_vector(5 downto 0);
signal VN76_sign_out : std_logic_vector(5 downto 0);
signal VN77_data_out : std_logic_vector(5 downto 0);
signal VN77_sign_out : std_logic_vector(5 downto 0);
signal VN78_data_out : std_logic_vector(5 downto 0);
signal VN78_sign_out : std_logic_vector(5 downto 0);
signal VN79_data_out : std_logic_vector(5 downto 0);
signal VN79_sign_out : std_logic_vector(5 downto 0);
signal VN80_data_out : std_logic_vector(5 downto 0);
signal VN80_sign_out : std_logic_vector(5 downto 0);
signal VN81_data_out : std_logic_vector(5 downto 0);
signal VN81_sign_out : std_logic_vector(5 downto 0);
signal VN82_data_out : std_logic_vector(5 downto 0);
signal VN82_sign_out : std_logic_vector(5 downto 0);
signal VN83_data_out : std_logic_vector(5 downto 0);
signal VN83_sign_out : std_logic_vector(5 downto 0);
signal VN84_data_out : std_logic_vector(5 downto 0);
signal VN84_sign_out : std_logic_vector(5 downto 0);
signal VN85_data_out : std_logic_vector(5 downto 0);
signal VN85_sign_out : std_logic_vector(5 downto 0);
signal VN86_data_out : std_logic_vector(5 downto 0);
signal VN86_sign_out : std_logic_vector(5 downto 0);
signal VN87_data_out : std_logic_vector(5 downto 0);
signal VN87_sign_out : std_logic_vector(5 downto 0);
signal VN88_data_out : std_logic_vector(5 downto 0);
signal VN88_sign_out : std_logic_vector(5 downto 0);
signal VN89_data_out : std_logic_vector(5 downto 0);
signal VN89_sign_out : std_logic_vector(5 downto 0);
signal VN90_data_out : std_logic_vector(5 downto 0);
signal VN90_sign_out : std_logic_vector(5 downto 0);
signal VN91_data_out : std_logic_vector(5 downto 0);
signal VN91_sign_out : std_logic_vector(5 downto 0);
signal VN92_data_out : std_logic_vector(5 downto 0);
signal VN92_sign_out : std_logic_vector(5 downto 0);
signal VN93_data_out : std_logic_vector(5 downto 0);
signal VN93_sign_out : std_logic_vector(5 downto 0);
signal VN94_data_out : std_logic_vector(5 downto 0);
signal VN94_sign_out : std_logic_vector(5 downto 0);
signal VN95_data_out : std_logic_vector(5 downto 0);
signal VN95_sign_out : std_logic_vector(5 downto 0);
signal VN96_data_out : std_logic_vector(5 downto 0);
signal VN96_sign_out : std_logic_vector(5 downto 0);
signal VN97_data_out : std_logic_vector(5 downto 0);
signal VN97_sign_out : std_logic_vector(5 downto 0);
signal VN98_data_out : std_logic_vector(5 downto 0);
signal VN98_sign_out : std_logic_vector(5 downto 0);
signal VN99_data_out : std_logic_vector(5 downto 0);
signal VN99_sign_out : std_logic_vector(5 downto 0);
signal VN100_data_out : std_logic_vector(5 downto 0);
signal VN100_sign_out : std_logic_vector(5 downto 0);
signal VN101_data_out : std_logic_vector(5 downto 0);
signal VN101_sign_out : std_logic_vector(5 downto 0);
signal VN102_data_out : std_logic_vector(5 downto 0);
signal VN102_sign_out : std_logic_vector(5 downto 0);
signal VN103_data_out : std_logic_vector(5 downto 0);
signal VN103_sign_out : std_logic_vector(5 downto 0);
signal VN104_data_out : std_logic_vector(5 downto 0);
signal VN104_sign_out : std_logic_vector(5 downto 0);
signal VN105_data_out : std_logic_vector(5 downto 0);
signal VN105_sign_out : std_logic_vector(5 downto 0);
signal VN106_data_out : std_logic_vector(5 downto 0);
signal VN106_sign_out : std_logic_vector(5 downto 0);
signal VN107_data_out : std_logic_vector(5 downto 0);
signal VN107_sign_out : std_logic_vector(5 downto 0);
signal VN108_data_out : std_logic_vector(5 downto 0);
signal VN108_sign_out : std_logic_vector(5 downto 0);
signal VN109_data_out : std_logic_vector(5 downto 0);
signal VN109_sign_out : std_logic_vector(5 downto 0);
signal VN110_data_out : std_logic_vector(5 downto 0);
signal VN110_sign_out : std_logic_vector(5 downto 0);
signal VN111_data_out : std_logic_vector(5 downto 0);
signal VN111_sign_out : std_logic_vector(5 downto 0);
signal VN112_data_out : std_logic_vector(5 downto 0);
signal VN112_sign_out : std_logic_vector(5 downto 0);
signal VN113_data_out : std_logic_vector(5 downto 0);
signal VN113_sign_out : std_logic_vector(5 downto 0);
signal VN114_data_out : std_logic_vector(5 downto 0);
signal VN114_sign_out : std_logic_vector(5 downto 0);
signal VN115_data_out : std_logic_vector(5 downto 0);
signal VN115_sign_out : std_logic_vector(5 downto 0);
signal VN116_data_out : std_logic_vector(5 downto 0);
signal VN116_sign_out : std_logic_vector(5 downto 0);
signal VN117_data_out : std_logic_vector(5 downto 0);
signal VN117_sign_out : std_logic_vector(5 downto 0);
signal VN118_data_out : std_logic_vector(5 downto 0);
signal VN118_sign_out : std_logic_vector(5 downto 0);
signal VN119_data_out : std_logic_vector(5 downto 0);
signal VN119_sign_out : std_logic_vector(5 downto 0);
signal VN120_data_out : std_logic_vector(5 downto 0);
signal VN120_sign_out : std_logic_vector(5 downto 0);
signal VN121_data_out : std_logic_vector(5 downto 0);
signal VN121_sign_out : std_logic_vector(5 downto 0);
signal VN122_data_out : std_logic_vector(5 downto 0);
signal VN122_sign_out : std_logic_vector(5 downto 0);
signal VN123_data_out : std_logic_vector(5 downto 0);
signal VN123_sign_out : std_logic_vector(5 downto 0);
signal VN124_data_out : std_logic_vector(5 downto 0);
signal VN124_sign_out : std_logic_vector(5 downto 0);
signal VN125_data_out : std_logic_vector(5 downto 0);
signal VN125_sign_out : std_logic_vector(5 downto 0);
signal VN126_data_out : std_logic_vector(5 downto 0);
signal VN126_sign_out : std_logic_vector(5 downto 0);
signal VN127_data_out : std_logic_vector(5 downto 0);
signal VN127_sign_out : std_logic_vector(5 downto 0);
signal VN128_data_out : std_logic_vector(5 downto 0);
signal VN128_sign_out : std_logic_vector(5 downto 0);
signal VN129_data_out : std_logic_vector(5 downto 0);
signal VN129_sign_out : std_logic_vector(5 downto 0);
signal VN130_data_out : std_logic_vector(5 downto 0);
signal VN130_sign_out : std_logic_vector(5 downto 0);
signal VN131_data_out : std_logic_vector(5 downto 0);
signal VN131_sign_out : std_logic_vector(5 downto 0);
signal VN132_data_out : std_logic_vector(5 downto 0);
signal VN132_sign_out : std_logic_vector(5 downto 0);
signal VN133_data_out : std_logic_vector(5 downto 0);
signal VN133_sign_out : std_logic_vector(5 downto 0);
signal VN134_data_out : std_logic_vector(5 downto 0);
signal VN134_sign_out : std_logic_vector(5 downto 0);
signal VN135_data_out : std_logic_vector(5 downto 0);
signal VN135_sign_out : std_logic_vector(5 downto 0);
signal VN136_data_out : std_logic_vector(5 downto 0);
signal VN136_sign_out : std_logic_vector(5 downto 0);
signal VN137_data_out : std_logic_vector(5 downto 0);
signal VN137_sign_out : std_logic_vector(5 downto 0);
signal VN138_data_out : std_logic_vector(5 downto 0);
signal VN138_sign_out : std_logic_vector(5 downto 0);
signal VN139_data_out : std_logic_vector(5 downto 0);
signal VN139_sign_out : std_logic_vector(5 downto 0);
signal VN140_data_out : std_logic_vector(5 downto 0);
signal VN140_sign_out : std_logic_vector(5 downto 0);
signal VN141_data_out : std_logic_vector(5 downto 0);
signal VN141_sign_out : std_logic_vector(5 downto 0);
signal VN142_data_out : std_logic_vector(5 downto 0);
signal VN142_sign_out : std_logic_vector(5 downto 0);
signal VN143_data_out : std_logic_vector(5 downto 0);
signal VN143_sign_out : std_logic_vector(5 downto 0);
signal VN144_data_out : std_logic_vector(5 downto 0);
signal VN144_sign_out : std_logic_vector(5 downto 0);
signal VN145_data_out : std_logic_vector(5 downto 0);
signal VN145_sign_out : std_logic_vector(5 downto 0);
signal VN146_data_out : std_logic_vector(5 downto 0);
signal VN146_sign_out : std_logic_vector(5 downto 0);
signal VN147_data_out : std_logic_vector(5 downto 0);
signal VN147_sign_out : std_logic_vector(5 downto 0);
signal VN148_data_out : std_logic_vector(5 downto 0);
signal VN148_sign_out : std_logic_vector(5 downto 0);
signal VN149_data_out : std_logic_vector(5 downto 0);
signal VN149_sign_out : std_logic_vector(5 downto 0);
signal VN150_data_out : std_logic_vector(5 downto 0);
signal VN150_sign_out : std_logic_vector(5 downto 0);
signal VN151_data_out : std_logic_vector(5 downto 0);
signal VN151_sign_out : std_logic_vector(5 downto 0);
signal VN152_data_out : std_logic_vector(5 downto 0);
signal VN152_sign_out : std_logic_vector(5 downto 0);
signal VN153_data_out : std_logic_vector(5 downto 0);
signal VN153_sign_out : std_logic_vector(5 downto 0);
signal VN154_data_out : std_logic_vector(5 downto 0);
signal VN154_sign_out : std_logic_vector(5 downto 0);
signal VN155_data_out : std_logic_vector(5 downto 0);
signal VN155_sign_out : std_logic_vector(5 downto 0);
signal VN156_data_out : std_logic_vector(5 downto 0);
signal VN156_sign_out : std_logic_vector(5 downto 0);
signal VN157_data_out : std_logic_vector(5 downto 0);
signal VN157_sign_out : std_logic_vector(5 downto 0);
signal VN158_data_out : std_logic_vector(5 downto 0);
signal VN158_sign_out : std_logic_vector(5 downto 0);
signal VN159_data_out : std_logic_vector(5 downto 0);
signal VN159_sign_out : std_logic_vector(5 downto 0);
signal VN160_data_out : std_logic_vector(5 downto 0);
signal VN160_sign_out : std_logic_vector(5 downto 0);
signal VN161_data_out : std_logic_vector(5 downto 0);
signal VN161_sign_out : std_logic_vector(5 downto 0);
signal VN162_data_out : std_logic_vector(5 downto 0);
signal VN162_sign_out : std_logic_vector(5 downto 0);
signal VN163_data_out : std_logic_vector(5 downto 0);
signal VN163_sign_out : std_logic_vector(5 downto 0);
signal VN164_data_out : std_logic_vector(5 downto 0);
signal VN164_sign_out : std_logic_vector(5 downto 0);
signal VN165_data_out : std_logic_vector(5 downto 0);
signal VN165_sign_out : std_logic_vector(5 downto 0);
signal VN166_data_out : std_logic_vector(5 downto 0);
signal VN166_sign_out : std_logic_vector(5 downto 0);
signal VN167_data_out : std_logic_vector(5 downto 0);
signal VN167_sign_out : std_logic_vector(5 downto 0);
signal VN168_data_out : std_logic_vector(5 downto 0);
signal VN168_sign_out : std_logic_vector(5 downto 0);
signal VN169_data_out : std_logic_vector(5 downto 0);
signal VN169_sign_out : std_logic_vector(5 downto 0);
signal VN170_data_out : std_logic_vector(5 downto 0);
signal VN170_sign_out : std_logic_vector(5 downto 0);
signal VN171_data_out : std_logic_vector(5 downto 0);
signal VN171_sign_out : std_logic_vector(5 downto 0);
signal VN172_data_out : std_logic_vector(5 downto 0);
signal VN172_sign_out : std_logic_vector(5 downto 0);
signal VN173_data_out : std_logic_vector(5 downto 0);
signal VN173_sign_out : std_logic_vector(5 downto 0);
signal VN174_data_out : std_logic_vector(5 downto 0);
signal VN174_sign_out : std_logic_vector(5 downto 0);
signal VN175_data_out : std_logic_vector(5 downto 0);
signal VN175_sign_out : std_logic_vector(5 downto 0);
signal VN176_data_out : std_logic_vector(5 downto 0);
signal VN176_sign_out : std_logic_vector(5 downto 0);
signal VN177_data_out : std_logic_vector(5 downto 0);
signal VN177_sign_out : std_logic_vector(5 downto 0);
signal VN178_data_out : std_logic_vector(5 downto 0);
signal VN178_sign_out : std_logic_vector(5 downto 0);
signal VN179_data_out : std_logic_vector(5 downto 0);
signal VN179_sign_out : std_logic_vector(5 downto 0);
signal VN180_data_out : std_logic_vector(5 downto 0);
signal VN180_sign_out : std_logic_vector(5 downto 0);
signal VN181_data_out : std_logic_vector(5 downto 0);
signal VN181_sign_out : std_logic_vector(5 downto 0);
signal VN182_data_out : std_logic_vector(5 downto 0);
signal VN182_sign_out : std_logic_vector(5 downto 0);
signal VN183_data_out : std_logic_vector(5 downto 0);
signal VN183_sign_out : std_logic_vector(5 downto 0);
signal VN184_data_out : std_logic_vector(5 downto 0);
signal VN184_sign_out : std_logic_vector(5 downto 0);
signal VN185_data_out : std_logic_vector(5 downto 0);
signal VN185_sign_out : std_logic_vector(5 downto 0);
signal VN186_data_out : std_logic_vector(5 downto 0);
signal VN186_sign_out : std_logic_vector(5 downto 0);
signal VN187_data_out : std_logic_vector(5 downto 0);
signal VN187_sign_out : std_logic_vector(5 downto 0);
signal VN188_data_out : std_logic_vector(5 downto 0);
signal VN188_sign_out : std_logic_vector(5 downto 0);
signal VN189_data_out : std_logic_vector(5 downto 0);
signal VN189_sign_out : std_logic_vector(5 downto 0);
signal VN190_data_out : std_logic_vector(5 downto 0);
signal VN190_sign_out : std_logic_vector(5 downto 0);
signal VN191_data_out : std_logic_vector(5 downto 0);
signal VN191_sign_out : std_logic_vector(5 downto 0);
signal VN192_data_out : std_logic_vector(5 downto 0);
signal VN192_sign_out : std_logic_vector(5 downto 0);
signal VN193_data_out : std_logic_vector(5 downto 0);
signal VN193_sign_out : std_logic_vector(5 downto 0);
signal VN194_data_out : std_logic_vector(5 downto 0);
signal VN194_sign_out : std_logic_vector(5 downto 0);
signal VN195_data_out : std_logic_vector(5 downto 0);
signal VN195_sign_out : std_logic_vector(5 downto 0);
signal VN196_data_out : std_logic_vector(5 downto 0);
signal VN196_sign_out : std_logic_vector(5 downto 0);
signal VN197_data_out : std_logic_vector(5 downto 0);
signal VN197_sign_out : std_logic_vector(5 downto 0);
signal VN198_data_out : std_logic_vector(5 downto 0);
signal VN198_sign_out : std_logic_vector(5 downto 0);
signal VN199_data_out : std_logic_vector(5 downto 0);
signal VN199_sign_out : std_logic_vector(5 downto 0);
signal VN200_data_out : std_logic_vector(5 downto 0);
signal VN200_sign_out : std_logic_vector(5 downto 0);
signal VN201_data_out : std_logic_vector(5 downto 0);
signal VN201_sign_out : std_logic_vector(5 downto 0);
signal VN202_data_out : std_logic_vector(5 downto 0);
signal VN202_sign_out : std_logic_vector(5 downto 0);
signal VN203_data_out : std_logic_vector(5 downto 0);
signal VN203_sign_out : std_logic_vector(5 downto 0);
signal VN204_data_out : std_logic_vector(5 downto 0);
signal VN204_sign_out : std_logic_vector(5 downto 0);
signal VN205_data_out : std_logic_vector(5 downto 0);
signal VN205_sign_out : std_logic_vector(5 downto 0);
signal VN206_data_out : std_logic_vector(5 downto 0);
signal VN206_sign_out : std_logic_vector(5 downto 0);
signal VN207_data_out : std_logic_vector(5 downto 0);
signal VN207_sign_out : std_logic_vector(5 downto 0);
signal VN208_data_out : std_logic_vector(5 downto 0);
signal VN208_sign_out : std_logic_vector(5 downto 0);
signal VN209_data_out : std_logic_vector(5 downto 0);
signal VN209_sign_out : std_logic_vector(5 downto 0);
signal VN210_data_out : std_logic_vector(5 downto 0);
signal VN210_sign_out : std_logic_vector(5 downto 0);
signal VN211_data_out : std_logic_vector(5 downto 0);
signal VN211_sign_out : std_logic_vector(5 downto 0);
signal VN212_data_out : std_logic_vector(5 downto 0);
signal VN212_sign_out : std_logic_vector(5 downto 0);
signal VN213_data_out : std_logic_vector(5 downto 0);
signal VN213_sign_out : std_logic_vector(5 downto 0);
signal VN214_data_out : std_logic_vector(5 downto 0);
signal VN214_sign_out : std_logic_vector(5 downto 0);
signal VN215_data_out : std_logic_vector(5 downto 0);
signal VN215_sign_out : std_logic_vector(5 downto 0);
signal VN216_data_out : std_logic_vector(5 downto 0);
signal VN216_sign_out : std_logic_vector(5 downto 0);
signal VN217_data_out : std_logic_vector(5 downto 0);
signal VN217_sign_out : std_logic_vector(5 downto 0);
signal VN218_data_out : std_logic_vector(5 downto 0);
signal VN218_sign_out : std_logic_vector(5 downto 0);
signal VN219_data_out : std_logic_vector(5 downto 0);
signal VN219_sign_out : std_logic_vector(5 downto 0);
signal VN220_data_out : std_logic_vector(5 downto 0);
signal VN220_sign_out : std_logic_vector(5 downto 0);
signal VN221_data_out : std_logic_vector(5 downto 0);
signal VN221_sign_out : std_logic_vector(5 downto 0);
signal VN222_data_out : std_logic_vector(5 downto 0);
signal VN222_sign_out : std_logic_vector(5 downto 0);
signal VN223_data_out : std_logic_vector(5 downto 0);
signal VN223_sign_out : std_logic_vector(5 downto 0);
signal VN224_data_out : std_logic_vector(5 downto 0);
signal VN224_sign_out : std_logic_vector(5 downto 0);
signal VN225_data_out : std_logic_vector(5 downto 0);
signal VN225_sign_out : std_logic_vector(5 downto 0);
signal VN226_data_out : std_logic_vector(5 downto 0);
signal VN226_sign_out : std_logic_vector(5 downto 0);
signal VN227_data_out : std_logic_vector(5 downto 0);
signal VN227_sign_out : std_logic_vector(5 downto 0);
signal VN228_data_out : std_logic_vector(5 downto 0);
signal VN228_sign_out : std_logic_vector(5 downto 0);
signal VN229_data_out : std_logic_vector(5 downto 0);
signal VN229_sign_out : std_logic_vector(5 downto 0);
signal VN230_data_out : std_logic_vector(5 downto 0);
signal VN230_sign_out : std_logic_vector(5 downto 0);
signal VN231_data_out : std_logic_vector(5 downto 0);
signal VN231_sign_out : std_logic_vector(5 downto 0);
signal VN232_data_out : std_logic_vector(5 downto 0);
signal VN232_sign_out : std_logic_vector(5 downto 0);
signal VN233_data_out : std_logic_vector(5 downto 0);
signal VN233_sign_out : std_logic_vector(5 downto 0);
signal VN234_data_out : std_logic_vector(5 downto 0);
signal VN234_sign_out : std_logic_vector(5 downto 0);
signal VN235_data_out : std_logic_vector(5 downto 0);
signal VN235_sign_out : std_logic_vector(5 downto 0);
signal VN236_data_out : std_logic_vector(5 downto 0);
signal VN236_sign_out : std_logic_vector(5 downto 0);
signal VN237_data_out : std_logic_vector(5 downto 0);
signal VN237_sign_out : std_logic_vector(5 downto 0);
signal VN238_data_out : std_logic_vector(5 downto 0);
signal VN238_sign_out : std_logic_vector(5 downto 0);
signal VN239_data_out : std_logic_vector(5 downto 0);
signal VN239_sign_out : std_logic_vector(5 downto 0);
signal VN240_data_out : std_logic_vector(5 downto 0);
signal VN240_sign_out : std_logic_vector(5 downto 0);
signal VN241_data_out : std_logic_vector(5 downto 0);
signal VN241_sign_out : std_logic_vector(5 downto 0);
signal VN242_data_out : std_logic_vector(5 downto 0);
signal VN242_sign_out : std_logic_vector(5 downto 0);
signal VN243_data_out : std_logic_vector(5 downto 0);
signal VN243_sign_out : std_logic_vector(5 downto 0);
signal VN244_data_out : std_logic_vector(5 downto 0);
signal VN244_sign_out : std_logic_vector(5 downto 0);
signal VN245_data_out : std_logic_vector(5 downto 0);
signal VN245_sign_out : std_logic_vector(5 downto 0);
signal VN246_data_out : std_logic_vector(5 downto 0);
signal VN246_sign_out : std_logic_vector(5 downto 0);
signal VN247_data_out : std_logic_vector(5 downto 0);
signal VN247_sign_out : std_logic_vector(5 downto 0);
signal VN248_data_out : std_logic_vector(5 downto 0);
signal VN248_sign_out : std_logic_vector(5 downto 0);
signal VN249_data_out : std_logic_vector(5 downto 0);
signal VN249_sign_out : std_logic_vector(5 downto 0);
signal VN250_data_out : std_logic_vector(5 downto 0);
signal VN250_sign_out : std_logic_vector(5 downto 0);
signal VN251_data_out : std_logic_vector(5 downto 0);
signal VN251_sign_out : std_logic_vector(5 downto 0);
signal VN252_data_out : std_logic_vector(5 downto 0);
signal VN252_sign_out : std_logic_vector(5 downto 0);
signal VN253_data_out : std_logic_vector(5 downto 0);
signal VN253_sign_out : std_logic_vector(5 downto 0);
signal VN254_data_out : std_logic_vector(5 downto 0);
signal VN254_sign_out : std_logic_vector(5 downto 0);
signal VN255_data_out : std_logic_vector(5 downto 0);
signal VN255_sign_out : std_logic_vector(5 downto 0);
signal VN256_data_out : std_logic_vector(5 downto 0);
signal VN256_sign_out : std_logic_vector(5 downto 0);
signal VN257_data_out : std_logic_vector(5 downto 0);
signal VN257_sign_out : std_logic_vector(5 downto 0);
signal VN258_data_out : std_logic_vector(5 downto 0);
signal VN258_sign_out : std_logic_vector(5 downto 0);
signal VN259_data_out : std_logic_vector(5 downto 0);
signal VN259_sign_out : std_logic_vector(5 downto 0);
signal VN260_data_out : std_logic_vector(5 downto 0);
signal VN260_sign_out : std_logic_vector(5 downto 0);
signal VN261_data_out : std_logic_vector(5 downto 0);
signal VN261_sign_out : std_logic_vector(5 downto 0);
signal VN262_data_out : std_logic_vector(5 downto 0);
signal VN262_sign_out : std_logic_vector(5 downto 0);
signal VN263_data_out : std_logic_vector(5 downto 0);
signal VN263_sign_out : std_logic_vector(5 downto 0);
signal VN264_data_out : std_logic_vector(5 downto 0);
signal VN264_sign_out : std_logic_vector(5 downto 0);
signal VN265_data_out : std_logic_vector(5 downto 0);
signal VN265_sign_out : std_logic_vector(5 downto 0);
signal VN266_data_out : std_logic_vector(5 downto 0);
signal VN266_sign_out : std_logic_vector(5 downto 0);
signal VN267_data_out : std_logic_vector(5 downto 0);
signal VN267_sign_out : std_logic_vector(5 downto 0);
signal VN268_data_out : std_logic_vector(5 downto 0);
signal VN268_sign_out : std_logic_vector(5 downto 0);
signal VN269_data_out : std_logic_vector(5 downto 0);
signal VN269_sign_out : std_logic_vector(5 downto 0);
signal VN270_data_out : std_logic_vector(5 downto 0);
signal VN270_sign_out : std_logic_vector(5 downto 0);
signal VN271_data_out : std_logic_vector(5 downto 0);
signal VN271_sign_out : std_logic_vector(5 downto 0);
signal VN272_data_out : std_logic_vector(5 downto 0);
signal VN272_sign_out : std_logic_vector(5 downto 0);
signal VN273_data_out : std_logic_vector(5 downto 0);
signal VN273_sign_out : std_logic_vector(5 downto 0);
signal VN274_data_out : std_logic_vector(5 downto 0);
signal VN274_sign_out : std_logic_vector(5 downto 0);
signal VN275_data_out : std_logic_vector(5 downto 0);
signal VN275_sign_out : std_logic_vector(5 downto 0);
signal VN276_data_out : std_logic_vector(5 downto 0);
signal VN276_sign_out : std_logic_vector(5 downto 0);
signal VN277_data_out : std_logic_vector(5 downto 0);
signal VN277_sign_out : std_logic_vector(5 downto 0);
signal VN278_data_out : std_logic_vector(5 downto 0);
signal VN278_sign_out : std_logic_vector(5 downto 0);
signal VN279_data_out : std_logic_vector(5 downto 0);
signal VN279_sign_out : std_logic_vector(5 downto 0);
signal VN280_data_out : std_logic_vector(5 downto 0);
signal VN280_sign_out : std_logic_vector(5 downto 0);
signal VN281_data_out : std_logic_vector(5 downto 0);
signal VN281_sign_out : std_logic_vector(5 downto 0);
signal VN282_data_out : std_logic_vector(5 downto 0);
signal VN282_sign_out : std_logic_vector(5 downto 0);
signal VN283_data_out : std_logic_vector(5 downto 0);
signal VN283_sign_out : std_logic_vector(5 downto 0);
signal VN284_data_out : std_logic_vector(5 downto 0);
signal VN284_sign_out : std_logic_vector(5 downto 0);
signal VN285_data_out : std_logic_vector(5 downto 0);
signal VN285_sign_out : std_logic_vector(5 downto 0);
signal VN286_data_out : std_logic_vector(5 downto 0);
signal VN286_sign_out : std_logic_vector(5 downto 0);
signal VN287_data_out : std_logic_vector(5 downto 0);
signal VN287_sign_out : std_logic_vector(5 downto 0);
signal VN288_data_out : std_logic_vector(5 downto 0);
signal VN288_sign_out : std_logic_vector(5 downto 0);
signal VN289_data_out : std_logic_vector(5 downto 0);
signal VN289_sign_out : std_logic_vector(5 downto 0);
signal VN290_data_out : std_logic_vector(5 downto 0);
signal VN290_sign_out : std_logic_vector(5 downto 0);
signal VN291_data_out : std_logic_vector(5 downto 0);
signal VN291_sign_out : std_logic_vector(5 downto 0);
signal VN292_data_out : std_logic_vector(5 downto 0);
signal VN292_sign_out : std_logic_vector(5 downto 0);
signal VN293_data_out : std_logic_vector(5 downto 0);
signal VN293_sign_out : std_logic_vector(5 downto 0);
signal VN294_data_out : std_logic_vector(5 downto 0);
signal VN294_sign_out : std_logic_vector(5 downto 0);
signal VN295_data_out : std_logic_vector(5 downto 0);
signal VN295_sign_out : std_logic_vector(5 downto 0);
signal VN296_data_out : std_logic_vector(5 downto 0);
signal VN296_sign_out : std_logic_vector(5 downto 0);
signal VN297_data_out : std_logic_vector(5 downto 0);
signal VN297_sign_out : std_logic_vector(5 downto 0);
signal VN298_data_out : std_logic_vector(5 downto 0);
signal VN298_sign_out : std_logic_vector(5 downto 0);
signal VN299_data_out : std_logic_vector(5 downto 0);
signal VN299_sign_out : std_logic_vector(5 downto 0);
signal VN300_data_out : std_logic_vector(5 downto 0);
signal VN300_sign_out : std_logic_vector(5 downto 0);
signal VN301_data_out : std_logic_vector(5 downto 0);
signal VN301_sign_out : std_logic_vector(5 downto 0);
signal VN302_data_out : std_logic_vector(5 downto 0);
signal VN302_sign_out : std_logic_vector(5 downto 0);
signal VN303_data_out : std_logic_vector(5 downto 0);
signal VN303_sign_out : std_logic_vector(5 downto 0);
signal VN304_data_out : std_logic_vector(5 downto 0);
signal VN304_sign_out : std_logic_vector(5 downto 0);
signal VN305_data_out : std_logic_vector(5 downto 0);
signal VN305_sign_out : std_logic_vector(5 downto 0);
signal VN306_data_out : std_logic_vector(5 downto 0);
signal VN306_sign_out : std_logic_vector(5 downto 0);
signal VN307_data_out : std_logic_vector(5 downto 0);
signal VN307_sign_out : std_logic_vector(5 downto 0);
signal VN308_data_out : std_logic_vector(5 downto 0);
signal VN308_sign_out : std_logic_vector(5 downto 0);
signal VN309_data_out : std_logic_vector(5 downto 0);
signal VN309_sign_out : std_logic_vector(5 downto 0);
signal VN310_data_out : std_logic_vector(5 downto 0);
signal VN310_sign_out : std_logic_vector(5 downto 0);
signal VN311_data_out : std_logic_vector(5 downto 0);
signal VN311_sign_out : std_logic_vector(5 downto 0);
signal VN312_data_out : std_logic_vector(5 downto 0);
signal VN312_sign_out : std_logic_vector(5 downto 0);
signal VN313_data_out : std_logic_vector(5 downto 0);
signal VN313_sign_out : std_logic_vector(5 downto 0);
signal VN314_data_out : std_logic_vector(5 downto 0);
signal VN314_sign_out : std_logic_vector(5 downto 0);
signal VN315_data_out : std_logic_vector(5 downto 0);
signal VN315_sign_out : std_logic_vector(5 downto 0);
signal VN316_data_out : std_logic_vector(5 downto 0);
signal VN316_sign_out : std_logic_vector(5 downto 0);
signal VN317_data_out : std_logic_vector(5 downto 0);
signal VN317_sign_out : std_logic_vector(5 downto 0);
signal VN318_data_out : std_logic_vector(5 downto 0);
signal VN318_sign_out : std_logic_vector(5 downto 0);
signal VN319_data_out : std_logic_vector(5 downto 0);
signal VN319_sign_out : std_logic_vector(5 downto 0);
signal VN320_data_out : std_logic_vector(5 downto 0);
signal VN320_sign_out : std_logic_vector(5 downto 0);
signal VN321_data_out : std_logic_vector(5 downto 0);
signal VN321_sign_out : std_logic_vector(5 downto 0);
signal VN322_data_out : std_logic_vector(5 downto 0);
signal VN322_sign_out : std_logic_vector(5 downto 0);
signal VN323_data_out : std_logic_vector(5 downto 0);
signal VN323_sign_out : std_logic_vector(5 downto 0);
signal VN324_data_out : std_logic_vector(5 downto 0);
signal VN324_sign_out : std_logic_vector(5 downto 0);
signal VN325_data_out : std_logic_vector(5 downto 0);
signal VN325_sign_out : std_logic_vector(5 downto 0);
signal VN326_data_out : std_logic_vector(5 downto 0);
signal VN326_sign_out : std_logic_vector(5 downto 0);
signal VN327_data_out : std_logic_vector(5 downto 0);
signal VN327_sign_out : std_logic_vector(5 downto 0);
signal VN328_data_out : std_logic_vector(5 downto 0);
signal VN328_sign_out : std_logic_vector(5 downto 0);
signal VN329_data_out : std_logic_vector(5 downto 0);
signal VN329_sign_out : std_logic_vector(5 downto 0);
signal VN330_data_out : std_logic_vector(5 downto 0);
signal VN330_sign_out : std_logic_vector(5 downto 0);
signal VN331_data_out : std_logic_vector(5 downto 0);
signal VN331_sign_out : std_logic_vector(5 downto 0);
signal VN332_data_out : std_logic_vector(5 downto 0);
signal VN332_sign_out : std_logic_vector(5 downto 0);
signal VN333_data_out : std_logic_vector(5 downto 0);
signal VN333_sign_out : std_logic_vector(5 downto 0);
signal VN334_data_out : std_logic_vector(5 downto 0);
signal VN334_sign_out : std_logic_vector(5 downto 0);
signal VN335_data_out : std_logic_vector(5 downto 0);
signal VN335_sign_out : std_logic_vector(5 downto 0);
signal VN336_data_out : std_logic_vector(5 downto 0);
signal VN336_sign_out : std_logic_vector(5 downto 0);
signal VN337_data_out : std_logic_vector(5 downto 0);
signal VN337_sign_out : std_logic_vector(5 downto 0);
signal VN338_data_out : std_logic_vector(5 downto 0);
signal VN338_sign_out : std_logic_vector(5 downto 0);
signal VN339_data_out : std_logic_vector(5 downto 0);
signal VN339_sign_out : std_logic_vector(5 downto 0);
signal VN340_data_out : std_logic_vector(5 downto 0);
signal VN340_sign_out : std_logic_vector(5 downto 0);
signal VN341_data_out : std_logic_vector(5 downto 0);
signal VN341_sign_out : std_logic_vector(5 downto 0);
signal VN342_data_out : std_logic_vector(5 downto 0);
signal VN342_sign_out : std_logic_vector(5 downto 0);
signal VN343_data_out : std_logic_vector(5 downto 0);
signal VN343_sign_out : std_logic_vector(5 downto 0);
signal VN344_data_out : std_logic_vector(5 downto 0);
signal VN344_sign_out : std_logic_vector(5 downto 0);
signal VN345_data_out : std_logic_vector(5 downto 0);
signal VN345_sign_out : std_logic_vector(5 downto 0);
signal VN346_data_out : std_logic_vector(5 downto 0);
signal VN346_sign_out : std_logic_vector(5 downto 0);
signal VN347_data_out : std_logic_vector(5 downto 0);
signal VN347_sign_out : std_logic_vector(5 downto 0);
signal VN348_data_out : std_logic_vector(5 downto 0);
signal VN348_sign_out : std_logic_vector(5 downto 0);
signal VN349_data_out : std_logic_vector(5 downto 0);
signal VN349_sign_out : std_logic_vector(5 downto 0);
signal VN350_data_out : std_logic_vector(5 downto 0);
signal VN350_sign_out : std_logic_vector(5 downto 0);
signal VN351_data_out : std_logic_vector(5 downto 0);
signal VN351_sign_out : std_logic_vector(5 downto 0);
signal VN352_data_out : std_logic_vector(5 downto 0);
signal VN352_sign_out : std_logic_vector(5 downto 0);
signal VN353_data_out : std_logic_vector(5 downto 0);
signal VN353_sign_out : std_logic_vector(5 downto 0);
signal VN354_data_out : std_logic_vector(5 downto 0);
signal VN354_sign_out : std_logic_vector(5 downto 0);
signal VN355_data_out : std_logic_vector(5 downto 0);
signal VN355_sign_out : std_logic_vector(5 downto 0);
signal VN356_data_out : std_logic_vector(5 downto 0);
signal VN356_sign_out : std_logic_vector(5 downto 0);
signal VN357_data_out : std_logic_vector(5 downto 0);
signal VN357_sign_out : std_logic_vector(5 downto 0);
signal VN358_data_out : std_logic_vector(5 downto 0);
signal VN358_sign_out : std_logic_vector(5 downto 0);
signal VN359_data_out : std_logic_vector(5 downto 0);
signal VN359_sign_out : std_logic_vector(5 downto 0);
signal VN360_data_out : std_logic_vector(5 downto 0);
signal VN360_sign_out : std_logic_vector(5 downto 0);
signal VN361_data_out : std_logic_vector(5 downto 0);
signal VN361_sign_out : std_logic_vector(5 downto 0);
signal VN362_data_out : std_logic_vector(5 downto 0);
signal VN362_sign_out : std_logic_vector(5 downto 0);
signal VN363_data_out : std_logic_vector(5 downto 0);
signal VN363_sign_out : std_logic_vector(5 downto 0);
signal VN364_data_out : std_logic_vector(5 downto 0);
signal VN364_sign_out : std_logic_vector(5 downto 0);
signal VN365_data_out : std_logic_vector(5 downto 0);
signal VN365_sign_out : std_logic_vector(5 downto 0);
signal VN366_data_out : std_logic_vector(5 downto 0);
signal VN366_sign_out : std_logic_vector(5 downto 0);
signal VN367_data_out : std_logic_vector(5 downto 0);
signal VN367_sign_out : std_logic_vector(5 downto 0);
signal VN368_data_out : std_logic_vector(5 downto 0);
signal VN368_sign_out : std_logic_vector(5 downto 0);
signal VN369_data_out : std_logic_vector(5 downto 0);
signal VN369_sign_out : std_logic_vector(5 downto 0);
signal VN370_data_out : std_logic_vector(5 downto 0);
signal VN370_sign_out : std_logic_vector(5 downto 0);
signal VN371_data_out : std_logic_vector(5 downto 0);
signal VN371_sign_out : std_logic_vector(5 downto 0);
signal VN372_data_out : std_logic_vector(5 downto 0);
signal VN372_sign_out : std_logic_vector(5 downto 0);
signal VN373_data_out : std_logic_vector(5 downto 0);
signal VN373_sign_out : std_logic_vector(5 downto 0);
signal VN374_data_out : std_logic_vector(5 downto 0);
signal VN374_sign_out : std_logic_vector(5 downto 0);
signal VN375_data_out : std_logic_vector(5 downto 0);
signal VN375_sign_out : std_logic_vector(5 downto 0);
signal VN376_data_out : std_logic_vector(5 downto 0);
signal VN376_sign_out : std_logic_vector(5 downto 0);
signal VN377_data_out : std_logic_vector(5 downto 0);
signal VN377_sign_out : std_logic_vector(5 downto 0);
signal VN378_data_out : std_logic_vector(5 downto 0);
signal VN378_sign_out : std_logic_vector(5 downto 0);
signal VN379_data_out : std_logic_vector(5 downto 0);
signal VN379_sign_out : std_logic_vector(5 downto 0);
signal VN380_data_out : std_logic_vector(5 downto 0);
signal VN380_sign_out : std_logic_vector(5 downto 0);
signal VN381_data_out : std_logic_vector(5 downto 0);
signal VN381_sign_out : std_logic_vector(5 downto 0);
signal VN382_data_out : std_logic_vector(5 downto 0);
signal VN382_sign_out : std_logic_vector(5 downto 0);
signal VN383_data_out : std_logic_vector(5 downto 0);
signal VN383_sign_out : std_logic_vector(5 downto 0);
signal VN384_data_out : std_logic_vector(5 downto 0);
signal VN384_sign_out : std_logic_vector(5 downto 0);
signal VN385_data_out : std_logic_vector(5 downto 0);
signal VN385_sign_out : std_logic_vector(5 downto 0);
signal VN386_data_out : std_logic_vector(5 downto 0);
signal VN386_sign_out : std_logic_vector(5 downto 0);
signal VN387_data_out : std_logic_vector(5 downto 0);
signal VN387_sign_out : std_logic_vector(5 downto 0);
signal VN388_data_out : std_logic_vector(5 downto 0);
signal VN388_sign_out : std_logic_vector(5 downto 0);
signal VN389_data_out : std_logic_vector(5 downto 0);
signal VN389_sign_out : std_logic_vector(5 downto 0);
signal VN390_data_out : std_logic_vector(5 downto 0);
signal VN390_sign_out : std_logic_vector(5 downto 0);
signal VN391_data_out : std_logic_vector(5 downto 0);
signal VN391_sign_out : std_logic_vector(5 downto 0);
signal VN392_data_out : std_logic_vector(5 downto 0);
signal VN392_sign_out : std_logic_vector(5 downto 0);
signal VN393_data_out : std_logic_vector(5 downto 0);
signal VN393_sign_out : std_logic_vector(5 downto 0);
signal VN394_data_out : std_logic_vector(5 downto 0);
signal VN394_sign_out : std_logic_vector(5 downto 0);
signal VN395_data_out : std_logic_vector(5 downto 0);
signal VN395_sign_out : std_logic_vector(5 downto 0);
signal VN396_data_out : std_logic_vector(5 downto 0);
signal VN396_sign_out : std_logic_vector(5 downto 0);
signal VN397_data_out : std_logic_vector(5 downto 0);
signal VN397_sign_out : std_logic_vector(5 downto 0);
signal VN398_data_out : std_logic_vector(5 downto 0);
signal VN398_sign_out : std_logic_vector(5 downto 0);
signal VN399_data_out : std_logic_vector(5 downto 0);
signal VN399_sign_out : std_logic_vector(5 downto 0);
signal VN400_data_out : std_logic_vector(5 downto 0);
signal VN400_sign_out : std_logic_vector(5 downto 0);
signal VN401_data_out : std_logic_vector(5 downto 0);
signal VN401_sign_out : std_logic_vector(5 downto 0);
signal VN402_data_out : std_logic_vector(5 downto 0);
signal VN402_sign_out : std_logic_vector(5 downto 0);
signal VN403_data_out : std_logic_vector(5 downto 0);
signal VN403_sign_out : std_logic_vector(5 downto 0);
signal VN404_data_out : std_logic_vector(5 downto 0);
signal VN404_sign_out : std_logic_vector(5 downto 0);
signal VN405_data_out : std_logic_vector(5 downto 0);
signal VN405_sign_out : std_logic_vector(5 downto 0);
signal VN406_data_out : std_logic_vector(5 downto 0);
signal VN406_sign_out : std_logic_vector(5 downto 0);
signal VN407_data_out : std_logic_vector(5 downto 0);
signal VN407_sign_out : std_logic_vector(5 downto 0);
signal VN408_data_out : std_logic_vector(5 downto 0);
signal VN408_sign_out : std_logic_vector(5 downto 0);
signal VN409_data_out : std_logic_vector(5 downto 0);
signal VN409_sign_out : std_logic_vector(5 downto 0);
signal VN410_data_out : std_logic_vector(5 downto 0);
signal VN410_sign_out : std_logic_vector(5 downto 0);
signal VN411_data_out : std_logic_vector(5 downto 0);
signal VN411_sign_out : std_logic_vector(5 downto 0);
signal VN412_data_out : std_logic_vector(5 downto 0);
signal VN412_sign_out : std_logic_vector(5 downto 0);
signal VN413_data_out : std_logic_vector(5 downto 0);
signal VN413_sign_out : std_logic_vector(5 downto 0);
signal VN414_data_out : std_logic_vector(5 downto 0);
signal VN414_sign_out : std_logic_vector(5 downto 0);
signal VN415_data_out : std_logic_vector(5 downto 0);
signal VN415_sign_out : std_logic_vector(5 downto 0);
signal VN416_data_out : std_logic_vector(5 downto 0);
signal VN416_sign_out : std_logic_vector(5 downto 0);
signal VN417_data_out : std_logic_vector(5 downto 0);
signal VN417_sign_out : std_logic_vector(5 downto 0);
signal VN418_data_out : std_logic_vector(5 downto 0);
signal VN418_sign_out : std_logic_vector(5 downto 0);
signal VN419_data_out : std_logic_vector(5 downto 0);
signal VN419_sign_out : std_logic_vector(5 downto 0);
signal VN420_data_out : std_logic_vector(5 downto 0);
signal VN420_sign_out : std_logic_vector(5 downto 0);
signal VN421_data_out : std_logic_vector(5 downto 0);
signal VN421_sign_out : std_logic_vector(5 downto 0);
signal VN422_data_out : std_logic_vector(5 downto 0);
signal VN422_sign_out : std_logic_vector(5 downto 0);
signal VN423_data_out : std_logic_vector(5 downto 0);
signal VN423_sign_out : std_logic_vector(5 downto 0);
signal VN424_data_out : std_logic_vector(5 downto 0);
signal VN424_sign_out : std_logic_vector(5 downto 0);
signal VN425_data_out : std_logic_vector(5 downto 0);
signal VN425_sign_out : std_logic_vector(5 downto 0);
signal VN426_data_out : std_logic_vector(5 downto 0);
signal VN426_sign_out : std_logic_vector(5 downto 0);
signal VN427_data_out : std_logic_vector(5 downto 0);
signal VN427_sign_out : std_logic_vector(5 downto 0);
signal VN428_data_out : std_logic_vector(5 downto 0);
signal VN428_sign_out : std_logic_vector(5 downto 0);
signal VN429_data_out : std_logic_vector(5 downto 0);
signal VN429_sign_out : std_logic_vector(5 downto 0);
signal VN430_data_out : std_logic_vector(5 downto 0);
signal VN430_sign_out : std_logic_vector(5 downto 0);
signal VN431_data_out : std_logic_vector(5 downto 0);
signal VN431_sign_out : std_logic_vector(5 downto 0);
signal VN432_data_out : std_logic_vector(5 downto 0);
signal VN432_sign_out : std_logic_vector(5 downto 0);
signal VN433_data_out : std_logic_vector(5 downto 0);
signal VN433_sign_out : std_logic_vector(5 downto 0);
signal VN434_data_out : std_logic_vector(5 downto 0);
signal VN434_sign_out : std_logic_vector(5 downto 0);
signal VN435_data_out : std_logic_vector(5 downto 0);
signal VN435_sign_out : std_logic_vector(5 downto 0);
signal VN436_data_out : std_logic_vector(5 downto 0);
signal VN436_sign_out : std_logic_vector(5 downto 0);
signal VN437_data_out : std_logic_vector(5 downto 0);
signal VN437_sign_out : std_logic_vector(5 downto 0);
signal VN438_data_out : std_logic_vector(5 downto 0);
signal VN438_sign_out : std_logic_vector(5 downto 0);
signal VN439_data_out : std_logic_vector(5 downto 0);
signal VN439_sign_out : std_logic_vector(5 downto 0);
signal VN440_data_out : std_logic_vector(5 downto 0);
signal VN440_sign_out : std_logic_vector(5 downto 0);
signal VN441_data_out : std_logic_vector(5 downto 0);
signal VN441_sign_out : std_logic_vector(5 downto 0);
signal VN442_data_out : std_logic_vector(5 downto 0);
signal VN442_sign_out : std_logic_vector(5 downto 0);
signal VN443_data_out : std_logic_vector(5 downto 0);
signal VN443_sign_out : std_logic_vector(5 downto 0);
signal VN444_data_out : std_logic_vector(5 downto 0);
signal VN444_sign_out : std_logic_vector(5 downto 0);
signal VN445_data_out : std_logic_vector(5 downto 0);
signal VN445_sign_out : std_logic_vector(5 downto 0);
signal VN446_data_out : std_logic_vector(5 downto 0);
signal VN446_sign_out : std_logic_vector(5 downto 0);
signal VN447_data_out : std_logic_vector(5 downto 0);
signal VN447_sign_out : std_logic_vector(5 downto 0);
signal VN448_data_out : std_logic_vector(5 downto 0);
signal VN448_sign_out : std_logic_vector(5 downto 0);
signal VN449_data_out : std_logic_vector(5 downto 0);
signal VN449_sign_out : std_logic_vector(5 downto 0);
signal VN450_data_out : std_logic_vector(5 downto 0);
signal VN450_sign_out : std_logic_vector(5 downto 0);
signal VN451_data_out : std_logic_vector(5 downto 0);
signal VN451_sign_out : std_logic_vector(5 downto 0);
signal VN452_data_out : std_logic_vector(5 downto 0);
signal VN452_sign_out : std_logic_vector(5 downto 0);
signal VN453_data_out : std_logic_vector(5 downto 0);
signal VN453_sign_out : std_logic_vector(5 downto 0);
signal VN454_data_out : std_logic_vector(5 downto 0);
signal VN454_sign_out : std_logic_vector(5 downto 0);
signal VN455_data_out : std_logic_vector(5 downto 0);
signal VN455_sign_out : std_logic_vector(5 downto 0);
signal VN456_data_out : std_logic_vector(5 downto 0);
signal VN456_sign_out : std_logic_vector(5 downto 0);
signal VN457_data_out : std_logic_vector(5 downto 0);
signal VN457_sign_out : std_logic_vector(5 downto 0);
signal VN458_data_out : std_logic_vector(5 downto 0);
signal VN458_sign_out : std_logic_vector(5 downto 0);
signal VN459_data_out : std_logic_vector(5 downto 0);
signal VN459_sign_out : std_logic_vector(5 downto 0);
signal VN460_data_out : std_logic_vector(5 downto 0);
signal VN460_sign_out : std_logic_vector(5 downto 0);
signal VN461_data_out : std_logic_vector(5 downto 0);
signal VN461_sign_out : std_logic_vector(5 downto 0);
signal VN462_data_out : std_logic_vector(5 downto 0);
signal VN462_sign_out : std_logic_vector(5 downto 0);
signal VN463_data_out : std_logic_vector(5 downto 0);
signal VN463_sign_out : std_logic_vector(5 downto 0);
signal VN464_data_out : std_logic_vector(5 downto 0);
signal VN464_sign_out : std_logic_vector(5 downto 0);
signal VN465_data_out : std_logic_vector(5 downto 0);
signal VN465_sign_out : std_logic_vector(5 downto 0);
signal VN466_data_out : std_logic_vector(5 downto 0);
signal VN466_sign_out : std_logic_vector(5 downto 0);
signal VN467_data_out : std_logic_vector(5 downto 0);
signal VN467_sign_out : std_logic_vector(5 downto 0);
signal VN468_data_out : std_logic_vector(5 downto 0);
signal VN468_sign_out : std_logic_vector(5 downto 0);
signal VN469_data_out : std_logic_vector(5 downto 0);
signal VN469_sign_out : std_logic_vector(5 downto 0);
signal VN470_data_out : std_logic_vector(5 downto 0);
signal VN470_sign_out : std_logic_vector(5 downto 0);
signal VN471_data_out : std_logic_vector(5 downto 0);
signal VN471_sign_out : std_logic_vector(5 downto 0);
signal VN472_data_out : std_logic_vector(5 downto 0);
signal VN472_sign_out : std_logic_vector(5 downto 0);
signal VN473_data_out : std_logic_vector(5 downto 0);
signal VN473_sign_out : std_logic_vector(5 downto 0);
signal VN474_data_out : std_logic_vector(5 downto 0);
signal VN474_sign_out : std_logic_vector(5 downto 0);
signal VN475_data_out : std_logic_vector(5 downto 0);
signal VN475_sign_out : std_logic_vector(5 downto 0);
signal VN476_data_out : std_logic_vector(5 downto 0);
signal VN476_sign_out : std_logic_vector(5 downto 0);
signal VN477_data_out : std_logic_vector(5 downto 0);
signal VN477_sign_out : std_logic_vector(5 downto 0);
signal VN478_data_out : std_logic_vector(5 downto 0);
signal VN478_sign_out : std_logic_vector(5 downto 0);
signal VN479_data_out : std_logic_vector(5 downto 0);
signal VN479_sign_out : std_logic_vector(5 downto 0);
signal VN480_data_out : std_logic_vector(5 downto 0);
signal VN480_sign_out : std_logic_vector(5 downto 0);
signal VN481_data_out : std_logic_vector(5 downto 0);
signal VN481_sign_out : std_logic_vector(5 downto 0);
signal VN482_data_out : std_logic_vector(5 downto 0);
signal VN482_sign_out : std_logic_vector(5 downto 0);
signal VN483_data_out : std_logic_vector(5 downto 0);
signal VN483_sign_out : std_logic_vector(5 downto 0);
signal VN484_data_out : std_logic_vector(5 downto 0);
signal VN484_sign_out : std_logic_vector(5 downto 0);
signal VN485_data_out : std_logic_vector(5 downto 0);
signal VN485_sign_out : std_logic_vector(5 downto 0);
signal VN486_data_out : std_logic_vector(5 downto 0);
signal VN486_sign_out : std_logic_vector(5 downto 0);
signal VN487_data_out : std_logic_vector(5 downto 0);
signal VN487_sign_out : std_logic_vector(5 downto 0);
signal VN488_data_out : std_logic_vector(5 downto 0);
signal VN488_sign_out : std_logic_vector(5 downto 0);
signal VN489_data_out : std_logic_vector(5 downto 0);
signal VN489_sign_out : std_logic_vector(5 downto 0);
signal VN490_data_out : std_logic_vector(5 downto 0);
signal VN490_sign_out : std_logic_vector(5 downto 0);
signal VN491_data_out : std_logic_vector(5 downto 0);
signal VN491_sign_out : std_logic_vector(5 downto 0);
signal VN492_data_out : std_logic_vector(5 downto 0);
signal VN492_sign_out : std_logic_vector(5 downto 0);
signal VN493_data_out : std_logic_vector(5 downto 0);
signal VN493_sign_out : std_logic_vector(5 downto 0);
signal VN494_data_out : std_logic_vector(5 downto 0);
signal VN494_sign_out : std_logic_vector(5 downto 0);
signal VN495_data_out : std_logic_vector(5 downto 0);
signal VN495_sign_out : std_logic_vector(5 downto 0);
signal VN496_data_out : std_logic_vector(5 downto 0);
signal VN496_sign_out : std_logic_vector(5 downto 0);
signal VN497_data_out : std_logic_vector(5 downto 0);
signal VN497_sign_out : std_logic_vector(5 downto 0);
signal VN498_data_out : std_logic_vector(5 downto 0);
signal VN498_sign_out : std_logic_vector(5 downto 0);
signal VN499_data_out : std_logic_vector(5 downto 0);
signal VN499_sign_out : std_logic_vector(5 downto 0);
signal VN500_data_out : std_logic_vector(5 downto 0);
signal VN500_sign_out : std_logic_vector(5 downto 0);
signal VN501_data_out : std_logic_vector(5 downto 0);
signal VN501_sign_out : std_logic_vector(5 downto 0);
signal VN502_data_out : std_logic_vector(5 downto 0);
signal VN502_sign_out : std_logic_vector(5 downto 0);
signal VN503_data_out : std_logic_vector(5 downto 0);
signal VN503_sign_out : std_logic_vector(5 downto 0);
signal VN504_data_out : std_logic_vector(5 downto 0);
signal VN504_sign_out : std_logic_vector(5 downto 0);
signal VN505_data_out : std_logic_vector(5 downto 0);
signal VN505_sign_out : std_logic_vector(5 downto 0);
signal VN506_data_out : std_logic_vector(5 downto 0);
signal VN506_sign_out : std_logic_vector(5 downto 0);
signal VN507_data_out : std_logic_vector(5 downto 0);
signal VN507_sign_out : std_logic_vector(5 downto 0);
signal VN508_data_out : std_logic_vector(5 downto 0);
signal VN508_sign_out : std_logic_vector(5 downto 0);
signal VN509_data_out : std_logic_vector(5 downto 0);
signal VN509_sign_out : std_logic_vector(5 downto 0);
signal VN510_data_out : std_logic_vector(5 downto 0);
signal VN510_sign_out : std_logic_vector(5 downto 0);
signal VN511_data_out : std_logic_vector(5 downto 0);
signal VN511_sign_out : std_logic_vector(5 downto 0);
signal VN512_data_out : std_logic_vector(5 downto 0);
signal VN512_sign_out : std_logic_vector(5 downto 0);
signal VN513_data_out : std_logic_vector(5 downto 0);
signal VN513_sign_out : std_logic_vector(5 downto 0);
signal VN514_data_out : std_logic_vector(5 downto 0);
signal VN514_sign_out : std_logic_vector(5 downto 0);
signal VN515_data_out : std_logic_vector(5 downto 0);
signal VN515_sign_out : std_logic_vector(5 downto 0);
signal VN516_data_out : std_logic_vector(5 downto 0);
signal VN516_sign_out : std_logic_vector(5 downto 0);
signal VN517_data_out : std_logic_vector(5 downto 0);
signal VN517_sign_out : std_logic_vector(5 downto 0);
signal VN518_data_out : std_logic_vector(5 downto 0);
signal VN518_sign_out : std_logic_vector(5 downto 0);
signal VN519_data_out : std_logic_vector(5 downto 0);
signal VN519_sign_out : std_logic_vector(5 downto 0);
signal VN520_data_out : std_logic_vector(5 downto 0);
signal VN520_sign_out : std_logic_vector(5 downto 0);
signal VN521_data_out : std_logic_vector(5 downto 0);
signal VN521_sign_out : std_logic_vector(5 downto 0);
signal VN522_data_out : std_logic_vector(5 downto 0);
signal VN522_sign_out : std_logic_vector(5 downto 0);
signal VN523_data_out : std_logic_vector(5 downto 0);
signal VN523_sign_out : std_logic_vector(5 downto 0);
signal VN524_data_out : std_logic_vector(5 downto 0);
signal VN524_sign_out : std_logic_vector(5 downto 0);
signal VN525_data_out : std_logic_vector(5 downto 0);
signal VN525_sign_out : std_logic_vector(5 downto 0);
signal VN526_data_out : std_logic_vector(5 downto 0);
signal VN526_sign_out : std_logic_vector(5 downto 0);
signal VN527_data_out : std_logic_vector(5 downto 0);
signal VN527_sign_out : std_logic_vector(5 downto 0);
signal VN528_data_out : std_logic_vector(5 downto 0);
signal VN528_sign_out : std_logic_vector(5 downto 0);
signal VN529_data_out : std_logic_vector(5 downto 0);
signal VN529_sign_out : std_logic_vector(5 downto 0);
signal VN530_data_out : std_logic_vector(5 downto 0);
signal VN530_sign_out : std_logic_vector(5 downto 0);
signal VN531_data_out : std_logic_vector(5 downto 0);
signal VN531_sign_out : std_logic_vector(5 downto 0);
signal VN532_data_out : std_logic_vector(5 downto 0);
signal VN532_sign_out : std_logic_vector(5 downto 0);
signal VN533_data_out : std_logic_vector(5 downto 0);
signal VN533_sign_out : std_logic_vector(5 downto 0);
signal VN534_data_out : std_logic_vector(5 downto 0);
signal VN534_sign_out : std_logic_vector(5 downto 0);
signal VN535_data_out : std_logic_vector(5 downto 0);
signal VN535_sign_out : std_logic_vector(5 downto 0);
signal VN536_data_out : std_logic_vector(5 downto 0);
signal VN536_sign_out : std_logic_vector(5 downto 0);
signal VN537_data_out : std_logic_vector(5 downto 0);
signal VN537_sign_out : std_logic_vector(5 downto 0);
signal VN538_data_out : std_logic_vector(5 downto 0);
signal VN538_sign_out : std_logic_vector(5 downto 0);
signal VN539_data_out : std_logic_vector(5 downto 0);
signal VN539_sign_out : std_logic_vector(5 downto 0);
signal VN540_data_out : std_logic_vector(5 downto 0);
signal VN540_sign_out : std_logic_vector(5 downto 0);
signal VN541_data_out : std_logic_vector(5 downto 0);
signal VN541_sign_out : std_logic_vector(5 downto 0);
signal VN542_data_out : std_logic_vector(5 downto 0);
signal VN542_sign_out : std_logic_vector(5 downto 0);
signal VN543_data_out : std_logic_vector(5 downto 0);
signal VN543_sign_out : std_logic_vector(5 downto 0);
signal VN544_data_out : std_logic_vector(5 downto 0);
signal VN544_sign_out : std_logic_vector(5 downto 0);
signal VN545_data_out : std_logic_vector(5 downto 0);
signal VN545_sign_out : std_logic_vector(5 downto 0);
signal VN546_data_out : std_logic_vector(5 downto 0);
signal VN546_sign_out : std_logic_vector(5 downto 0);
signal VN547_data_out : std_logic_vector(5 downto 0);
signal VN547_sign_out : std_logic_vector(5 downto 0);
signal VN548_data_out : std_logic_vector(5 downto 0);
signal VN548_sign_out : std_logic_vector(5 downto 0);
signal VN549_data_out : std_logic_vector(5 downto 0);
signal VN549_sign_out : std_logic_vector(5 downto 0);
signal VN550_data_out : std_logic_vector(5 downto 0);
signal VN550_sign_out : std_logic_vector(5 downto 0);
signal VN551_data_out : std_logic_vector(5 downto 0);
signal VN551_sign_out : std_logic_vector(5 downto 0);
signal VN552_data_out : std_logic_vector(5 downto 0);
signal VN552_sign_out : std_logic_vector(5 downto 0);
signal VN553_data_out : std_logic_vector(5 downto 0);
signal VN553_sign_out : std_logic_vector(5 downto 0);
signal VN554_data_out : std_logic_vector(5 downto 0);
signal VN554_sign_out : std_logic_vector(5 downto 0);
signal VN555_data_out : std_logic_vector(5 downto 0);
signal VN555_sign_out : std_logic_vector(5 downto 0);
signal VN556_data_out : std_logic_vector(5 downto 0);
signal VN556_sign_out : std_logic_vector(5 downto 0);
signal VN557_data_out : std_logic_vector(5 downto 0);
signal VN557_sign_out : std_logic_vector(5 downto 0);
signal VN558_data_out : std_logic_vector(5 downto 0);
signal VN558_sign_out : std_logic_vector(5 downto 0);
signal VN559_data_out : std_logic_vector(5 downto 0);
signal VN559_sign_out : std_logic_vector(5 downto 0);
signal VN560_data_out : std_logic_vector(5 downto 0);
signal VN560_sign_out : std_logic_vector(5 downto 0);
signal VN561_data_out : std_logic_vector(5 downto 0);
signal VN561_sign_out : std_logic_vector(5 downto 0);
signal VN562_data_out : std_logic_vector(5 downto 0);
signal VN562_sign_out : std_logic_vector(5 downto 0);
signal VN563_data_out : std_logic_vector(5 downto 0);
signal VN563_sign_out : std_logic_vector(5 downto 0);
signal VN564_data_out : std_logic_vector(5 downto 0);
signal VN564_sign_out : std_logic_vector(5 downto 0);
signal VN565_data_out : std_logic_vector(5 downto 0);
signal VN565_sign_out : std_logic_vector(5 downto 0);
signal VN566_data_out : std_logic_vector(5 downto 0);
signal VN566_sign_out : std_logic_vector(5 downto 0);
signal VN567_data_out : std_logic_vector(5 downto 0);
signal VN567_sign_out : std_logic_vector(5 downto 0);
signal VN568_data_out : std_logic_vector(5 downto 0);
signal VN568_sign_out : std_logic_vector(5 downto 0);
signal VN569_data_out : std_logic_vector(5 downto 0);
signal VN569_sign_out : std_logic_vector(5 downto 0);
signal VN570_data_out : std_logic_vector(5 downto 0);
signal VN570_sign_out : std_logic_vector(5 downto 0);
signal VN571_data_out : std_logic_vector(5 downto 0);
signal VN571_sign_out : std_logic_vector(5 downto 0);
signal VN572_data_out : std_logic_vector(5 downto 0);
signal VN572_sign_out : std_logic_vector(5 downto 0);
signal VN573_data_out : std_logic_vector(5 downto 0);
signal VN573_sign_out : std_logic_vector(5 downto 0);
signal VN574_data_out : std_logic_vector(5 downto 0);
signal VN574_sign_out : std_logic_vector(5 downto 0);
signal VN575_data_out : std_logic_vector(5 downto 0);
signal VN575_sign_out : std_logic_vector(5 downto 0);
signal VN576_data_out : std_logic_vector(5 downto 0);
signal VN576_sign_out : std_logic_vector(5 downto 0);
signal VN577_data_out : std_logic_vector(5 downto 0);
signal VN577_sign_out : std_logic_vector(5 downto 0);
signal VN578_data_out : std_logic_vector(5 downto 0);
signal VN578_sign_out : std_logic_vector(5 downto 0);
signal VN579_data_out : std_logic_vector(5 downto 0);
signal VN579_sign_out : std_logic_vector(5 downto 0);
signal VN580_data_out : std_logic_vector(5 downto 0);
signal VN580_sign_out : std_logic_vector(5 downto 0);
signal VN581_data_out : std_logic_vector(5 downto 0);
signal VN581_sign_out : std_logic_vector(5 downto 0);
signal VN582_data_out : std_logic_vector(5 downto 0);
signal VN582_sign_out : std_logic_vector(5 downto 0);
signal VN583_data_out : std_logic_vector(5 downto 0);
signal VN583_sign_out : std_logic_vector(5 downto 0);
signal VN584_data_out : std_logic_vector(5 downto 0);
signal VN584_sign_out : std_logic_vector(5 downto 0);
signal VN585_data_out : std_logic_vector(5 downto 0);
signal VN585_sign_out : std_logic_vector(5 downto 0);
signal VN586_data_out : std_logic_vector(5 downto 0);
signal VN586_sign_out : std_logic_vector(5 downto 0);
signal VN587_data_out : std_logic_vector(5 downto 0);
signal VN587_sign_out : std_logic_vector(5 downto 0);
signal VN588_data_out : std_logic_vector(5 downto 0);
signal VN588_sign_out : std_logic_vector(5 downto 0);
signal VN589_data_out : std_logic_vector(5 downto 0);
signal VN589_sign_out : std_logic_vector(5 downto 0);
signal VN590_data_out : std_logic_vector(5 downto 0);
signal VN590_sign_out : std_logic_vector(5 downto 0);
signal VN591_data_out : std_logic_vector(5 downto 0);
signal VN591_sign_out : std_logic_vector(5 downto 0);
signal VN592_data_out : std_logic_vector(5 downto 0);
signal VN592_sign_out : std_logic_vector(5 downto 0);
signal VN593_data_out : std_logic_vector(5 downto 0);
signal VN593_sign_out : std_logic_vector(5 downto 0);
signal VN594_data_out : std_logic_vector(5 downto 0);
signal VN594_sign_out : std_logic_vector(5 downto 0);
signal VN595_data_out : std_logic_vector(5 downto 0);
signal VN595_sign_out : std_logic_vector(5 downto 0);
signal VN596_data_out : std_logic_vector(5 downto 0);
signal VN596_sign_out : std_logic_vector(5 downto 0);
signal VN597_data_out : std_logic_vector(5 downto 0);
signal VN597_sign_out : std_logic_vector(5 downto 0);
signal VN598_data_out : std_logic_vector(5 downto 0);
signal VN598_sign_out : std_logic_vector(5 downto 0);
signal VN599_data_out : std_logic_vector(5 downto 0);
signal VN599_sign_out : std_logic_vector(5 downto 0);
signal VN600_data_out : std_logic_vector(5 downto 0);
signal VN600_sign_out : std_logic_vector(5 downto 0);
signal VN601_data_out : std_logic_vector(5 downto 0);
signal VN601_sign_out : std_logic_vector(5 downto 0);
signal VN602_data_out : std_logic_vector(5 downto 0);
signal VN602_sign_out : std_logic_vector(5 downto 0);
signal VN603_data_out : std_logic_vector(5 downto 0);
signal VN603_sign_out : std_logic_vector(5 downto 0);
signal VN604_data_out : std_logic_vector(5 downto 0);
signal VN604_sign_out : std_logic_vector(5 downto 0);
signal VN605_data_out : std_logic_vector(5 downto 0);
signal VN605_sign_out : std_logic_vector(5 downto 0);
signal VN606_data_out : std_logic_vector(5 downto 0);
signal VN606_sign_out : std_logic_vector(5 downto 0);
signal VN607_data_out : std_logic_vector(5 downto 0);
signal VN607_sign_out : std_logic_vector(5 downto 0);
signal VN608_data_out : std_logic_vector(5 downto 0);
signal VN608_sign_out : std_logic_vector(5 downto 0);
signal VN609_data_out : std_logic_vector(5 downto 0);
signal VN609_sign_out : std_logic_vector(5 downto 0);
signal VN610_data_out : std_logic_vector(5 downto 0);
signal VN610_sign_out : std_logic_vector(5 downto 0);
signal VN611_data_out : std_logic_vector(5 downto 0);
signal VN611_sign_out : std_logic_vector(5 downto 0);
signal VN612_data_out : std_logic_vector(5 downto 0);
signal VN612_sign_out : std_logic_vector(5 downto 0);
signal VN613_data_out : std_logic_vector(5 downto 0);
signal VN613_sign_out : std_logic_vector(5 downto 0);
signal VN614_data_out : std_logic_vector(5 downto 0);
signal VN614_sign_out : std_logic_vector(5 downto 0);
signal VN615_data_out : std_logic_vector(5 downto 0);
signal VN615_sign_out : std_logic_vector(5 downto 0);
signal VN616_data_out : std_logic_vector(5 downto 0);
signal VN616_sign_out : std_logic_vector(5 downto 0);
signal VN617_data_out : std_logic_vector(5 downto 0);
signal VN617_sign_out : std_logic_vector(5 downto 0);
signal VN618_data_out : std_logic_vector(5 downto 0);
signal VN618_sign_out : std_logic_vector(5 downto 0);
signal VN619_data_out : std_logic_vector(5 downto 0);
signal VN619_sign_out : std_logic_vector(5 downto 0);
signal VN620_data_out : std_logic_vector(5 downto 0);
signal VN620_sign_out : std_logic_vector(5 downto 0);
signal VN621_data_out : std_logic_vector(5 downto 0);
signal VN621_sign_out : std_logic_vector(5 downto 0);
signal VN622_data_out : std_logic_vector(5 downto 0);
signal VN622_sign_out : std_logic_vector(5 downto 0);
signal VN623_data_out : std_logic_vector(5 downto 0);
signal VN623_sign_out : std_logic_vector(5 downto 0);
signal VN624_data_out : std_logic_vector(5 downto 0);
signal VN624_sign_out : std_logic_vector(5 downto 0);
signal VN625_data_out : std_logic_vector(5 downto 0);
signal VN625_sign_out : std_logic_vector(5 downto 0);
signal VN626_data_out : std_logic_vector(5 downto 0);
signal VN626_sign_out : std_logic_vector(5 downto 0);
signal VN627_data_out : std_logic_vector(5 downto 0);
signal VN627_sign_out : std_logic_vector(5 downto 0);
signal VN628_data_out : std_logic_vector(5 downto 0);
signal VN628_sign_out : std_logic_vector(5 downto 0);
signal VN629_data_out : std_logic_vector(5 downto 0);
signal VN629_sign_out : std_logic_vector(5 downto 0);
signal VN630_data_out : std_logic_vector(5 downto 0);
signal VN630_sign_out : std_logic_vector(5 downto 0);
signal VN631_data_out : std_logic_vector(5 downto 0);
signal VN631_sign_out : std_logic_vector(5 downto 0);
signal VN632_data_out : std_logic_vector(5 downto 0);
signal VN632_sign_out : std_logic_vector(5 downto 0);
signal VN633_data_out : std_logic_vector(5 downto 0);
signal VN633_sign_out : std_logic_vector(5 downto 0);
signal VN634_data_out : std_logic_vector(5 downto 0);
signal VN634_sign_out : std_logic_vector(5 downto 0);
signal VN635_data_out : std_logic_vector(5 downto 0);
signal VN635_sign_out : std_logic_vector(5 downto 0);
signal VN636_data_out : std_logic_vector(5 downto 0);
signal VN636_sign_out : std_logic_vector(5 downto 0);
signal VN637_data_out : std_logic_vector(5 downto 0);
signal VN637_sign_out : std_logic_vector(5 downto 0);
signal VN638_data_out : std_logic_vector(5 downto 0);
signal VN638_sign_out : std_logic_vector(5 downto 0);
signal VN639_data_out : std_logic_vector(5 downto 0);
signal VN639_sign_out : std_logic_vector(5 downto 0);
signal VN640_data_out : std_logic_vector(5 downto 0);
signal VN640_sign_out : std_logic_vector(5 downto 0);
signal VN641_data_out : std_logic_vector(5 downto 0);
signal VN641_sign_out : std_logic_vector(5 downto 0);
signal VN642_data_out : std_logic_vector(5 downto 0);
signal VN642_sign_out : std_logic_vector(5 downto 0);
signal VN643_data_out : std_logic_vector(5 downto 0);
signal VN643_sign_out : std_logic_vector(5 downto 0);
signal VN644_data_out : std_logic_vector(5 downto 0);
signal VN644_sign_out : std_logic_vector(5 downto 0);
signal VN645_data_out : std_logic_vector(5 downto 0);
signal VN645_sign_out : std_logic_vector(5 downto 0);
signal VN646_data_out : std_logic_vector(5 downto 0);
signal VN646_sign_out : std_logic_vector(5 downto 0);
signal VN647_data_out : std_logic_vector(5 downto 0);
signal VN647_sign_out : std_logic_vector(5 downto 0);
signal VN648_data_out : std_logic_vector(5 downto 0);
signal VN648_sign_out : std_logic_vector(5 downto 0);
signal VN649_data_out : std_logic_vector(5 downto 0);
signal VN649_sign_out : std_logic_vector(5 downto 0);
signal VN650_data_out : std_logic_vector(5 downto 0);
signal VN650_sign_out : std_logic_vector(5 downto 0);
signal VN651_data_out : std_logic_vector(5 downto 0);
signal VN651_sign_out : std_logic_vector(5 downto 0);
signal VN652_data_out : std_logic_vector(5 downto 0);
signal VN652_sign_out : std_logic_vector(5 downto 0);
signal VN653_data_out : std_logic_vector(5 downto 0);
signal VN653_sign_out : std_logic_vector(5 downto 0);
signal VN654_data_out : std_logic_vector(5 downto 0);
signal VN654_sign_out : std_logic_vector(5 downto 0);
signal VN655_data_out : std_logic_vector(5 downto 0);
signal VN655_sign_out : std_logic_vector(5 downto 0);
signal VN656_data_out : std_logic_vector(5 downto 0);
signal VN656_sign_out : std_logic_vector(5 downto 0);
signal VN657_data_out : std_logic_vector(5 downto 0);
signal VN657_sign_out : std_logic_vector(5 downto 0);
signal VN658_data_out : std_logic_vector(5 downto 0);
signal VN658_sign_out : std_logic_vector(5 downto 0);
signal VN659_data_out : std_logic_vector(5 downto 0);
signal VN659_sign_out : std_logic_vector(5 downto 0);
signal VN660_data_out : std_logic_vector(5 downto 0);
signal VN660_sign_out : std_logic_vector(5 downto 0);
signal VN661_data_out : std_logic_vector(5 downto 0);
signal VN661_sign_out : std_logic_vector(5 downto 0);
signal VN662_data_out : std_logic_vector(5 downto 0);
signal VN662_sign_out : std_logic_vector(5 downto 0);
signal VN663_data_out : std_logic_vector(5 downto 0);
signal VN663_sign_out : std_logic_vector(5 downto 0);
signal VN664_data_out : std_logic_vector(5 downto 0);
signal VN664_sign_out : std_logic_vector(5 downto 0);
signal VN665_data_out : std_logic_vector(5 downto 0);
signal VN665_sign_out : std_logic_vector(5 downto 0);
signal VN666_data_out : std_logic_vector(5 downto 0);
signal VN666_sign_out : std_logic_vector(5 downto 0);
signal VN667_data_out : std_logic_vector(5 downto 0);
signal VN667_sign_out : std_logic_vector(5 downto 0);
signal VN668_data_out : std_logic_vector(5 downto 0);
signal VN668_sign_out : std_logic_vector(5 downto 0);
signal VN669_data_out : std_logic_vector(5 downto 0);
signal VN669_sign_out : std_logic_vector(5 downto 0);
signal VN670_data_out : std_logic_vector(5 downto 0);
signal VN670_sign_out : std_logic_vector(5 downto 0);
signal VN671_data_out : std_logic_vector(5 downto 0);
signal VN671_sign_out : std_logic_vector(5 downto 0);
signal VN672_data_out : std_logic_vector(5 downto 0);
signal VN672_sign_out : std_logic_vector(5 downto 0);
signal VN673_data_out : std_logic_vector(5 downto 0);
signal VN673_sign_out : std_logic_vector(5 downto 0);
signal VN674_data_out : std_logic_vector(5 downto 0);
signal VN674_sign_out : std_logic_vector(5 downto 0);
signal VN675_data_out : std_logic_vector(5 downto 0);
signal VN675_sign_out : std_logic_vector(5 downto 0);
signal VN676_data_out : std_logic_vector(5 downto 0);
signal VN676_sign_out : std_logic_vector(5 downto 0);
signal VN677_data_out : std_logic_vector(5 downto 0);
signal VN677_sign_out : std_logic_vector(5 downto 0);
signal VN678_data_out : std_logic_vector(5 downto 0);
signal VN678_sign_out : std_logic_vector(5 downto 0);
signal VN679_data_out : std_logic_vector(5 downto 0);
signal VN679_sign_out : std_logic_vector(5 downto 0);
signal VN680_data_out : std_logic_vector(5 downto 0);
signal VN680_sign_out : std_logic_vector(5 downto 0);
signal VN681_data_out : std_logic_vector(5 downto 0);
signal VN681_sign_out : std_logic_vector(5 downto 0);
signal VN682_data_out : std_logic_vector(5 downto 0);
signal VN682_sign_out : std_logic_vector(5 downto 0);
signal VN683_data_out : std_logic_vector(5 downto 0);
signal VN683_sign_out : std_logic_vector(5 downto 0);
signal VN684_data_out : std_logic_vector(5 downto 0);
signal VN684_sign_out : std_logic_vector(5 downto 0);
signal VN685_data_out : std_logic_vector(5 downto 0);
signal VN685_sign_out : std_logic_vector(5 downto 0);
signal VN686_data_out : std_logic_vector(5 downto 0);
signal VN686_sign_out : std_logic_vector(5 downto 0);
signal VN687_data_out : std_logic_vector(5 downto 0);
signal VN687_sign_out : std_logic_vector(5 downto 0);
signal VN688_data_out : std_logic_vector(5 downto 0);
signal VN688_sign_out : std_logic_vector(5 downto 0);
signal VN689_data_out : std_logic_vector(5 downto 0);
signal VN689_sign_out : std_logic_vector(5 downto 0);
signal VN690_data_out : std_logic_vector(5 downto 0);
signal VN690_sign_out : std_logic_vector(5 downto 0);
signal VN691_data_out : std_logic_vector(5 downto 0);
signal VN691_sign_out : std_logic_vector(5 downto 0);
signal VN692_data_out : std_logic_vector(5 downto 0);
signal VN692_sign_out : std_logic_vector(5 downto 0);
signal VN693_data_out : std_logic_vector(5 downto 0);
signal VN693_sign_out : std_logic_vector(5 downto 0);
signal VN694_data_out : std_logic_vector(5 downto 0);
signal VN694_sign_out : std_logic_vector(5 downto 0);
signal VN695_data_out : std_logic_vector(5 downto 0);
signal VN695_sign_out : std_logic_vector(5 downto 0);
signal VN696_data_out : std_logic_vector(5 downto 0);
signal VN696_sign_out : std_logic_vector(5 downto 0);
signal VN697_data_out : std_logic_vector(5 downto 0);
signal VN697_sign_out : std_logic_vector(5 downto 0);
signal VN698_data_out : std_logic_vector(5 downto 0);
signal VN698_sign_out : std_logic_vector(5 downto 0);
signal VN699_data_out : std_logic_vector(5 downto 0);
signal VN699_sign_out : std_logic_vector(5 downto 0);
signal VN700_data_out : std_logic_vector(5 downto 0);
signal VN700_sign_out : std_logic_vector(5 downto 0);
signal VN701_data_out : std_logic_vector(5 downto 0);
signal VN701_sign_out : std_logic_vector(5 downto 0);
signal VN702_data_out : std_logic_vector(5 downto 0);
signal VN702_sign_out : std_logic_vector(5 downto 0);
signal VN703_data_out : std_logic_vector(5 downto 0);
signal VN703_sign_out : std_logic_vector(5 downto 0);
signal VN704_data_out : std_logic_vector(5 downto 0);
signal VN704_sign_out : std_logic_vector(5 downto 0);
signal VN705_data_out : std_logic_vector(5 downto 0);
signal VN705_sign_out : std_logic_vector(5 downto 0);
signal VN706_data_out : std_logic_vector(5 downto 0);
signal VN706_sign_out : std_logic_vector(5 downto 0);
signal VN707_data_out : std_logic_vector(5 downto 0);
signal VN707_sign_out : std_logic_vector(5 downto 0);
signal VN708_data_out : std_logic_vector(5 downto 0);
signal VN708_sign_out : std_logic_vector(5 downto 0);
signal VN709_data_out : std_logic_vector(5 downto 0);
signal VN709_sign_out : std_logic_vector(5 downto 0);
signal VN710_data_out : std_logic_vector(5 downto 0);
signal VN710_sign_out : std_logic_vector(5 downto 0);
signal VN711_data_out : std_logic_vector(5 downto 0);
signal VN711_sign_out : std_logic_vector(5 downto 0);
signal VN712_data_out : std_logic_vector(5 downto 0);
signal VN712_sign_out : std_logic_vector(5 downto 0);
signal VN713_data_out : std_logic_vector(5 downto 0);
signal VN713_sign_out : std_logic_vector(5 downto 0);
signal VN714_data_out : std_logic_vector(5 downto 0);
signal VN714_sign_out : std_logic_vector(5 downto 0);
signal VN715_data_out : std_logic_vector(5 downto 0);
signal VN715_sign_out : std_logic_vector(5 downto 0);
signal VN716_data_out : std_logic_vector(5 downto 0);
signal VN716_sign_out : std_logic_vector(5 downto 0);
signal VN717_data_out : std_logic_vector(5 downto 0);
signal VN717_sign_out : std_logic_vector(5 downto 0);
signal VN718_data_out : std_logic_vector(5 downto 0);
signal VN718_sign_out : std_logic_vector(5 downto 0);
signal VN719_data_out : std_logic_vector(5 downto 0);
signal VN719_sign_out : std_logic_vector(5 downto 0);
signal VN720_data_out : std_logic_vector(5 downto 0);
signal VN720_sign_out : std_logic_vector(5 downto 0);
signal VN721_data_out : std_logic_vector(5 downto 0);
signal VN721_sign_out : std_logic_vector(5 downto 0);
signal VN722_data_out : std_logic_vector(5 downto 0);
signal VN722_sign_out : std_logic_vector(5 downto 0);
signal VN723_data_out : std_logic_vector(5 downto 0);
signal VN723_sign_out : std_logic_vector(5 downto 0);
signal VN724_data_out : std_logic_vector(5 downto 0);
signal VN724_sign_out : std_logic_vector(5 downto 0);
signal VN725_data_out : std_logic_vector(5 downto 0);
signal VN725_sign_out : std_logic_vector(5 downto 0);
signal VN726_data_out : std_logic_vector(5 downto 0);
signal VN726_sign_out : std_logic_vector(5 downto 0);
signal VN727_data_out : std_logic_vector(5 downto 0);
signal VN727_sign_out : std_logic_vector(5 downto 0);
signal VN728_data_out : std_logic_vector(5 downto 0);
signal VN728_sign_out : std_logic_vector(5 downto 0);
signal VN729_data_out : std_logic_vector(5 downto 0);
signal VN729_sign_out : std_logic_vector(5 downto 0);
signal VN730_data_out : std_logic_vector(5 downto 0);
signal VN730_sign_out : std_logic_vector(5 downto 0);
signal VN731_data_out : std_logic_vector(5 downto 0);
signal VN731_sign_out : std_logic_vector(5 downto 0);
signal VN732_data_out : std_logic_vector(5 downto 0);
signal VN732_sign_out : std_logic_vector(5 downto 0);
signal VN733_data_out : std_logic_vector(5 downto 0);
signal VN733_sign_out : std_logic_vector(5 downto 0);
signal VN734_data_out : std_logic_vector(5 downto 0);
signal VN734_sign_out : std_logic_vector(5 downto 0);
signal VN735_data_out : std_logic_vector(5 downto 0);
signal VN735_sign_out : std_logic_vector(5 downto 0);
signal VN736_data_out : std_logic_vector(5 downto 0);
signal VN736_sign_out : std_logic_vector(5 downto 0);
signal VN737_data_out : std_logic_vector(5 downto 0);
signal VN737_sign_out : std_logic_vector(5 downto 0);
signal VN738_data_out : std_logic_vector(5 downto 0);
signal VN738_sign_out : std_logic_vector(5 downto 0);
signal VN739_data_out : std_logic_vector(5 downto 0);
signal VN739_sign_out : std_logic_vector(5 downto 0);
signal VN740_data_out : std_logic_vector(5 downto 0);
signal VN740_sign_out : std_logic_vector(5 downto 0);
signal VN741_data_out : std_logic_vector(5 downto 0);
signal VN741_sign_out : std_logic_vector(5 downto 0);
signal VN742_data_out : std_logic_vector(5 downto 0);
signal VN742_sign_out : std_logic_vector(5 downto 0);
signal VN743_data_out : std_logic_vector(5 downto 0);
signal VN743_sign_out : std_logic_vector(5 downto 0);
signal VN744_data_out : std_logic_vector(5 downto 0);
signal VN744_sign_out : std_logic_vector(5 downto 0);
signal VN745_data_out : std_logic_vector(5 downto 0);
signal VN745_sign_out : std_logic_vector(5 downto 0);
signal VN746_data_out : std_logic_vector(5 downto 0);
signal VN746_sign_out : std_logic_vector(5 downto 0);
signal VN747_data_out : std_logic_vector(5 downto 0);
signal VN747_sign_out : std_logic_vector(5 downto 0);
signal VN748_data_out : std_logic_vector(5 downto 0);
signal VN748_sign_out : std_logic_vector(5 downto 0);
signal VN749_data_out : std_logic_vector(5 downto 0);
signal VN749_sign_out : std_logic_vector(5 downto 0);
signal VN750_data_out : std_logic_vector(5 downto 0);
signal VN750_sign_out : std_logic_vector(5 downto 0);
signal VN751_data_out : std_logic_vector(5 downto 0);
signal VN751_sign_out : std_logic_vector(5 downto 0);
signal VN752_data_out : std_logic_vector(5 downto 0);
signal VN752_sign_out : std_logic_vector(5 downto 0);
signal VN753_data_out : std_logic_vector(5 downto 0);
signal VN753_sign_out : std_logic_vector(5 downto 0);
signal VN754_data_out : std_logic_vector(5 downto 0);
signal VN754_sign_out : std_logic_vector(5 downto 0);
signal VN755_data_out : std_logic_vector(5 downto 0);
signal VN755_sign_out : std_logic_vector(5 downto 0);
signal VN756_data_out : std_logic_vector(5 downto 0);
signal VN756_sign_out : std_logic_vector(5 downto 0);
signal VN757_data_out : std_logic_vector(5 downto 0);
signal VN757_sign_out : std_logic_vector(5 downto 0);
signal VN758_data_out : std_logic_vector(5 downto 0);
signal VN758_sign_out : std_logic_vector(5 downto 0);
signal VN759_data_out : std_logic_vector(5 downto 0);
signal VN759_sign_out : std_logic_vector(5 downto 0);
signal VN760_data_out : std_logic_vector(5 downto 0);
signal VN760_sign_out : std_logic_vector(5 downto 0);
signal VN761_data_out : std_logic_vector(5 downto 0);
signal VN761_sign_out : std_logic_vector(5 downto 0);
signal VN762_data_out : std_logic_vector(5 downto 0);
signal VN762_sign_out : std_logic_vector(5 downto 0);
signal VN763_data_out : std_logic_vector(5 downto 0);
signal VN763_sign_out : std_logic_vector(5 downto 0);
signal VN764_data_out : std_logic_vector(5 downto 0);
signal VN764_sign_out : std_logic_vector(5 downto 0);
signal VN765_data_out : std_logic_vector(5 downto 0);
signal VN765_sign_out : std_logic_vector(5 downto 0);
signal VN766_data_out : std_logic_vector(5 downto 0);
signal VN766_sign_out : std_logic_vector(5 downto 0);
signal VN767_data_out : std_logic_vector(5 downto 0);
signal VN767_sign_out : std_logic_vector(5 downto 0);
signal VN768_data_out : std_logic_vector(5 downto 0);
signal VN768_sign_out : std_logic_vector(5 downto 0);
signal VN769_data_out : std_logic_vector(5 downto 0);
signal VN769_sign_out : std_logic_vector(5 downto 0);
signal VN770_data_out : std_logic_vector(5 downto 0);
signal VN770_sign_out : std_logic_vector(5 downto 0);
signal VN771_data_out : std_logic_vector(5 downto 0);
signal VN771_sign_out : std_logic_vector(5 downto 0);
signal VN772_data_out : std_logic_vector(5 downto 0);
signal VN772_sign_out : std_logic_vector(5 downto 0);
signal VN773_data_out : std_logic_vector(5 downto 0);
signal VN773_sign_out : std_logic_vector(5 downto 0);
signal VN774_data_out : std_logic_vector(5 downto 0);
signal VN774_sign_out : std_logic_vector(5 downto 0);
signal VN775_data_out : std_logic_vector(5 downto 0);
signal VN775_sign_out : std_logic_vector(5 downto 0);
signal VN776_data_out : std_logic_vector(5 downto 0);
signal VN776_sign_out : std_logic_vector(5 downto 0);
signal VN777_data_out : std_logic_vector(5 downto 0);
signal VN777_sign_out : std_logic_vector(5 downto 0);
signal VN778_data_out : std_logic_vector(5 downto 0);
signal VN778_sign_out : std_logic_vector(5 downto 0);
signal VN779_data_out : std_logic_vector(5 downto 0);
signal VN779_sign_out : std_logic_vector(5 downto 0);
signal VN780_data_out : std_logic_vector(5 downto 0);
signal VN780_sign_out : std_logic_vector(5 downto 0);
signal VN781_data_out : std_logic_vector(5 downto 0);
signal VN781_sign_out : std_logic_vector(5 downto 0);
signal VN782_data_out : std_logic_vector(5 downto 0);
signal VN782_sign_out : std_logic_vector(5 downto 0);
signal VN783_data_out : std_logic_vector(5 downto 0);
signal VN783_sign_out : std_logic_vector(5 downto 0);
signal VN784_data_out : std_logic_vector(5 downto 0);
signal VN784_sign_out : std_logic_vector(5 downto 0);
signal VN785_data_out : std_logic_vector(5 downto 0);
signal VN785_sign_out : std_logic_vector(5 downto 0);
signal VN786_data_out : std_logic_vector(5 downto 0);
signal VN786_sign_out : std_logic_vector(5 downto 0);
signal VN787_data_out : std_logic_vector(5 downto 0);
signal VN787_sign_out : std_logic_vector(5 downto 0);
signal VN788_data_out : std_logic_vector(5 downto 0);
signal VN788_sign_out : std_logic_vector(5 downto 0);
signal VN789_data_out : std_logic_vector(5 downto 0);
signal VN789_sign_out : std_logic_vector(5 downto 0);
signal VN790_data_out : std_logic_vector(5 downto 0);
signal VN790_sign_out : std_logic_vector(5 downto 0);
signal VN791_data_out : std_logic_vector(5 downto 0);
signal VN791_sign_out : std_logic_vector(5 downto 0);
signal VN792_data_out : std_logic_vector(5 downto 0);
signal VN792_sign_out : std_logic_vector(5 downto 0);
signal VN793_data_out : std_logic_vector(5 downto 0);
signal VN793_sign_out : std_logic_vector(5 downto 0);
signal VN794_data_out : std_logic_vector(5 downto 0);
signal VN794_sign_out : std_logic_vector(5 downto 0);
signal VN795_data_out : std_logic_vector(5 downto 0);
signal VN795_sign_out : std_logic_vector(5 downto 0);
signal VN796_data_out : std_logic_vector(5 downto 0);
signal VN796_sign_out : std_logic_vector(5 downto 0);
signal VN797_data_out : std_logic_vector(5 downto 0);
signal VN797_sign_out : std_logic_vector(5 downto 0);
signal VN798_data_out : std_logic_vector(5 downto 0);
signal VN798_sign_out : std_logic_vector(5 downto 0);
signal VN799_data_out : std_logic_vector(5 downto 0);
signal VN799_sign_out : std_logic_vector(5 downto 0);
signal VN800_data_out : std_logic_vector(5 downto 0);
signal VN800_sign_out : std_logic_vector(5 downto 0);
signal VN801_data_out : std_logic_vector(5 downto 0);
signal VN801_sign_out : std_logic_vector(5 downto 0);
signal VN802_data_out : std_logic_vector(5 downto 0);
signal VN802_sign_out : std_logic_vector(5 downto 0);
signal VN803_data_out : std_logic_vector(5 downto 0);
signal VN803_sign_out : std_logic_vector(5 downto 0);
signal VN804_data_out : std_logic_vector(5 downto 0);
signal VN804_sign_out : std_logic_vector(5 downto 0);
signal VN805_data_out : std_logic_vector(5 downto 0);
signal VN805_sign_out : std_logic_vector(5 downto 0);
signal VN806_data_out : std_logic_vector(5 downto 0);
signal VN806_sign_out : std_logic_vector(5 downto 0);
signal VN807_data_out : std_logic_vector(5 downto 0);
signal VN807_sign_out : std_logic_vector(5 downto 0);
signal VN808_data_out : std_logic_vector(5 downto 0);
signal VN808_sign_out : std_logic_vector(5 downto 0);
signal VN809_data_out : std_logic_vector(5 downto 0);
signal VN809_sign_out : std_logic_vector(5 downto 0);
signal VN810_data_out : std_logic_vector(5 downto 0);
signal VN810_sign_out : std_logic_vector(5 downto 0);
signal VN811_data_out : std_logic_vector(5 downto 0);
signal VN811_sign_out : std_logic_vector(5 downto 0);
signal VN812_data_out : std_logic_vector(5 downto 0);
signal VN812_sign_out : std_logic_vector(5 downto 0);
signal VN813_data_out : std_logic_vector(5 downto 0);
signal VN813_sign_out : std_logic_vector(5 downto 0);
signal VN814_data_out : std_logic_vector(5 downto 0);
signal VN814_sign_out : std_logic_vector(5 downto 0);
signal VN815_data_out : std_logic_vector(5 downto 0);
signal VN815_sign_out : std_logic_vector(5 downto 0);
signal VN816_data_out : std_logic_vector(5 downto 0);
signal VN816_sign_out : std_logic_vector(5 downto 0);
signal VN817_data_out : std_logic_vector(5 downto 0);
signal VN817_sign_out : std_logic_vector(5 downto 0);
signal VN818_data_out : std_logic_vector(5 downto 0);
signal VN818_sign_out : std_logic_vector(5 downto 0);
signal VN819_data_out : std_logic_vector(5 downto 0);
signal VN819_sign_out : std_logic_vector(5 downto 0);
signal VN820_data_out : std_logic_vector(5 downto 0);
signal VN820_sign_out : std_logic_vector(5 downto 0);
signal VN821_data_out : std_logic_vector(5 downto 0);
signal VN821_sign_out : std_logic_vector(5 downto 0);
signal VN822_data_out : std_logic_vector(5 downto 0);
signal VN822_sign_out : std_logic_vector(5 downto 0);
signal VN823_data_out : std_logic_vector(5 downto 0);
signal VN823_sign_out : std_logic_vector(5 downto 0);
signal VN824_data_out : std_logic_vector(5 downto 0);
signal VN824_sign_out : std_logic_vector(5 downto 0);
signal VN825_data_out : std_logic_vector(5 downto 0);
signal VN825_sign_out : std_logic_vector(5 downto 0);
signal VN826_data_out : std_logic_vector(5 downto 0);
signal VN826_sign_out : std_logic_vector(5 downto 0);
signal VN827_data_out : std_logic_vector(5 downto 0);
signal VN827_sign_out : std_logic_vector(5 downto 0);
signal VN828_data_out : std_logic_vector(5 downto 0);
signal VN828_sign_out : std_logic_vector(5 downto 0);
signal VN829_data_out : std_logic_vector(5 downto 0);
signal VN829_sign_out : std_logic_vector(5 downto 0);
signal VN830_data_out : std_logic_vector(5 downto 0);
signal VN830_sign_out : std_logic_vector(5 downto 0);
signal VN831_data_out : std_logic_vector(5 downto 0);
signal VN831_sign_out : std_logic_vector(5 downto 0);
signal VN832_data_out : std_logic_vector(5 downto 0);
signal VN832_sign_out : std_logic_vector(5 downto 0);
signal VN833_data_out : std_logic_vector(5 downto 0);
signal VN833_sign_out : std_logic_vector(5 downto 0);
signal VN834_data_out : std_logic_vector(5 downto 0);
signal VN834_sign_out : std_logic_vector(5 downto 0);
signal VN835_data_out : std_logic_vector(5 downto 0);
signal VN835_sign_out : std_logic_vector(5 downto 0);
signal VN836_data_out : std_logic_vector(5 downto 0);
signal VN836_sign_out : std_logic_vector(5 downto 0);
signal VN837_data_out : std_logic_vector(5 downto 0);
signal VN837_sign_out : std_logic_vector(5 downto 0);
signal VN838_data_out : std_logic_vector(5 downto 0);
signal VN838_sign_out : std_logic_vector(5 downto 0);
signal VN839_data_out : std_logic_vector(5 downto 0);
signal VN839_sign_out : std_logic_vector(5 downto 0);
signal VN840_data_out : std_logic_vector(5 downto 0);
signal VN840_sign_out : std_logic_vector(5 downto 0);
signal VN841_data_out : std_logic_vector(5 downto 0);
signal VN841_sign_out : std_logic_vector(5 downto 0);
signal VN842_data_out : std_logic_vector(5 downto 0);
signal VN842_sign_out : std_logic_vector(5 downto 0);
signal VN843_data_out : std_logic_vector(5 downto 0);
signal VN843_sign_out : std_logic_vector(5 downto 0);
signal VN844_data_out : std_logic_vector(5 downto 0);
signal VN844_sign_out : std_logic_vector(5 downto 0);
signal VN845_data_out : std_logic_vector(5 downto 0);
signal VN845_sign_out : std_logic_vector(5 downto 0);
signal VN846_data_out : std_logic_vector(5 downto 0);
signal VN846_sign_out : std_logic_vector(5 downto 0);
signal VN847_data_out : std_logic_vector(5 downto 0);
signal VN847_sign_out : std_logic_vector(5 downto 0);
signal VN848_data_out : std_logic_vector(5 downto 0);
signal VN848_sign_out : std_logic_vector(5 downto 0);
signal VN849_data_out : std_logic_vector(5 downto 0);
signal VN849_sign_out : std_logic_vector(5 downto 0);
signal VN850_data_out : std_logic_vector(5 downto 0);
signal VN850_sign_out : std_logic_vector(5 downto 0);
signal VN851_data_out : std_logic_vector(5 downto 0);
signal VN851_sign_out : std_logic_vector(5 downto 0);
signal VN852_data_out : std_logic_vector(5 downto 0);
signal VN852_sign_out : std_logic_vector(5 downto 0);
signal VN853_data_out : std_logic_vector(5 downto 0);
signal VN853_sign_out : std_logic_vector(5 downto 0);
signal VN854_data_out : std_logic_vector(5 downto 0);
signal VN854_sign_out : std_logic_vector(5 downto 0);
signal VN855_data_out : std_logic_vector(5 downto 0);
signal VN855_sign_out : std_logic_vector(5 downto 0);
signal VN856_data_out : std_logic_vector(5 downto 0);
signal VN856_sign_out : std_logic_vector(5 downto 0);
signal VN857_data_out : std_logic_vector(5 downto 0);
signal VN857_sign_out : std_logic_vector(5 downto 0);
signal VN858_data_out : std_logic_vector(5 downto 0);
signal VN858_sign_out : std_logic_vector(5 downto 0);
signal VN859_data_out : std_logic_vector(5 downto 0);
signal VN859_sign_out : std_logic_vector(5 downto 0);
signal VN860_data_out : std_logic_vector(5 downto 0);
signal VN860_sign_out : std_logic_vector(5 downto 0);
signal VN861_data_out : std_logic_vector(5 downto 0);
signal VN861_sign_out : std_logic_vector(5 downto 0);
signal VN862_data_out : std_logic_vector(5 downto 0);
signal VN862_sign_out : std_logic_vector(5 downto 0);
signal VN863_data_out : std_logic_vector(5 downto 0);
signal VN863_sign_out : std_logic_vector(5 downto 0);
signal VN864_data_out : std_logic_vector(5 downto 0);
signal VN864_sign_out : std_logic_vector(5 downto 0);
signal VN865_data_out : std_logic_vector(5 downto 0);
signal VN865_sign_out : std_logic_vector(5 downto 0);
signal VN866_data_out : std_logic_vector(5 downto 0);
signal VN866_sign_out : std_logic_vector(5 downto 0);
signal VN867_data_out : std_logic_vector(5 downto 0);
signal VN867_sign_out : std_logic_vector(5 downto 0);
signal VN868_data_out : std_logic_vector(5 downto 0);
signal VN868_sign_out : std_logic_vector(5 downto 0);
signal VN869_data_out : std_logic_vector(5 downto 0);
signal VN869_sign_out : std_logic_vector(5 downto 0);
signal VN870_data_out : std_logic_vector(5 downto 0);
signal VN870_sign_out : std_logic_vector(5 downto 0);
signal VN871_data_out : std_logic_vector(5 downto 0);
signal VN871_sign_out : std_logic_vector(5 downto 0);
signal VN872_data_out : std_logic_vector(5 downto 0);
signal VN872_sign_out : std_logic_vector(5 downto 0);
signal VN873_data_out : std_logic_vector(5 downto 0);
signal VN873_sign_out : std_logic_vector(5 downto 0);
signal VN874_data_out : std_logic_vector(5 downto 0);
signal VN874_sign_out : std_logic_vector(5 downto 0);
signal VN875_data_out : std_logic_vector(5 downto 0);
signal VN875_sign_out : std_logic_vector(5 downto 0);
signal VN876_data_out : std_logic_vector(5 downto 0);
signal VN876_sign_out : std_logic_vector(5 downto 0);
signal VN877_data_out : std_logic_vector(5 downto 0);
signal VN877_sign_out : std_logic_vector(5 downto 0);
signal VN878_data_out : std_logic_vector(5 downto 0);
signal VN878_sign_out : std_logic_vector(5 downto 0);
signal VN879_data_out : std_logic_vector(5 downto 0);
signal VN879_sign_out : std_logic_vector(5 downto 0);
signal VN880_data_out : std_logic_vector(5 downto 0);
signal VN880_sign_out : std_logic_vector(5 downto 0);
signal VN881_data_out : std_logic_vector(5 downto 0);
signal VN881_sign_out : std_logic_vector(5 downto 0);
signal VN882_data_out : std_logic_vector(5 downto 0);
signal VN882_sign_out : std_logic_vector(5 downto 0);
signal VN883_data_out : std_logic_vector(5 downto 0);
signal VN883_sign_out : std_logic_vector(5 downto 0);
signal VN884_data_out : std_logic_vector(5 downto 0);
signal VN884_sign_out : std_logic_vector(5 downto 0);
signal VN885_data_out : std_logic_vector(5 downto 0);
signal VN885_sign_out : std_logic_vector(5 downto 0);
signal VN886_data_out : std_logic_vector(5 downto 0);
signal VN886_sign_out : std_logic_vector(5 downto 0);
signal VN887_data_out : std_logic_vector(5 downto 0);
signal VN887_sign_out : std_logic_vector(5 downto 0);
signal VN888_data_out : std_logic_vector(5 downto 0);
signal VN888_sign_out : std_logic_vector(5 downto 0);
signal VN889_data_out : std_logic_vector(5 downto 0);
signal VN889_sign_out : std_logic_vector(5 downto 0);
signal VN890_data_out : std_logic_vector(5 downto 0);
signal VN890_sign_out : std_logic_vector(5 downto 0);
signal VN891_data_out : std_logic_vector(5 downto 0);
signal VN891_sign_out : std_logic_vector(5 downto 0);
signal VN892_data_out : std_logic_vector(5 downto 0);
signal VN892_sign_out : std_logic_vector(5 downto 0);
signal VN893_data_out : std_logic_vector(5 downto 0);
signal VN893_sign_out : std_logic_vector(5 downto 0);
signal VN894_data_out : std_logic_vector(5 downto 0);
signal VN894_sign_out : std_logic_vector(5 downto 0);
signal VN895_data_out : std_logic_vector(5 downto 0);
signal VN895_sign_out : std_logic_vector(5 downto 0);
signal VN896_data_out : std_logic_vector(5 downto 0);
signal VN896_sign_out : std_logic_vector(5 downto 0);
signal VN897_data_out : std_logic_vector(5 downto 0);
signal VN897_sign_out : std_logic_vector(5 downto 0);
signal VN898_data_out : std_logic_vector(5 downto 0);
signal VN898_sign_out : std_logic_vector(5 downto 0);
signal VN899_data_out : std_logic_vector(5 downto 0);
signal VN899_sign_out : std_logic_vector(5 downto 0);
signal VN900_data_out : std_logic_vector(5 downto 0);
signal VN900_sign_out : std_logic_vector(5 downto 0);
signal VN901_data_out : std_logic_vector(5 downto 0);
signal VN901_sign_out : std_logic_vector(5 downto 0);
signal VN902_data_out : std_logic_vector(5 downto 0);
signal VN902_sign_out : std_logic_vector(5 downto 0);
signal VN903_data_out : std_logic_vector(5 downto 0);
signal VN903_sign_out : std_logic_vector(5 downto 0);
signal VN904_data_out : std_logic_vector(5 downto 0);
signal VN904_sign_out : std_logic_vector(5 downto 0);
signal VN905_data_out : std_logic_vector(5 downto 0);
signal VN905_sign_out : std_logic_vector(5 downto 0);
signal VN906_data_out : std_logic_vector(5 downto 0);
signal VN906_sign_out : std_logic_vector(5 downto 0);
signal VN907_data_out : std_logic_vector(5 downto 0);
signal VN907_sign_out : std_logic_vector(5 downto 0);
signal VN908_data_out : std_logic_vector(5 downto 0);
signal VN908_sign_out : std_logic_vector(5 downto 0);
signal VN909_data_out : std_logic_vector(5 downto 0);
signal VN909_sign_out : std_logic_vector(5 downto 0);
signal VN910_data_out : std_logic_vector(5 downto 0);
signal VN910_sign_out : std_logic_vector(5 downto 0);
signal VN911_data_out : std_logic_vector(5 downto 0);
signal VN911_sign_out : std_logic_vector(5 downto 0);
signal VN912_data_out : std_logic_vector(5 downto 0);
signal VN912_sign_out : std_logic_vector(5 downto 0);
signal VN913_data_out : std_logic_vector(5 downto 0);
signal VN913_sign_out : std_logic_vector(5 downto 0);
signal VN914_data_out : std_logic_vector(5 downto 0);
signal VN914_sign_out : std_logic_vector(5 downto 0);
signal VN915_data_out : std_logic_vector(5 downto 0);
signal VN915_sign_out : std_logic_vector(5 downto 0);
signal VN916_data_out : std_logic_vector(5 downto 0);
signal VN916_sign_out : std_logic_vector(5 downto 0);
signal VN917_data_out : std_logic_vector(5 downto 0);
signal VN917_sign_out : std_logic_vector(5 downto 0);
signal VN918_data_out : std_logic_vector(5 downto 0);
signal VN918_sign_out : std_logic_vector(5 downto 0);
signal VN919_data_out : std_logic_vector(5 downto 0);
signal VN919_sign_out : std_logic_vector(5 downto 0);
signal VN920_data_out : std_logic_vector(5 downto 0);
signal VN920_sign_out : std_logic_vector(5 downto 0);
signal VN921_data_out : std_logic_vector(5 downto 0);
signal VN921_sign_out : std_logic_vector(5 downto 0);
signal VN922_data_out : std_logic_vector(5 downto 0);
signal VN922_sign_out : std_logic_vector(5 downto 0);
signal VN923_data_out : std_logic_vector(5 downto 0);
signal VN923_sign_out : std_logic_vector(5 downto 0);
signal VN924_data_out : std_logic_vector(5 downto 0);
signal VN924_sign_out : std_logic_vector(5 downto 0);
signal VN925_data_out : std_logic_vector(5 downto 0);
signal VN925_sign_out : std_logic_vector(5 downto 0);
signal VN926_data_out : std_logic_vector(5 downto 0);
signal VN926_sign_out : std_logic_vector(5 downto 0);
signal VN927_data_out : std_logic_vector(5 downto 0);
signal VN927_sign_out : std_logic_vector(5 downto 0);
signal VN928_data_out : std_logic_vector(5 downto 0);
signal VN928_sign_out : std_logic_vector(5 downto 0);
signal VN929_data_out : std_logic_vector(5 downto 0);
signal VN929_sign_out : std_logic_vector(5 downto 0);
signal VN930_data_out : std_logic_vector(5 downto 0);
signal VN930_sign_out : std_logic_vector(5 downto 0);
signal VN931_data_out : std_logic_vector(5 downto 0);
signal VN931_sign_out : std_logic_vector(5 downto 0);
signal VN932_data_out : std_logic_vector(5 downto 0);
signal VN932_sign_out : std_logic_vector(5 downto 0);
signal VN933_data_out : std_logic_vector(5 downto 0);
signal VN933_sign_out : std_logic_vector(5 downto 0);
signal VN934_data_out : std_logic_vector(5 downto 0);
signal VN934_sign_out : std_logic_vector(5 downto 0);
signal VN935_data_out : std_logic_vector(5 downto 0);
signal VN935_sign_out : std_logic_vector(5 downto 0);
signal VN936_data_out : std_logic_vector(5 downto 0);
signal VN936_sign_out : std_logic_vector(5 downto 0);
signal VN937_data_out : std_logic_vector(5 downto 0);
signal VN937_sign_out : std_logic_vector(5 downto 0);
signal VN938_data_out : std_logic_vector(5 downto 0);
signal VN938_sign_out : std_logic_vector(5 downto 0);
signal VN939_data_out : std_logic_vector(5 downto 0);
signal VN939_sign_out : std_logic_vector(5 downto 0);
signal VN940_data_out : std_logic_vector(5 downto 0);
signal VN940_sign_out : std_logic_vector(5 downto 0);
signal VN941_data_out : std_logic_vector(5 downto 0);
signal VN941_sign_out : std_logic_vector(5 downto 0);
signal VN942_data_out : std_logic_vector(5 downto 0);
signal VN942_sign_out : std_logic_vector(5 downto 0);
signal VN943_data_out : std_logic_vector(5 downto 0);
signal VN943_sign_out : std_logic_vector(5 downto 0);
signal VN944_data_out : std_logic_vector(5 downto 0);
signal VN944_sign_out : std_logic_vector(5 downto 0);
signal VN945_data_out : std_logic_vector(5 downto 0);
signal VN945_sign_out : std_logic_vector(5 downto 0);
signal VN946_data_out : std_logic_vector(5 downto 0);
signal VN946_sign_out : std_logic_vector(5 downto 0);
signal VN947_data_out : std_logic_vector(5 downto 0);
signal VN947_sign_out : std_logic_vector(5 downto 0);
signal VN948_data_out : std_logic_vector(5 downto 0);
signal VN948_sign_out : std_logic_vector(5 downto 0);
signal VN949_data_out : std_logic_vector(5 downto 0);
signal VN949_sign_out : std_logic_vector(5 downto 0);
signal VN950_data_out : std_logic_vector(5 downto 0);
signal VN950_sign_out : std_logic_vector(5 downto 0);
signal VN951_data_out : std_logic_vector(5 downto 0);
signal VN951_sign_out : std_logic_vector(5 downto 0);
signal VN952_data_out : std_logic_vector(5 downto 0);
signal VN952_sign_out : std_logic_vector(5 downto 0);
signal VN953_data_out : std_logic_vector(5 downto 0);
signal VN953_sign_out : std_logic_vector(5 downto 0);
signal VN954_data_out : std_logic_vector(5 downto 0);
signal VN954_sign_out : std_logic_vector(5 downto 0);
signal VN955_data_out : std_logic_vector(5 downto 0);
signal VN955_sign_out : std_logic_vector(5 downto 0);
signal VN956_data_out : std_logic_vector(5 downto 0);
signal VN956_sign_out : std_logic_vector(5 downto 0);
signal VN957_data_out : std_logic_vector(5 downto 0);
signal VN957_sign_out : std_logic_vector(5 downto 0);
signal VN958_data_out : std_logic_vector(5 downto 0);
signal VN958_sign_out : std_logic_vector(5 downto 0);
signal VN959_data_out : std_logic_vector(5 downto 0);
signal VN959_sign_out : std_logic_vector(5 downto 0);
signal VN960_data_out : std_logic_vector(5 downto 0);
signal VN960_sign_out : std_logic_vector(5 downto 0);
signal VN961_data_out : std_logic_vector(5 downto 0);
signal VN961_sign_out : std_logic_vector(5 downto 0);
signal VN962_data_out : std_logic_vector(5 downto 0);
signal VN962_sign_out : std_logic_vector(5 downto 0);
signal VN963_data_out : std_logic_vector(5 downto 0);
signal VN963_sign_out : std_logic_vector(5 downto 0);
signal VN964_data_out : std_logic_vector(5 downto 0);
signal VN964_sign_out : std_logic_vector(5 downto 0);
signal VN965_data_out : std_logic_vector(5 downto 0);
signal VN965_sign_out : std_logic_vector(5 downto 0);
signal VN966_data_out : std_logic_vector(5 downto 0);
signal VN966_sign_out : std_logic_vector(5 downto 0);
signal VN967_data_out : std_logic_vector(5 downto 0);
signal VN967_sign_out : std_logic_vector(5 downto 0);
signal VN968_data_out : std_logic_vector(5 downto 0);
signal VN968_sign_out : std_logic_vector(5 downto 0);
signal VN969_data_out : std_logic_vector(5 downto 0);
signal VN969_sign_out : std_logic_vector(5 downto 0);
signal VN970_data_out : std_logic_vector(5 downto 0);
signal VN970_sign_out : std_logic_vector(5 downto 0);
signal VN971_data_out : std_logic_vector(5 downto 0);
signal VN971_sign_out : std_logic_vector(5 downto 0);
signal VN972_data_out : std_logic_vector(5 downto 0);
signal VN972_sign_out : std_logic_vector(5 downto 0);
signal VN973_data_out : std_logic_vector(5 downto 0);
signal VN973_sign_out : std_logic_vector(5 downto 0);
signal VN974_data_out : std_logic_vector(5 downto 0);
signal VN974_sign_out : std_logic_vector(5 downto 0);
signal VN975_data_out : std_logic_vector(5 downto 0);
signal VN975_sign_out : std_logic_vector(5 downto 0);
signal VN976_data_out : std_logic_vector(5 downto 0);
signal VN976_sign_out : std_logic_vector(5 downto 0);
signal VN977_data_out : std_logic_vector(5 downto 0);
signal VN977_sign_out : std_logic_vector(5 downto 0);
signal VN978_data_out : std_logic_vector(5 downto 0);
signal VN978_sign_out : std_logic_vector(5 downto 0);
signal VN979_data_out : std_logic_vector(5 downto 0);
signal VN979_sign_out : std_logic_vector(5 downto 0);
signal VN980_data_out : std_logic_vector(5 downto 0);
signal VN980_sign_out : std_logic_vector(5 downto 0);
signal VN981_data_out : std_logic_vector(5 downto 0);
signal VN981_sign_out : std_logic_vector(5 downto 0);
signal VN982_data_out : std_logic_vector(5 downto 0);
signal VN982_sign_out : std_logic_vector(5 downto 0);
signal VN983_data_out : std_logic_vector(5 downto 0);
signal VN983_sign_out : std_logic_vector(5 downto 0);
signal VN984_data_out : std_logic_vector(5 downto 0);
signal VN984_sign_out : std_logic_vector(5 downto 0);
signal VN985_data_out : std_logic_vector(5 downto 0);
signal VN985_sign_out : std_logic_vector(5 downto 0);
signal VN986_data_out : std_logic_vector(5 downto 0);
signal VN986_sign_out : std_logic_vector(5 downto 0);
signal VN987_data_out : std_logic_vector(5 downto 0);
signal VN987_sign_out : std_logic_vector(5 downto 0);
signal VN988_data_out : std_logic_vector(5 downto 0);
signal VN988_sign_out : std_logic_vector(5 downto 0);
signal VN989_data_out : std_logic_vector(5 downto 0);
signal VN989_sign_out : std_logic_vector(5 downto 0);
signal VN990_data_out : std_logic_vector(5 downto 0);
signal VN990_sign_out : std_logic_vector(5 downto 0);
signal VN991_data_out : std_logic_vector(5 downto 0);
signal VN991_sign_out : std_logic_vector(5 downto 0);
signal VN992_data_out : std_logic_vector(5 downto 0);
signal VN992_sign_out : std_logic_vector(5 downto 0);
signal VN993_data_out : std_logic_vector(5 downto 0);
signal VN993_sign_out : std_logic_vector(5 downto 0);
signal VN994_data_out : std_logic_vector(5 downto 0);
signal VN994_sign_out : std_logic_vector(5 downto 0);
signal VN995_data_out : std_logic_vector(5 downto 0);
signal VN995_sign_out : std_logic_vector(5 downto 0);
signal VN996_data_out : std_logic_vector(5 downto 0);
signal VN996_sign_out : std_logic_vector(5 downto 0);
signal VN997_data_out : std_logic_vector(5 downto 0);
signal VN997_sign_out : std_logic_vector(5 downto 0);
signal VN998_data_out : std_logic_vector(5 downto 0);
signal VN998_sign_out : std_logic_vector(5 downto 0);
signal VN999_data_out : std_logic_vector(5 downto 0);
signal VN999_sign_out : std_logic_vector(5 downto 0);
signal VN1000_data_out : std_logic_vector(5 downto 0);
signal VN1000_sign_out : std_logic_vector(5 downto 0);
signal VN1001_data_out : std_logic_vector(5 downto 0);
signal VN1001_sign_out : std_logic_vector(5 downto 0);
signal VN1002_data_out : std_logic_vector(5 downto 0);
signal VN1002_sign_out : std_logic_vector(5 downto 0);
signal VN1003_data_out : std_logic_vector(5 downto 0);
signal VN1003_sign_out : std_logic_vector(5 downto 0);
signal VN1004_data_out : std_logic_vector(5 downto 0);
signal VN1004_sign_out : std_logic_vector(5 downto 0);
signal VN1005_data_out : std_logic_vector(5 downto 0);
signal VN1005_sign_out : std_logic_vector(5 downto 0);
signal VN1006_data_out : std_logic_vector(5 downto 0);
signal VN1006_sign_out : std_logic_vector(5 downto 0);
signal VN1007_data_out : std_logic_vector(5 downto 0);
signal VN1007_sign_out : std_logic_vector(5 downto 0);
signal VN1008_data_out : std_logic_vector(5 downto 0);
signal VN1008_sign_out : std_logic_vector(5 downto 0);
signal VN1009_data_out : std_logic_vector(5 downto 0);
signal VN1009_sign_out : std_logic_vector(5 downto 0);
signal VN1010_data_out : std_logic_vector(5 downto 0);
signal VN1010_sign_out : std_logic_vector(5 downto 0);
signal VN1011_data_out : std_logic_vector(5 downto 0);
signal VN1011_sign_out : std_logic_vector(5 downto 0);
signal VN1012_data_out : std_logic_vector(5 downto 0);
signal VN1012_sign_out : std_logic_vector(5 downto 0);
signal VN1013_data_out : std_logic_vector(5 downto 0);
signal VN1013_sign_out : std_logic_vector(5 downto 0);
signal VN1014_data_out : std_logic_vector(5 downto 0);
signal VN1014_sign_out : std_logic_vector(5 downto 0);
signal VN1015_data_out : std_logic_vector(5 downto 0);
signal VN1015_sign_out : std_logic_vector(5 downto 0);
signal VN1016_data_out : std_logic_vector(5 downto 0);
signal VN1016_sign_out : std_logic_vector(5 downto 0);
signal VN1017_data_out : std_logic_vector(5 downto 0);
signal VN1017_sign_out : std_logic_vector(5 downto 0);
signal VN1018_data_out : std_logic_vector(5 downto 0);
signal VN1018_sign_out : std_logic_vector(5 downto 0);
signal VN1019_data_out : std_logic_vector(5 downto 0);
signal VN1019_sign_out : std_logic_vector(5 downto 0);
signal VN1020_data_out : std_logic_vector(5 downto 0);
signal VN1020_sign_out : std_logic_vector(5 downto 0);
signal VN1021_data_out : std_logic_vector(5 downto 0);
signal VN1021_sign_out : std_logic_vector(5 downto 0);
signal VN1022_data_out : std_logic_vector(5 downto 0);
signal VN1022_sign_out : std_logic_vector(5 downto 0);
signal VN1023_data_out : std_logic_vector(5 downto 0);
signal VN1023_sign_out : std_logic_vector(5 downto 0);
signal VN1024_data_out : std_logic_vector(5 downto 0);
signal VN1024_sign_out : std_logic_vector(5 downto 0);
signal VN1025_data_out : std_logic_vector(5 downto 0);
signal VN1025_sign_out : std_logic_vector(5 downto 0);
signal VN1026_data_out : std_logic_vector(5 downto 0);
signal VN1026_sign_out : std_logic_vector(5 downto 0);
signal VN1027_data_out : std_logic_vector(5 downto 0);
signal VN1027_sign_out : std_logic_vector(5 downto 0);
signal VN1028_data_out : std_logic_vector(5 downto 0);
signal VN1028_sign_out : std_logic_vector(5 downto 0);
signal VN1029_data_out : std_logic_vector(5 downto 0);
signal VN1029_sign_out : std_logic_vector(5 downto 0);
signal VN1030_data_out : std_logic_vector(5 downto 0);
signal VN1030_sign_out : std_logic_vector(5 downto 0);
signal VN1031_data_out : std_logic_vector(5 downto 0);
signal VN1031_sign_out : std_logic_vector(5 downto 0);
signal VN1032_data_out : std_logic_vector(5 downto 0);
signal VN1032_sign_out : std_logic_vector(5 downto 0);
signal VN1033_data_out : std_logic_vector(5 downto 0);
signal VN1033_sign_out : std_logic_vector(5 downto 0);
signal VN1034_data_out : std_logic_vector(5 downto 0);
signal VN1034_sign_out : std_logic_vector(5 downto 0);
signal VN1035_data_out : std_logic_vector(5 downto 0);
signal VN1035_sign_out : std_logic_vector(5 downto 0);
signal VN1036_data_out : std_logic_vector(5 downto 0);
signal VN1036_sign_out : std_logic_vector(5 downto 0);
signal VN1037_data_out : std_logic_vector(5 downto 0);
signal VN1037_sign_out : std_logic_vector(5 downto 0);
signal VN1038_data_out : std_logic_vector(5 downto 0);
signal VN1038_sign_out : std_logic_vector(5 downto 0);
signal VN1039_data_out : std_logic_vector(5 downto 0);
signal VN1039_sign_out : std_logic_vector(5 downto 0);
signal VN1040_data_out : std_logic_vector(5 downto 0);
signal VN1040_sign_out : std_logic_vector(5 downto 0);
signal VN1041_data_out : std_logic_vector(5 downto 0);
signal VN1041_sign_out : std_logic_vector(5 downto 0);
signal VN1042_data_out : std_logic_vector(5 downto 0);
signal VN1042_sign_out : std_logic_vector(5 downto 0);
signal VN1043_data_out : std_logic_vector(5 downto 0);
signal VN1043_sign_out : std_logic_vector(5 downto 0);
signal VN1044_data_out : std_logic_vector(5 downto 0);
signal VN1044_sign_out : std_logic_vector(5 downto 0);
signal VN1045_data_out : std_logic_vector(5 downto 0);
signal VN1045_sign_out : std_logic_vector(5 downto 0);
signal VN1046_data_out : std_logic_vector(5 downto 0);
signal VN1046_sign_out : std_logic_vector(5 downto 0);
signal VN1047_data_out : std_logic_vector(5 downto 0);
signal VN1047_sign_out : std_logic_vector(5 downto 0);
signal VN1048_data_out : std_logic_vector(5 downto 0);
signal VN1048_sign_out : std_logic_vector(5 downto 0);
signal VN1049_data_out : std_logic_vector(5 downto 0);
signal VN1049_sign_out : std_logic_vector(5 downto 0);
signal VN1050_data_out : std_logic_vector(5 downto 0);
signal VN1050_sign_out : std_logic_vector(5 downto 0);
signal VN1051_data_out : std_logic_vector(5 downto 0);
signal VN1051_sign_out : std_logic_vector(5 downto 0);
signal VN1052_data_out : std_logic_vector(5 downto 0);
signal VN1052_sign_out : std_logic_vector(5 downto 0);
signal VN1053_data_out : std_logic_vector(5 downto 0);
signal VN1053_sign_out : std_logic_vector(5 downto 0);
signal VN1054_data_out : std_logic_vector(5 downto 0);
signal VN1054_sign_out : std_logic_vector(5 downto 0);
signal VN1055_data_out : std_logic_vector(5 downto 0);
signal VN1055_sign_out : std_logic_vector(5 downto 0);
signal VN1056_data_out : std_logic_vector(5 downto 0);
signal VN1056_sign_out : std_logic_vector(5 downto 0);
signal VN1057_data_out : std_logic_vector(5 downto 0);
signal VN1057_sign_out : std_logic_vector(5 downto 0);
signal VN1058_data_out : std_logic_vector(5 downto 0);
signal VN1058_sign_out : std_logic_vector(5 downto 0);
signal VN1059_data_out : std_logic_vector(5 downto 0);
signal VN1059_sign_out : std_logic_vector(5 downto 0);
signal VN1060_data_out : std_logic_vector(5 downto 0);
signal VN1060_sign_out : std_logic_vector(5 downto 0);
signal VN1061_data_out : std_logic_vector(5 downto 0);
signal VN1061_sign_out : std_logic_vector(5 downto 0);
signal VN1062_data_out : std_logic_vector(5 downto 0);
signal VN1062_sign_out : std_logic_vector(5 downto 0);
signal VN1063_data_out : std_logic_vector(5 downto 0);
signal VN1063_sign_out : std_logic_vector(5 downto 0);
signal VN1064_data_out : std_logic_vector(5 downto 0);
signal VN1064_sign_out : std_logic_vector(5 downto 0);
signal VN1065_data_out : std_logic_vector(5 downto 0);
signal VN1065_sign_out : std_logic_vector(5 downto 0);
signal VN1066_data_out : std_logic_vector(5 downto 0);
signal VN1066_sign_out : std_logic_vector(5 downto 0);
signal VN1067_data_out : std_logic_vector(5 downto 0);
signal VN1067_sign_out : std_logic_vector(5 downto 0);
signal VN1068_data_out : std_logic_vector(5 downto 0);
signal VN1068_sign_out : std_logic_vector(5 downto 0);
signal VN1069_data_out : std_logic_vector(5 downto 0);
signal VN1069_sign_out : std_logic_vector(5 downto 0);
signal VN1070_data_out : std_logic_vector(5 downto 0);
signal VN1070_sign_out : std_logic_vector(5 downto 0);
signal VN1071_data_out : std_logic_vector(5 downto 0);
signal VN1071_sign_out : std_logic_vector(5 downto 0);
signal VN1072_data_out : std_logic_vector(5 downto 0);
signal VN1072_sign_out : std_logic_vector(5 downto 0);
signal VN1073_data_out : std_logic_vector(5 downto 0);
signal VN1073_sign_out : std_logic_vector(5 downto 0);
signal VN1074_data_out : std_logic_vector(5 downto 0);
signal VN1074_sign_out : std_logic_vector(5 downto 0);
signal VN1075_data_out : std_logic_vector(5 downto 0);
signal VN1075_sign_out : std_logic_vector(5 downto 0);
signal VN1076_data_out : std_logic_vector(5 downto 0);
signal VN1076_sign_out : std_logic_vector(5 downto 0);
signal VN1077_data_out : std_logic_vector(5 downto 0);
signal VN1077_sign_out : std_logic_vector(5 downto 0);
signal VN1078_data_out : std_logic_vector(5 downto 0);
signal VN1078_sign_out : std_logic_vector(5 downto 0);
signal VN1079_data_out : std_logic_vector(5 downto 0);
signal VN1079_sign_out : std_logic_vector(5 downto 0);
signal VN1080_data_out : std_logic_vector(5 downto 0);
signal VN1080_sign_out : std_logic_vector(5 downto 0);
signal VN1081_data_out : std_logic_vector(5 downto 0);
signal VN1081_sign_out : std_logic_vector(5 downto 0);
signal VN1082_data_out : std_logic_vector(5 downto 0);
signal VN1082_sign_out : std_logic_vector(5 downto 0);
signal VN1083_data_out : std_logic_vector(5 downto 0);
signal VN1083_sign_out : std_logic_vector(5 downto 0);
signal VN1084_data_out : std_logic_vector(5 downto 0);
signal VN1084_sign_out : std_logic_vector(5 downto 0);
signal VN1085_data_out : std_logic_vector(5 downto 0);
signal VN1085_sign_out : std_logic_vector(5 downto 0);
signal VN1086_data_out : std_logic_vector(5 downto 0);
signal VN1086_sign_out : std_logic_vector(5 downto 0);
signal VN1087_data_out : std_logic_vector(5 downto 0);
signal VN1087_sign_out : std_logic_vector(5 downto 0);
signal VN1088_data_out : std_logic_vector(5 downto 0);
signal VN1088_sign_out : std_logic_vector(5 downto 0);
signal VN1089_data_out : std_logic_vector(5 downto 0);
signal VN1089_sign_out : std_logic_vector(5 downto 0);
signal VN1090_data_out : std_logic_vector(5 downto 0);
signal VN1090_sign_out : std_logic_vector(5 downto 0);
signal VN1091_data_out : std_logic_vector(5 downto 0);
signal VN1091_sign_out : std_logic_vector(5 downto 0);
signal VN1092_data_out : std_logic_vector(5 downto 0);
signal VN1092_sign_out : std_logic_vector(5 downto 0);
signal VN1093_data_out : std_logic_vector(5 downto 0);
signal VN1093_sign_out : std_logic_vector(5 downto 0);
signal VN1094_data_out : std_logic_vector(5 downto 0);
signal VN1094_sign_out : std_logic_vector(5 downto 0);
signal VN1095_data_out : std_logic_vector(5 downto 0);
signal VN1095_sign_out : std_logic_vector(5 downto 0);
signal VN1096_data_out : std_logic_vector(5 downto 0);
signal VN1096_sign_out : std_logic_vector(5 downto 0);
signal VN1097_data_out : std_logic_vector(5 downto 0);
signal VN1097_sign_out : std_logic_vector(5 downto 0);
signal VN1098_data_out : std_logic_vector(5 downto 0);
signal VN1098_sign_out : std_logic_vector(5 downto 0);
signal VN1099_data_out : std_logic_vector(5 downto 0);
signal VN1099_sign_out : std_logic_vector(5 downto 0);
signal VN1100_data_out : std_logic_vector(5 downto 0);
signal VN1100_sign_out : std_logic_vector(5 downto 0);
signal VN1101_data_out : std_logic_vector(5 downto 0);
signal VN1101_sign_out : std_logic_vector(5 downto 0);
signal VN1102_data_out : std_logic_vector(5 downto 0);
signal VN1102_sign_out : std_logic_vector(5 downto 0);
signal VN1103_data_out : std_logic_vector(5 downto 0);
signal VN1103_sign_out : std_logic_vector(5 downto 0);
signal VN1104_data_out : std_logic_vector(5 downto 0);
signal VN1104_sign_out : std_logic_vector(5 downto 0);
signal VN1105_data_out : std_logic_vector(5 downto 0);
signal VN1105_sign_out : std_logic_vector(5 downto 0);
signal VN1106_data_out : std_logic_vector(5 downto 0);
signal VN1106_sign_out : std_logic_vector(5 downto 0);
signal VN1107_data_out : std_logic_vector(5 downto 0);
signal VN1107_sign_out : std_logic_vector(5 downto 0);
signal VN1108_data_out : std_logic_vector(5 downto 0);
signal VN1108_sign_out : std_logic_vector(5 downto 0);
signal VN1109_data_out : std_logic_vector(5 downto 0);
signal VN1109_sign_out : std_logic_vector(5 downto 0);
signal VN1110_data_out : std_logic_vector(5 downto 0);
signal VN1110_sign_out : std_logic_vector(5 downto 0);
signal VN1111_data_out : std_logic_vector(5 downto 0);
signal VN1111_sign_out : std_logic_vector(5 downto 0);
signal VN1112_data_out : std_logic_vector(5 downto 0);
signal VN1112_sign_out : std_logic_vector(5 downto 0);
signal VN1113_data_out : std_logic_vector(5 downto 0);
signal VN1113_sign_out : std_logic_vector(5 downto 0);
signal VN1114_data_out : std_logic_vector(5 downto 0);
signal VN1114_sign_out : std_logic_vector(5 downto 0);
signal VN1115_data_out : std_logic_vector(5 downto 0);
signal VN1115_sign_out : std_logic_vector(5 downto 0);
signal VN1116_data_out : std_logic_vector(5 downto 0);
signal VN1116_sign_out : std_logic_vector(5 downto 0);
signal VN1117_data_out : std_logic_vector(5 downto 0);
signal VN1117_sign_out : std_logic_vector(5 downto 0);
signal VN1118_data_out : std_logic_vector(5 downto 0);
signal VN1118_sign_out : std_logic_vector(5 downto 0);
signal VN1119_data_out : std_logic_vector(5 downto 0);
signal VN1119_sign_out : std_logic_vector(5 downto 0);
signal VN1120_data_out : std_logic_vector(5 downto 0);
signal VN1120_sign_out : std_logic_vector(5 downto 0);
signal VN1121_data_out : std_logic_vector(5 downto 0);
signal VN1121_sign_out : std_logic_vector(5 downto 0);
signal VN1122_data_out : std_logic_vector(5 downto 0);
signal VN1122_sign_out : std_logic_vector(5 downto 0);
signal VN1123_data_out : std_logic_vector(5 downto 0);
signal VN1123_sign_out : std_logic_vector(5 downto 0);
signal VN1124_data_out : std_logic_vector(5 downto 0);
signal VN1124_sign_out : std_logic_vector(5 downto 0);
signal VN1125_data_out : std_logic_vector(5 downto 0);
signal VN1125_sign_out : std_logic_vector(5 downto 0);
signal VN1126_data_out : std_logic_vector(5 downto 0);
signal VN1126_sign_out : std_logic_vector(5 downto 0);
signal VN1127_data_out : std_logic_vector(5 downto 0);
signal VN1127_sign_out : std_logic_vector(5 downto 0);
signal VN1128_data_out : std_logic_vector(5 downto 0);
signal VN1128_sign_out : std_logic_vector(5 downto 0);
signal VN1129_data_out : std_logic_vector(5 downto 0);
signal VN1129_sign_out : std_logic_vector(5 downto 0);
signal VN1130_data_out : std_logic_vector(5 downto 0);
signal VN1130_sign_out : std_logic_vector(5 downto 0);
signal VN1131_data_out : std_logic_vector(5 downto 0);
signal VN1131_sign_out : std_logic_vector(5 downto 0);
signal VN1132_data_out : std_logic_vector(5 downto 0);
signal VN1132_sign_out : std_logic_vector(5 downto 0);
signal VN1133_data_out : std_logic_vector(5 downto 0);
signal VN1133_sign_out : std_logic_vector(5 downto 0);
signal VN1134_data_out : std_logic_vector(5 downto 0);
signal VN1134_sign_out : std_logic_vector(5 downto 0);
signal VN1135_data_out : std_logic_vector(5 downto 0);
signal VN1135_sign_out : std_logic_vector(5 downto 0);
signal VN1136_data_out : std_logic_vector(5 downto 0);
signal VN1136_sign_out : std_logic_vector(5 downto 0);
signal VN1137_data_out : std_logic_vector(5 downto 0);
signal VN1137_sign_out : std_logic_vector(5 downto 0);
signal VN1138_data_out : std_logic_vector(5 downto 0);
signal VN1138_sign_out : std_logic_vector(5 downto 0);
signal VN1139_data_out : std_logic_vector(5 downto 0);
signal VN1139_sign_out : std_logic_vector(5 downto 0);
signal VN1140_data_out : std_logic_vector(5 downto 0);
signal VN1140_sign_out : std_logic_vector(5 downto 0);
signal VN1141_data_out : std_logic_vector(5 downto 0);
signal VN1141_sign_out : std_logic_vector(5 downto 0);
signal VN1142_data_out : std_logic_vector(5 downto 0);
signal VN1142_sign_out : std_logic_vector(5 downto 0);
signal VN1143_data_out : std_logic_vector(5 downto 0);
signal VN1143_sign_out : std_logic_vector(5 downto 0);
signal VN1144_data_out : std_logic_vector(5 downto 0);
signal VN1144_sign_out : std_logic_vector(5 downto 0);
signal VN1145_data_out : std_logic_vector(5 downto 0);
signal VN1145_sign_out : std_logic_vector(5 downto 0);
signal VN1146_data_out : std_logic_vector(5 downto 0);
signal VN1146_sign_out : std_logic_vector(5 downto 0);
signal VN1147_data_out : std_logic_vector(5 downto 0);
signal VN1147_sign_out : std_logic_vector(5 downto 0);
signal VN1148_data_out : std_logic_vector(5 downto 0);
signal VN1148_sign_out : std_logic_vector(5 downto 0);
signal VN1149_data_out : std_logic_vector(5 downto 0);
signal VN1149_sign_out : std_logic_vector(5 downto 0);
signal VN1150_data_out : std_logic_vector(5 downto 0);
signal VN1150_sign_out : std_logic_vector(5 downto 0);
signal VN1151_data_out : std_logic_vector(5 downto 0);
signal VN1151_sign_out : std_logic_vector(5 downto 0);
signal VN1152_data_out : std_logic_vector(5 downto 0);
signal VN1152_sign_out : std_logic_vector(5 downto 0);
signal VN1153_data_out : std_logic_vector(5 downto 0);
signal VN1153_sign_out : std_logic_vector(5 downto 0);
signal VN1154_data_out : std_logic_vector(5 downto 0);
signal VN1154_sign_out : std_logic_vector(5 downto 0);
signal VN1155_data_out : std_logic_vector(5 downto 0);
signal VN1155_sign_out : std_logic_vector(5 downto 0);
signal VN1156_data_out : std_logic_vector(5 downto 0);
signal VN1156_sign_out : std_logic_vector(5 downto 0);
signal VN1157_data_out : std_logic_vector(5 downto 0);
signal VN1157_sign_out : std_logic_vector(5 downto 0);
signal VN1158_data_out : std_logic_vector(5 downto 0);
signal VN1158_sign_out : std_logic_vector(5 downto 0);
signal VN1159_data_out : std_logic_vector(5 downto 0);
signal VN1159_sign_out : std_logic_vector(5 downto 0);
signal VN1160_data_out : std_logic_vector(5 downto 0);
signal VN1160_sign_out : std_logic_vector(5 downto 0);
signal VN1161_data_out : std_logic_vector(5 downto 0);
signal VN1161_sign_out : std_logic_vector(5 downto 0);
signal VN1162_data_out : std_logic_vector(5 downto 0);
signal VN1162_sign_out : std_logic_vector(5 downto 0);
signal VN1163_data_out : std_logic_vector(5 downto 0);
signal VN1163_sign_out : std_logic_vector(5 downto 0);
signal VN1164_data_out : std_logic_vector(5 downto 0);
signal VN1164_sign_out : std_logic_vector(5 downto 0);
signal VN1165_data_out : std_logic_vector(5 downto 0);
signal VN1165_sign_out : std_logic_vector(5 downto 0);
signal VN1166_data_out : std_logic_vector(5 downto 0);
signal VN1166_sign_out : std_logic_vector(5 downto 0);
signal VN1167_data_out : std_logic_vector(5 downto 0);
signal VN1167_sign_out : std_logic_vector(5 downto 0);
signal VN1168_data_out : std_logic_vector(5 downto 0);
signal VN1168_sign_out : std_logic_vector(5 downto 0);
signal VN1169_data_out : std_logic_vector(5 downto 0);
signal VN1169_sign_out : std_logic_vector(5 downto 0);
signal VN1170_data_out : std_logic_vector(5 downto 0);
signal VN1170_sign_out : std_logic_vector(5 downto 0);
signal VN1171_data_out : std_logic_vector(5 downto 0);
signal VN1171_sign_out : std_logic_vector(5 downto 0);
signal VN1172_data_out : std_logic_vector(5 downto 0);
signal VN1172_sign_out : std_logic_vector(5 downto 0);
signal VN1173_data_out : std_logic_vector(5 downto 0);
signal VN1173_sign_out : std_logic_vector(5 downto 0);
signal VN1174_data_out : std_logic_vector(5 downto 0);
signal VN1174_sign_out : std_logic_vector(5 downto 0);
signal VN1175_data_out : std_logic_vector(5 downto 0);
signal VN1175_sign_out : std_logic_vector(5 downto 0);
signal VN1176_data_out : std_logic_vector(5 downto 0);
signal VN1176_sign_out : std_logic_vector(5 downto 0);
signal VN1177_data_out : std_logic_vector(5 downto 0);
signal VN1177_sign_out : std_logic_vector(5 downto 0);
signal VN1178_data_out : std_logic_vector(5 downto 0);
signal VN1178_sign_out : std_logic_vector(5 downto 0);
signal VN1179_data_out : std_logic_vector(5 downto 0);
signal VN1179_sign_out : std_logic_vector(5 downto 0);
signal VN1180_data_out : std_logic_vector(5 downto 0);
signal VN1180_sign_out : std_logic_vector(5 downto 0);
signal VN1181_data_out : std_logic_vector(5 downto 0);
signal VN1181_sign_out : std_logic_vector(5 downto 0);
signal VN1182_data_out : std_logic_vector(5 downto 0);
signal VN1182_sign_out : std_logic_vector(5 downto 0);
signal VN1183_data_out : std_logic_vector(5 downto 0);
signal VN1183_sign_out : std_logic_vector(5 downto 0);
signal VN1184_data_out : std_logic_vector(5 downto 0);
signal VN1184_sign_out : std_logic_vector(5 downto 0);
signal VN1185_data_out : std_logic_vector(5 downto 0);
signal VN1185_sign_out : std_logic_vector(5 downto 0);
signal VN1186_data_out : std_logic_vector(5 downto 0);
signal VN1186_sign_out : std_logic_vector(5 downto 0);
signal VN1187_data_out : std_logic_vector(5 downto 0);
signal VN1187_sign_out : std_logic_vector(5 downto 0);
signal VN1188_data_out : std_logic_vector(5 downto 0);
signal VN1188_sign_out : std_logic_vector(5 downto 0);
signal VN1189_data_out : std_logic_vector(5 downto 0);
signal VN1189_sign_out : std_logic_vector(5 downto 0);
signal VN1190_data_out : std_logic_vector(5 downto 0);
signal VN1190_sign_out : std_logic_vector(5 downto 0);
signal VN1191_data_out : std_logic_vector(5 downto 0);
signal VN1191_sign_out : std_logic_vector(5 downto 0);
signal VN1192_data_out : std_logic_vector(5 downto 0);
signal VN1192_sign_out : std_logic_vector(5 downto 0);
signal VN1193_data_out : std_logic_vector(5 downto 0);
signal VN1193_sign_out : std_logic_vector(5 downto 0);
signal VN1194_data_out : std_logic_vector(5 downto 0);
signal VN1194_sign_out : std_logic_vector(5 downto 0);
signal VN1195_data_out : std_logic_vector(5 downto 0);
signal VN1195_sign_out : std_logic_vector(5 downto 0);
signal VN1196_data_out : std_logic_vector(5 downto 0);
signal VN1196_sign_out : std_logic_vector(5 downto 0);
signal VN1197_data_out : std_logic_vector(5 downto 0);
signal VN1197_sign_out : std_logic_vector(5 downto 0);
signal VN1198_data_out : std_logic_vector(5 downto 0);
signal VN1198_sign_out : std_logic_vector(5 downto 0);
signal VN1199_data_out : std_logic_vector(5 downto 0);
signal VN1199_sign_out : std_logic_vector(5 downto 0);
signal VN1200_data_out : std_logic_vector(5 downto 0);
signal VN1200_sign_out : std_logic_vector(5 downto 0);
signal VN1201_data_out : std_logic_vector(5 downto 0);
signal VN1201_sign_out : std_logic_vector(5 downto 0);
signal VN1202_data_out : std_logic_vector(5 downto 0);
signal VN1202_sign_out : std_logic_vector(5 downto 0);
signal VN1203_data_out : std_logic_vector(5 downto 0);
signal VN1203_sign_out : std_logic_vector(5 downto 0);
signal VN1204_data_out : std_logic_vector(5 downto 0);
signal VN1204_sign_out : std_logic_vector(5 downto 0);
signal VN1205_data_out : std_logic_vector(5 downto 0);
signal VN1205_sign_out : std_logic_vector(5 downto 0);
signal VN1206_data_out : std_logic_vector(5 downto 0);
signal VN1206_sign_out : std_logic_vector(5 downto 0);
signal VN1207_data_out : std_logic_vector(5 downto 0);
signal VN1207_sign_out : std_logic_vector(5 downto 0);
signal VN1208_data_out : std_logic_vector(5 downto 0);
signal VN1208_sign_out : std_logic_vector(5 downto 0);
signal VN1209_data_out : std_logic_vector(5 downto 0);
signal VN1209_sign_out : std_logic_vector(5 downto 0);
signal VN1210_data_out : std_logic_vector(5 downto 0);
signal VN1210_sign_out : std_logic_vector(5 downto 0);
signal VN1211_data_out : std_logic_vector(5 downto 0);
signal VN1211_sign_out : std_logic_vector(5 downto 0);
signal VN1212_data_out : std_logic_vector(5 downto 0);
signal VN1212_sign_out : std_logic_vector(5 downto 0);
signal VN1213_data_out : std_logic_vector(5 downto 0);
signal VN1213_sign_out : std_logic_vector(5 downto 0);
signal VN1214_data_out : std_logic_vector(5 downto 0);
signal VN1214_sign_out : std_logic_vector(5 downto 0);
signal VN1215_data_out : std_logic_vector(5 downto 0);
signal VN1215_sign_out : std_logic_vector(5 downto 0);
signal VN1216_data_out : std_logic_vector(5 downto 0);
signal VN1216_sign_out : std_logic_vector(5 downto 0);
signal VN1217_data_out : std_logic_vector(5 downto 0);
signal VN1217_sign_out : std_logic_vector(5 downto 0);
signal VN1218_data_out : std_logic_vector(5 downto 0);
signal VN1218_sign_out : std_logic_vector(5 downto 0);
signal VN1219_data_out : std_logic_vector(5 downto 0);
signal VN1219_sign_out : std_logic_vector(5 downto 0);
signal VN1220_data_out : std_logic_vector(5 downto 0);
signal VN1220_sign_out : std_logic_vector(5 downto 0);
signal VN1221_data_out : std_logic_vector(5 downto 0);
signal VN1221_sign_out : std_logic_vector(5 downto 0);
signal VN1222_data_out : std_logic_vector(5 downto 0);
signal VN1222_sign_out : std_logic_vector(5 downto 0);
signal VN1223_data_out : std_logic_vector(5 downto 0);
signal VN1223_sign_out : std_logic_vector(5 downto 0);
signal VN1224_data_out : std_logic_vector(5 downto 0);
signal VN1224_sign_out : std_logic_vector(5 downto 0);
signal VN1225_data_out : std_logic_vector(5 downto 0);
signal VN1225_sign_out : std_logic_vector(5 downto 0);
signal VN1226_data_out : std_logic_vector(5 downto 0);
signal VN1226_sign_out : std_logic_vector(5 downto 0);
signal VN1227_data_out : std_logic_vector(5 downto 0);
signal VN1227_sign_out : std_logic_vector(5 downto 0);
signal VN1228_data_out : std_logic_vector(5 downto 0);
signal VN1228_sign_out : std_logic_vector(5 downto 0);
signal VN1229_data_out : std_logic_vector(5 downto 0);
signal VN1229_sign_out : std_logic_vector(5 downto 0);
signal VN1230_data_out : std_logic_vector(5 downto 0);
signal VN1230_sign_out : std_logic_vector(5 downto 0);
signal VN1231_data_out : std_logic_vector(5 downto 0);
signal VN1231_sign_out : std_logic_vector(5 downto 0);
signal VN1232_data_out : std_logic_vector(5 downto 0);
signal VN1232_sign_out : std_logic_vector(5 downto 0);
signal VN1233_data_out : std_logic_vector(5 downto 0);
signal VN1233_sign_out : std_logic_vector(5 downto 0);
signal VN1234_data_out : std_logic_vector(5 downto 0);
signal VN1234_sign_out : std_logic_vector(5 downto 0);
signal VN1235_data_out : std_logic_vector(5 downto 0);
signal VN1235_sign_out : std_logic_vector(5 downto 0);
signal VN1236_data_out : std_logic_vector(5 downto 0);
signal VN1236_sign_out : std_logic_vector(5 downto 0);
signal VN1237_data_out : std_logic_vector(5 downto 0);
signal VN1237_sign_out : std_logic_vector(5 downto 0);
signal VN1238_data_out : std_logic_vector(5 downto 0);
signal VN1238_sign_out : std_logic_vector(5 downto 0);
signal VN1239_data_out : std_logic_vector(5 downto 0);
signal VN1239_sign_out : std_logic_vector(5 downto 0);
signal VN1240_data_out : std_logic_vector(5 downto 0);
signal VN1240_sign_out : std_logic_vector(5 downto 0);
signal VN1241_data_out : std_logic_vector(5 downto 0);
signal VN1241_sign_out : std_logic_vector(5 downto 0);
signal VN1242_data_out : std_logic_vector(5 downto 0);
signal VN1242_sign_out : std_logic_vector(5 downto 0);
signal VN1243_data_out : std_logic_vector(5 downto 0);
signal VN1243_sign_out : std_logic_vector(5 downto 0);
signal VN1244_data_out : std_logic_vector(5 downto 0);
signal VN1244_sign_out : std_logic_vector(5 downto 0);
signal VN1245_data_out : std_logic_vector(5 downto 0);
signal VN1245_sign_out : std_logic_vector(5 downto 0);
signal VN1246_data_out : std_logic_vector(5 downto 0);
signal VN1246_sign_out : std_logic_vector(5 downto 0);
signal VN1247_data_out : std_logic_vector(5 downto 0);
signal VN1247_sign_out : std_logic_vector(5 downto 0);
signal VN1248_data_out : std_logic_vector(5 downto 0);
signal VN1248_sign_out : std_logic_vector(5 downto 0);
signal VN1249_data_out : std_logic_vector(5 downto 0);
signal VN1249_sign_out : std_logic_vector(5 downto 0);
signal VN1250_data_out : std_logic_vector(5 downto 0);
signal VN1250_sign_out : std_logic_vector(5 downto 0);
signal VN1251_data_out : std_logic_vector(5 downto 0);
signal VN1251_sign_out : std_logic_vector(5 downto 0);
signal VN1252_data_out : std_logic_vector(5 downto 0);
signal VN1252_sign_out : std_logic_vector(5 downto 0);
signal VN1253_data_out : std_logic_vector(5 downto 0);
signal VN1253_sign_out : std_logic_vector(5 downto 0);
signal VN1254_data_out : std_logic_vector(5 downto 0);
signal VN1254_sign_out : std_logic_vector(5 downto 0);
signal VN1255_data_out : std_logic_vector(5 downto 0);
signal VN1255_sign_out : std_logic_vector(5 downto 0);
signal VN1256_data_out : std_logic_vector(5 downto 0);
signal VN1256_sign_out : std_logic_vector(5 downto 0);
signal VN1257_data_out : std_logic_vector(5 downto 0);
signal VN1257_sign_out : std_logic_vector(5 downto 0);
signal VN1258_data_out : std_logic_vector(5 downto 0);
signal VN1258_sign_out : std_logic_vector(5 downto 0);
signal VN1259_data_out : std_logic_vector(5 downto 0);
signal VN1259_sign_out : std_logic_vector(5 downto 0);
signal VN1260_data_out : std_logic_vector(5 downto 0);
signal VN1260_sign_out : std_logic_vector(5 downto 0);
signal VN1261_data_out : std_logic_vector(5 downto 0);
signal VN1261_sign_out : std_logic_vector(5 downto 0);
signal VN1262_data_out : std_logic_vector(5 downto 0);
signal VN1262_sign_out : std_logic_vector(5 downto 0);
signal VN1263_data_out : std_logic_vector(5 downto 0);
signal VN1263_sign_out : std_logic_vector(5 downto 0);
signal VN1264_data_out : std_logic_vector(5 downto 0);
signal VN1264_sign_out : std_logic_vector(5 downto 0);
signal VN1265_data_out : std_logic_vector(5 downto 0);
signal VN1265_sign_out : std_logic_vector(5 downto 0);
signal VN1266_data_out : std_logic_vector(5 downto 0);
signal VN1266_sign_out : std_logic_vector(5 downto 0);
signal VN1267_data_out : std_logic_vector(5 downto 0);
signal VN1267_sign_out : std_logic_vector(5 downto 0);
signal VN1268_data_out : std_logic_vector(5 downto 0);
signal VN1268_sign_out : std_logic_vector(5 downto 0);
signal VN1269_data_out : std_logic_vector(5 downto 0);
signal VN1269_sign_out : std_logic_vector(5 downto 0);
signal VN1270_data_out : std_logic_vector(5 downto 0);
signal VN1270_sign_out : std_logic_vector(5 downto 0);
signal VN1271_data_out : std_logic_vector(5 downto 0);
signal VN1271_sign_out : std_logic_vector(5 downto 0);
signal VN1272_data_out : std_logic_vector(5 downto 0);
signal VN1272_sign_out : std_logic_vector(5 downto 0);
signal VN1273_data_out : std_logic_vector(5 downto 0);
signal VN1273_sign_out : std_logic_vector(5 downto 0);
signal VN1274_data_out : std_logic_vector(5 downto 0);
signal VN1274_sign_out : std_logic_vector(5 downto 0);
signal VN1275_data_out : std_logic_vector(5 downto 0);
signal VN1275_sign_out : std_logic_vector(5 downto 0);
signal VN1276_data_out : std_logic_vector(5 downto 0);
signal VN1276_sign_out : std_logic_vector(5 downto 0);
signal VN1277_data_out : std_logic_vector(5 downto 0);
signal VN1277_sign_out : std_logic_vector(5 downto 0);
signal VN1278_data_out : std_logic_vector(5 downto 0);
signal VN1278_sign_out : std_logic_vector(5 downto 0);
signal VN1279_data_out : std_logic_vector(5 downto 0);
signal VN1279_sign_out : std_logic_vector(5 downto 0);
signal VN1280_data_out : std_logic_vector(5 downto 0);
signal VN1280_sign_out : std_logic_vector(5 downto 0);
signal VN1281_data_out : std_logic_vector(5 downto 0);
signal VN1281_sign_out : std_logic_vector(5 downto 0);
signal VN1282_data_out : std_logic_vector(5 downto 0);
signal VN1282_sign_out : std_logic_vector(5 downto 0);
signal VN1283_data_out : std_logic_vector(5 downto 0);
signal VN1283_sign_out : std_logic_vector(5 downto 0);
signal VN1284_data_out : std_logic_vector(5 downto 0);
signal VN1284_sign_out : std_logic_vector(5 downto 0);
signal VN1285_data_out : std_logic_vector(5 downto 0);
signal VN1285_sign_out : std_logic_vector(5 downto 0);
signal VN1286_data_out : std_logic_vector(5 downto 0);
signal VN1286_sign_out : std_logic_vector(5 downto 0);
signal VN1287_data_out : std_logic_vector(5 downto 0);
signal VN1287_sign_out : std_logic_vector(5 downto 0);
signal VN1288_data_out : std_logic_vector(5 downto 0);
signal VN1288_sign_out : std_logic_vector(5 downto 0);
signal VN1289_data_out : std_logic_vector(5 downto 0);
signal VN1289_sign_out : std_logic_vector(5 downto 0);
signal VN1290_data_out : std_logic_vector(5 downto 0);
signal VN1290_sign_out : std_logic_vector(5 downto 0);
signal VN1291_data_out : std_logic_vector(5 downto 0);
signal VN1291_sign_out : std_logic_vector(5 downto 0);
signal VN1292_data_out : std_logic_vector(5 downto 0);
signal VN1292_sign_out : std_logic_vector(5 downto 0);
signal VN1293_data_out : std_logic_vector(5 downto 0);
signal VN1293_sign_out : std_logic_vector(5 downto 0);
signal VN1294_data_out : std_logic_vector(5 downto 0);
signal VN1294_sign_out : std_logic_vector(5 downto 0);
signal VN1295_data_out : std_logic_vector(5 downto 0);
signal VN1295_sign_out : std_logic_vector(5 downto 0);
signal VN1296_data_out : std_logic_vector(5 downto 0);
signal VN1296_sign_out : std_logic_vector(5 downto 0);
signal VN1297_data_out : std_logic_vector(5 downto 0);
signal VN1297_sign_out : std_logic_vector(5 downto 0);
signal VN1298_data_out : std_logic_vector(5 downto 0);
signal VN1298_sign_out : std_logic_vector(5 downto 0);
signal VN1299_data_out : std_logic_vector(5 downto 0);
signal VN1299_sign_out : std_logic_vector(5 downto 0);
signal VN1300_data_out : std_logic_vector(5 downto 0);
signal VN1300_sign_out : std_logic_vector(5 downto 0);
signal VN1301_data_out : std_logic_vector(5 downto 0);
signal VN1301_sign_out : std_logic_vector(5 downto 0);
signal VN1302_data_out : std_logic_vector(5 downto 0);
signal VN1302_sign_out : std_logic_vector(5 downto 0);
signal VN1303_data_out : std_logic_vector(5 downto 0);
signal VN1303_sign_out : std_logic_vector(5 downto 0);
signal VN1304_data_out : std_logic_vector(5 downto 0);
signal VN1304_sign_out : std_logic_vector(5 downto 0);
signal VN1305_data_out : std_logic_vector(5 downto 0);
signal VN1305_sign_out : std_logic_vector(5 downto 0);
signal VN1306_data_out : std_logic_vector(5 downto 0);
signal VN1306_sign_out : std_logic_vector(5 downto 0);
signal VN1307_data_out : std_logic_vector(5 downto 0);
signal VN1307_sign_out : std_logic_vector(5 downto 0);
signal VN1308_data_out : std_logic_vector(5 downto 0);
signal VN1308_sign_out : std_logic_vector(5 downto 0);
signal VN1309_data_out : std_logic_vector(5 downto 0);
signal VN1309_sign_out : std_logic_vector(5 downto 0);
signal VN1310_data_out : std_logic_vector(5 downto 0);
signal VN1310_sign_out : std_logic_vector(5 downto 0);
signal VN1311_data_out : std_logic_vector(5 downto 0);
signal VN1311_sign_out : std_logic_vector(5 downto 0);
signal VN1312_data_out : std_logic_vector(5 downto 0);
signal VN1312_sign_out : std_logic_vector(5 downto 0);
signal VN1313_data_out : std_logic_vector(5 downto 0);
signal VN1313_sign_out : std_logic_vector(5 downto 0);
signal VN1314_data_out : std_logic_vector(5 downto 0);
signal VN1314_sign_out : std_logic_vector(5 downto 0);
signal VN1315_data_out : std_logic_vector(5 downto 0);
signal VN1315_sign_out : std_logic_vector(5 downto 0);
signal VN1316_data_out : std_logic_vector(5 downto 0);
signal VN1316_sign_out : std_logic_vector(5 downto 0);
signal VN1317_data_out : std_logic_vector(5 downto 0);
signal VN1317_sign_out : std_logic_vector(5 downto 0);
signal VN1318_data_out : std_logic_vector(5 downto 0);
signal VN1318_sign_out : std_logic_vector(5 downto 0);
signal VN1319_data_out : std_logic_vector(5 downto 0);
signal VN1319_sign_out : std_logic_vector(5 downto 0);
signal VN1320_data_out : std_logic_vector(5 downto 0);
signal VN1320_sign_out : std_logic_vector(5 downto 0);
signal VN1321_data_out : std_logic_vector(5 downto 0);
signal VN1321_sign_out : std_logic_vector(5 downto 0);
signal VN1322_data_out : std_logic_vector(5 downto 0);
signal VN1322_sign_out : std_logic_vector(5 downto 0);
signal VN1323_data_out : std_logic_vector(5 downto 0);
signal VN1323_sign_out : std_logic_vector(5 downto 0);
signal VN1324_data_out : std_logic_vector(5 downto 0);
signal VN1324_sign_out : std_logic_vector(5 downto 0);
signal VN1325_data_out : std_logic_vector(5 downto 0);
signal VN1325_sign_out : std_logic_vector(5 downto 0);
signal VN1326_data_out : std_logic_vector(5 downto 0);
signal VN1326_sign_out : std_logic_vector(5 downto 0);
signal VN1327_data_out : std_logic_vector(5 downto 0);
signal VN1327_sign_out : std_logic_vector(5 downto 0);
signal VN1328_data_out : std_logic_vector(5 downto 0);
signal VN1328_sign_out : std_logic_vector(5 downto 0);
signal VN1329_data_out : std_logic_vector(5 downto 0);
signal VN1329_sign_out : std_logic_vector(5 downto 0);
signal VN1330_data_out : std_logic_vector(5 downto 0);
signal VN1330_sign_out : std_logic_vector(5 downto 0);
signal VN1331_data_out : std_logic_vector(5 downto 0);
signal VN1331_sign_out : std_logic_vector(5 downto 0);
signal VN1332_data_out : std_logic_vector(5 downto 0);
signal VN1332_sign_out : std_logic_vector(5 downto 0);
signal VN1333_data_out : std_logic_vector(5 downto 0);
signal VN1333_sign_out : std_logic_vector(5 downto 0);
signal VN1334_data_out : std_logic_vector(5 downto 0);
signal VN1334_sign_out : std_logic_vector(5 downto 0);
signal VN1335_data_out : std_logic_vector(5 downto 0);
signal VN1335_sign_out : std_logic_vector(5 downto 0);
signal VN1336_data_out : std_logic_vector(5 downto 0);
signal VN1336_sign_out : std_logic_vector(5 downto 0);
signal VN1337_data_out : std_logic_vector(5 downto 0);
signal VN1337_sign_out : std_logic_vector(5 downto 0);
signal VN1338_data_out : std_logic_vector(5 downto 0);
signal VN1338_sign_out : std_logic_vector(5 downto 0);
signal VN1339_data_out : std_logic_vector(5 downto 0);
signal VN1339_sign_out : std_logic_vector(5 downto 0);
signal VN1340_data_out : std_logic_vector(5 downto 0);
signal VN1340_sign_out : std_logic_vector(5 downto 0);
signal VN1341_data_out : std_logic_vector(5 downto 0);
signal VN1341_sign_out : std_logic_vector(5 downto 0);
signal VN1342_data_out : std_logic_vector(5 downto 0);
signal VN1342_sign_out : std_logic_vector(5 downto 0);
signal VN1343_data_out : std_logic_vector(5 downto 0);
signal VN1343_sign_out : std_logic_vector(5 downto 0);
signal VN1344_data_out : std_logic_vector(5 downto 0);
signal VN1344_sign_out : std_logic_vector(5 downto 0);
signal VN1345_data_out : std_logic_vector(5 downto 0);
signal VN1345_sign_out : std_logic_vector(5 downto 0);
signal VN1346_data_out : std_logic_vector(5 downto 0);
signal VN1346_sign_out : std_logic_vector(5 downto 0);
signal VN1347_data_out : std_logic_vector(5 downto 0);
signal VN1347_sign_out : std_logic_vector(5 downto 0);
signal VN1348_data_out : std_logic_vector(5 downto 0);
signal VN1348_sign_out : std_logic_vector(5 downto 0);
signal VN1349_data_out : std_logic_vector(5 downto 0);
signal VN1349_sign_out : std_logic_vector(5 downto 0);
signal VN1350_data_out : std_logic_vector(5 downto 0);
signal VN1350_sign_out : std_logic_vector(5 downto 0);
signal VN1351_data_out : std_logic_vector(5 downto 0);
signal VN1351_sign_out : std_logic_vector(5 downto 0);
signal VN1352_data_out : std_logic_vector(5 downto 0);
signal VN1352_sign_out : std_logic_vector(5 downto 0);
signal VN1353_data_out : std_logic_vector(5 downto 0);
signal VN1353_sign_out : std_logic_vector(5 downto 0);
signal VN1354_data_out : std_logic_vector(5 downto 0);
signal VN1354_sign_out : std_logic_vector(5 downto 0);
signal VN1355_data_out : std_logic_vector(5 downto 0);
signal VN1355_sign_out : std_logic_vector(5 downto 0);
signal VN1356_data_out : std_logic_vector(5 downto 0);
signal VN1356_sign_out : std_logic_vector(5 downto 0);
signal VN1357_data_out : std_logic_vector(5 downto 0);
signal VN1357_sign_out : std_logic_vector(5 downto 0);
signal VN1358_data_out : std_logic_vector(5 downto 0);
signal VN1358_sign_out : std_logic_vector(5 downto 0);
signal VN1359_data_out : std_logic_vector(5 downto 0);
signal VN1359_sign_out : std_logic_vector(5 downto 0);
signal VN1360_data_out : std_logic_vector(5 downto 0);
signal VN1360_sign_out : std_logic_vector(5 downto 0);
signal VN1361_data_out : std_logic_vector(5 downto 0);
signal VN1361_sign_out : std_logic_vector(5 downto 0);
signal VN1362_data_out : std_logic_vector(5 downto 0);
signal VN1362_sign_out : std_logic_vector(5 downto 0);
signal VN1363_data_out : std_logic_vector(5 downto 0);
signal VN1363_sign_out : std_logic_vector(5 downto 0);
signal VN1364_data_out : std_logic_vector(5 downto 0);
signal VN1364_sign_out : std_logic_vector(5 downto 0);
signal VN1365_data_out : std_logic_vector(5 downto 0);
signal VN1365_sign_out : std_logic_vector(5 downto 0);
signal VN1366_data_out : std_logic_vector(5 downto 0);
signal VN1366_sign_out : std_logic_vector(5 downto 0);
signal VN1367_data_out : std_logic_vector(5 downto 0);
signal VN1367_sign_out : std_logic_vector(5 downto 0);
signal VN1368_data_out : std_logic_vector(5 downto 0);
signal VN1368_sign_out : std_logic_vector(5 downto 0);
signal VN1369_data_out : std_logic_vector(5 downto 0);
signal VN1369_sign_out : std_logic_vector(5 downto 0);
signal VN1370_data_out : std_logic_vector(5 downto 0);
signal VN1370_sign_out : std_logic_vector(5 downto 0);
signal VN1371_data_out : std_logic_vector(5 downto 0);
signal VN1371_sign_out : std_logic_vector(5 downto 0);
signal VN1372_data_out : std_logic_vector(5 downto 0);
signal VN1372_sign_out : std_logic_vector(5 downto 0);
signal VN1373_data_out : std_logic_vector(5 downto 0);
signal VN1373_sign_out : std_logic_vector(5 downto 0);
signal VN1374_data_out : std_logic_vector(5 downto 0);
signal VN1374_sign_out : std_logic_vector(5 downto 0);
signal VN1375_data_out : std_logic_vector(5 downto 0);
signal VN1375_sign_out : std_logic_vector(5 downto 0);
signal VN1376_data_out : std_logic_vector(5 downto 0);
signal VN1376_sign_out : std_logic_vector(5 downto 0);
signal VN1377_data_out : std_logic_vector(5 downto 0);
signal VN1377_sign_out : std_logic_vector(5 downto 0);
signal VN1378_data_out : std_logic_vector(5 downto 0);
signal VN1378_sign_out : std_logic_vector(5 downto 0);
signal VN1379_data_out : std_logic_vector(5 downto 0);
signal VN1379_sign_out : std_logic_vector(5 downto 0);
signal VN1380_data_out : std_logic_vector(5 downto 0);
signal VN1380_sign_out : std_logic_vector(5 downto 0);
signal VN1381_data_out : std_logic_vector(5 downto 0);
signal VN1381_sign_out : std_logic_vector(5 downto 0);
signal VN1382_data_out : std_logic_vector(5 downto 0);
signal VN1382_sign_out : std_logic_vector(5 downto 0);
signal VN1383_data_out : std_logic_vector(5 downto 0);
signal VN1383_sign_out : std_logic_vector(5 downto 0);
signal VN1384_data_out : std_logic_vector(5 downto 0);
signal VN1384_sign_out : std_logic_vector(5 downto 0);
signal VN1385_data_out : std_logic_vector(5 downto 0);
signal VN1385_sign_out : std_logic_vector(5 downto 0);
signal VN1386_data_out : std_logic_vector(5 downto 0);
signal VN1386_sign_out : std_logic_vector(5 downto 0);
signal VN1387_data_out : std_logic_vector(5 downto 0);
signal VN1387_sign_out : std_logic_vector(5 downto 0);
signal VN1388_data_out : std_logic_vector(5 downto 0);
signal VN1388_sign_out : std_logic_vector(5 downto 0);
signal VN1389_data_out : std_logic_vector(5 downto 0);
signal VN1389_sign_out : std_logic_vector(5 downto 0);
signal VN1390_data_out : std_logic_vector(5 downto 0);
signal VN1390_sign_out : std_logic_vector(5 downto 0);
signal VN1391_data_out : std_logic_vector(5 downto 0);
signal VN1391_sign_out : std_logic_vector(5 downto 0);
signal VN1392_data_out : std_logic_vector(5 downto 0);
signal VN1392_sign_out : std_logic_vector(5 downto 0);
signal VN1393_data_out : std_logic_vector(5 downto 0);
signal VN1393_sign_out : std_logic_vector(5 downto 0);
signal VN1394_data_out : std_logic_vector(5 downto 0);
signal VN1394_sign_out : std_logic_vector(5 downto 0);
signal VN1395_data_out : std_logic_vector(5 downto 0);
signal VN1395_sign_out : std_logic_vector(5 downto 0);
signal VN1396_data_out : std_logic_vector(5 downto 0);
signal VN1396_sign_out : std_logic_vector(5 downto 0);
signal VN1397_data_out : std_logic_vector(5 downto 0);
signal VN1397_sign_out : std_logic_vector(5 downto 0);
signal VN1398_data_out : std_logic_vector(5 downto 0);
signal VN1398_sign_out : std_logic_vector(5 downto 0);
signal VN1399_data_out : std_logic_vector(5 downto 0);
signal VN1399_sign_out : std_logic_vector(5 downto 0);
signal VN1400_data_out : std_logic_vector(5 downto 0);
signal VN1400_sign_out : std_logic_vector(5 downto 0);
signal VN1401_data_out : std_logic_vector(5 downto 0);
signal VN1401_sign_out : std_logic_vector(5 downto 0);
signal VN1402_data_out : std_logic_vector(5 downto 0);
signal VN1402_sign_out : std_logic_vector(5 downto 0);
signal VN1403_data_out : std_logic_vector(5 downto 0);
signal VN1403_sign_out : std_logic_vector(5 downto 0);
signal VN1404_data_out : std_logic_vector(5 downto 0);
signal VN1404_sign_out : std_logic_vector(5 downto 0);
signal VN1405_data_out : std_logic_vector(5 downto 0);
signal VN1405_sign_out : std_logic_vector(5 downto 0);
signal VN1406_data_out : std_logic_vector(5 downto 0);
signal VN1406_sign_out : std_logic_vector(5 downto 0);
signal VN1407_data_out : std_logic_vector(5 downto 0);
signal VN1407_sign_out : std_logic_vector(5 downto 0);
signal VN1408_data_out : std_logic_vector(5 downto 0);
signal VN1408_sign_out : std_logic_vector(5 downto 0);
signal VN1409_data_out : std_logic_vector(5 downto 0);
signal VN1409_sign_out : std_logic_vector(5 downto 0);
signal VN1410_data_out : std_logic_vector(5 downto 0);
signal VN1410_sign_out : std_logic_vector(5 downto 0);
signal VN1411_data_out : std_logic_vector(5 downto 0);
signal VN1411_sign_out : std_logic_vector(5 downto 0);
signal VN1412_data_out : std_logic_vector(5 downto 0);
signal VN1412_sign_out : std_logic_vector(5 downto 0);
signal VN1413_data_out : std_logic_vector(5 downto 0);
signal VN1413_sign_out : std_logic_vector(5 downto 0);
signal VN1414_data_out : std_logic_vector(5 downto 0);
signal VN1414_sign_out : std_logic_vector(5 downto 0);
signal VN1415_data_out : std_logic_vector(5 downto 0);
signal VN1415_sign_out : std_logic_vector(5 downto 0);
signal VN1416_data_out : std_logic_vector(5 downto 0);
signal VN1416_sign_out : std_logic_vector(5 downto 0);
signal VN1417_data_out : std_logic_vector(5 downto 0);
signal VN1417_sign_out : std_logic_vector(5 downto 0);
signal VN1418_data_out : std_logic_vector(5 downto 0);
signal VN1418_sign_out : std_logic_vector(5 downto 0);
signal VN1419_data_out : std_logic_vector(5 downto 0);
signal VN1419_sign_out : std_logic_vector(5 downto 0);
signal VN1420_data_out : std_logic_vector(5 downto 0);
signal VN1420_sign_out : std_logic_vector(5 downto 0);
signal VN1421_data_out : std_logic_vector(5 downto 0);
signal VN1421_sign_out : std_logic_vector(5 downto 0);
signal VN1422_data_out : std_logic_vector(5 downto 0);
signal VN1422_sign_out : std_logic_vector(5 downto 0);
signal VN1423_data_out : std_logic_vector(5 downto 0);
signal VN1423_sign_out : std_logic_vector(5 downto 0);
signal VN1424_data_out : std_logic_vector(5 downto 0);
signal VN1424_sign_out : std_logic_vector(5 downto 0);
signal VN1425_data_out : std_logic_vector(5 downto 0);
signal VN1425_sign_out : std_logic_vector(5 downto 0);
signal VN1426_data_out : std_logic_vector(5 downto 0);
signal VN1426_sign_out : std_logic_vector(5 downto 0);
signal VN1427_data_out : std_logic_vector(5 downto 0);
signal VN1427_sign_out : std_logic_vector(5 downto 0);
signal VN1428_data_out : std_logic_vector(5 downto 0);
signal VN1428_sign_out : std_logic_vector(5 downto 0);
signal VN1429_data_out : std_logic_vector(5 downto 0);
signal VN1429_sign_out : std_logic_vector(5 downto 0);
signal VN1430_data_out : std_logic_vector(5 downto 0);
signal VN1430_sign_out : std_logic_vector(5 downto 0);
signal VN1431_data_out : std_logic_vector(5 downto 0);
signal VN1431_sign_out : std_logic_vector(5 downto 0);
signal VN1432_data_out : std_logic_vector(5 downto 0);
signal VN1432_sign_out : std_logic_vector(5 downto 0);
signal VN1433_data_out : std_logic_vector(5 downto 0);
signal VN1433_sign_out : std_logic_vector(5 downto 0);
signal VN1434_data_out : std_logic_vector(5 downto 0);
signal VN1434_sign_out : std_logic_vector(5 downto 0);
signal VN1435_data_out : std_logic_vector(5 downto 0);
signal VN1435_sign_out : std_logic_vector(5 downto 0);
signal VN1436_data_out : std_logic_vector(5 downto 0);
signal VN1436_sign_out : std_logic_vector(5 downto 0);
signal VN1437_data_out : std_logic_vector(5 downto 0);
signal VN1437_sign_out : std_logic_vector(5 downto 0);
signal VN1438_data_out : std_logic_vector(5 downto 0);
signal VN1438_sign_out : std_logic_vector(5 downto 0);
signal VN1439_data_out : std_logic_vector(5 downto 0);
signal VN1439_sign_out : std_logic_vector(5 downto 0);
signal VN1440_data_out : std_logic_vector(5 downto 0);
signal VN1440_sign_out : std_logic_vector(5 downto 0);
signal VN1441_data_out : std_logic_vector(5 downto 0);
signal VN1441_sign_out : std_logic_vector(5 downto 0);
signal VN1442_data_out : std_logic_vector(5 downto 0);
signal VN1442_sign_out : std_logic_vector(5 downto 0);
signal VN1443_data_out : std_logic_vector(5 downto 0);
signal VN1443_sign_out : std_logic_vector(5 downto 0);
signal VN1444_data_out : std_logic_vector(5 downto 0);
signal VN1444_sign_out : std_logic_vector(5 downto 0);
signal VN1445_data_out : std_logic_vector(5 downto 0);
signal VN1445_sign_out : std_logic_vector(5 downto 0);
signal VN1446_data_out : std_logic_vector(5 downto 0);
signal VN1446_sign_out : std_logic_vector(5 downto 0);
signal VN1447_data_out : std_logic_vector(5 downto 0);
signal VN1447_sign_out : std_logic_vector(5 downto 0);
signal VN1448_data_out : std_logic_vector(5 downto 0);
signal VN1448_sign_out : std_logic_vector(5 downto 0);
signal VN1449_data_out : std_logic_vector(5 downto 0);
signal VN1449_sign_out : std_logic_vector(5 downto 0);
signal VN1450_data_out : std_logic_vector(5 downto 0);
signal VN1450_sign_out : std_logic_vector(5 downto 0);
signal VN1451_data_out : std_logic_vector(5 downto 0);
signal VN1451_sign_out : std_logic_vector(5 downto 0);
signal VN1452_data_out : std_logic_vector(5 downto 0);
signal VN1452_sign_out : std_logic_vector(5 downto 0);
signal VN1453_data_out : std_logic_vector(5 downto 0);
signal VN1453_sign_out : std_logic_vector(5 downto 0);
signal VN1454_data_out : std_logic_vector(5 downto 0);
signal VN1454_sign_out : std_logic_vector(5 downto 0);
signal VN1455_data_out : std_logic_vector(5 downto 0);
signal VN1455_sign_out : std_logic_vector(5 downto 0);
signal VN1456_data_out : std_logic_vector(5 downto 0);
signal VN1456_sign_out : std_logic_vector(5 downto 0);
signal VN1457_data_out : std_logic_vector(5 downto 0);
signal VN1457_sign_out : std_logic_vector(5 downto 0);
signal VN1458_data_out : std_logic_vector(5 downto 0);
signal VN1458_sign_out : std_logic_vector(5 downto 0);
signal VN1459_data_out : std_logic_vector(5 downto 0);
signal VN1459_sign_out : std_logic_vector(5 downto 0);
signal VN1460_data_out : std_logic_vector(5 downto 0);
signal VN1460_sign_out : std_logic_vector(5 downto 0);
signal VN1461_data_out : std_logic_vector(5 downto 0);
signal VN1461_sign_out : std_logic_vector(5 downto 0);
signal VN1462_data_out : std_logic_vector(5 downto 0);
signal VN1462_sign_out : std_logic_vector(5 downto 0);
signal VN1463_data_out : std_logic_vector(5 downto 0);
signal VN1463_sign_out : std_logic_vector(5 downto 0);
signal VN1464_data_out : std_logic_vector(5 downto 0);
signal VN1464_sign_out : std_logic_vector(5 downto 0);
signal VN1465_data_out : std_logic_vector(5 downto 0);
signal VN1465_sign_out : std_logic_vector(5 downto 0);
signal VN1466_data_out : std_logic_vector(5 downto 0);
signal VN1466_sign_out : std_logic_vector(5 downto 0);
signal VN1467_data_out : std_logic_vector(5 downto 0);
signal VN1467_sign_out : std_logic_vector(5 downto 0);
signal VN1468_data_out : std_logic_vector(5 downto 0);
signal VN1468_sign_out : std_logic_vector(5 downto 0);
signal VN1469_data_out : std_logic_vector(5 downto 0);
signal VN1469_sign_out : std_logic_vector(5 downto 0);
signal VN1470_data_out : std_logic_vector(5 downto 0);
signal VN1470_sign_out : std_logic_vector(5 downto 0);
signal VN1471_data_out : std_logic_vector(5 downto 0);
signal VN1471_sign_out : std_logic_vector(5 downto 0);
signal VN1472_data_out : std_logic_vector(5 downto 0);
signal VN1472_sign_out : std_logic_vector(5 downto 0);
signal VN1473_data_out : std_logic_vector(5 downto 0);
signal VN1473_sign_out : std_logic_vector(5 downto 0);
signal VN1474_data_out : std_logic_vector(5 downto 0);
signal VN1474_sign_out : std_logic_vector(5 downto 0);
signal VN1475_data_out : std_logic_vector(5 downto 0);
signal VN1475_sign_out : std_logic_vector(5 downto 0);
signal VN1476_data_out : std_logic_vector(5 downto 0);
signal VN1476_sign_out : std_logic_vector(5 downto 0);
signal VN1477_data_out : std_logic_vector(5 downto 0);
signal VN1477_sign_out : std_logic_vector(5 downto 0);
signal VN1478_data_out : std_logic_vector(5 downto 0);
signal VN1478_sign_out : std_logic_vector(5 downto 0);
signal VN1479_data_out : std_logic_vector(5 downto 0);
signal VN1479_sign_out : std_logic_vector(5 downto 0);
signal VN1480_data_out : std_logic_vector(5 downto 0);
signal VN1480_sign_out : std_logic_vector(5 downto 0);
signal VN1481_data_out : std_logic_vector(5 downto 0);
signal VN1481_sign_out : std_logic_vector(5 downto 0);
signal VN1482_data_out : std_logic_vector(5 downto 0);
signal VN1482_sign_out : std_logic_vector(5 downto 0);
signal VN1483_data_out : std_logic_vector(5 downto 0);
signal VN1483_sign_out : std_logic_vector(5 downto 0);
signal VN1484_data_out : std_logic_vector(5 downto 0);
signal VN1484_sign_out : std_logic_vector(5 downto 0);
signal VN1485_data_out : std_logic_vector(5 downto 0);
signal VN1485_sign_out : std_logic_vector(5 downto 0);
signal VN1486_data_out : std_logic_vector(5 downto 0);
signal VN1486_sign_out : std_logic_vector(5 downto 0);
signal VN1487_data_out : std_logic_vector(5 downto 0);
signal VN1487_sign_out : std_logic_vector(5 downto 0);
signal VN1488_data_out : std_logic_vector(5 downto 0);
signal VN1488_sign_out : std_logic_vector(5 downto 0);
signal VN1489_data_out : std_logic_vector(5 downto 0);
signal VN1489_sign_out : std_logic_vector(5 downto 0);
signal VN1490_data_out : std_logic_vector(5 downto 0);
signal VN1490_sign_out : std_logic_vector(5 downto 0);
signal VN1491_data_out : std_logic_vector(5 downto 0);
signal VN1491_sign_out : std_logic_vector(5 downto 0);
signal VN1492_data_out : std_logic_vector(5 downto 0);
signal VN1492_sign_out : std_logic_vector(5 downto 0);
signal VN1493_data_out : std_logic_vector(5 downto 0);
signal VN1493_sign_out : std_logic_vector(5 downto 0);
signal VN1494_data_out : std_logic_vector(5 downto 0);
signal VN1494_sign_out : std_logic_vector(5 downto 0);
signal VN1495_data_out : std_logic_vector(5 downto 0);
signal VN1495_sign_out : std_logic_vector(5 downto 0);
signal VN1496_data_out : std_logic_vector(5 downto 0);
signal VN1496_sign_out : std_logic_vector(5 downto 0);
signal VN1497_data_out : std_logic_vector(5 downto 0);
signal VN1497_sign_out : std_logic_vector(5 downto 0);
signal VN1498_data_out : std_logic_vector(5 downto 0);
signal VN1498_sign_out : std_logic_vector(5 downto 0);
signal VN1499_data_out : std_logic_vector(5 downto 0);
signal VN1499_sign_out : std_logic_vector(5 downto 0);
signal VN1500_data_out : std_logic_vector(5 downto 0);
signal VN1500_sign_out : std_logic_vector(5 downto 0);
signal VN1501_data_out : std_logic_vector(5 downto 0);
signal VN1501_sign_out : std_logic_vector(5 downto 0);
signal VN1502_data_out : std_logic_vector(5 downto 0);
signal VN1502_sign_out : std_logic_vector(5 downto 0);
signal VN1503_data_out : std_logic_vector(5 downto 0);
signal VN1503_sign_out : std_logic_vector(5 downto 0);
signal VN1504_data_out : std_logic_vector(5 downto 0);
signal VN1504_sign_out : std_logic_vector(5 downto 0);
signal VN1505_data_out : std_logic_vector(5 downto 0);
signal VN1505_sign_out : std_logic_vector(5 downto 0);
signal VN1506_data_out : std_logic_vector(5 downto 0);
signal VN1506_sign_out : std_logic_vector(5 downto 0);
signal VN1507_data_out : std_logic_vector(5 downto 0);
signal VN1507_sign_out : std_logic_vector(5 downto 0);
signal VN1508_data_out : std_logic_vector(5 downto 0);
signal VN1508_sign_out : std_logic_vector(5 downto 0);
signal VN1509_data_out : std_logic_vector(5 downto 0);
signal VN1509_sign_out : std_logic_vector(5 downto 0);
signal VN1510_data_out : std_logic_vector(5 downto 0);
signal VN1510_sign_out : std_logic_vector(5 downto 0);
signal VN1511_data_out : std_logic_vector(5 downto 0);
signal VN1511_sign_out : std_logic_vector(5 downto 0);
signal VN1512_data_out : std_logic_vector(5 downto 0);
signal VN1512_sign_out : std_logic_vector(5 downto 0);
signal VN1513_data_out : std_logic_vector(5 downto 0);
signal VN1513_sign_out : std_logic_vector(5 downto 0);
signal VN1514_data_out : std_logic_vector(5 downto 0);
signal VN1514_sign_out : std_logic_vector(5 downto 0);
signal VN1515_data_out : std_logic_vector(5 downto 0);
signal VN1515_sign_out : std_logic_vector(5 downto 0);
signal VN1516_data_out : std_logic_vector(5 downto 0);
signal VN1516_sign_out : std_logic_vector(5 downto 0);
signal VN1517_data_out : std_logic_vector(5 downto 0);
signal VN1517_sign_out : std_logic_vector(5 downto 0);
signal VN1518_data_out : std_logic_vector(5 downto 0);
signal VN1518_sign_out : std_logic_vector(5 downto 0);
signal VN1519_data_out : std_logic_vector(5 downto 0);
signal VN1519_sign_out : std_logic_vector(5 downto 0);
signal VN1520_data_out : std_logic_vector(5 downto 0);
signal VN1520_sign_out : std_logic_vector(5 downto 0);
signal VN1521_data_out : std_logic_vector(5 downto 0);
signal VN1521_sign_out : std_logic_vector(5 downto 0);
signal VN1522_data_out : std_logic_vector(5 downto 0);
signal VN1522_sign_out : std_logic_vector(5 downto 0);
signal VN1523_data_out : std_logic_vector(5 downto 0);
signal VN1523_sign_out : std_logic_vector(5 downto 0);
signal VN1524_data_out : std_logic_vector(5 downto 0);
signal VN1524_sign_out : std_logic_vector(5 downto 0);
signal VN1525_data_out : std_logic_vector(5 downto 0);
signal VN1525_sign_out : std_logic_vector(5 downto 0);
signal VN1526_data_out : std_logic_vector(5 downto 0);
signal VN1526_sign_out : std_logic_vector(5 downto 0);
signal VN1527_data_out : std_logic_vector(5 downto 0);
signal VN1527_sign_out : std_logic_vector(5 downto 0);
signal VN1528_data_out : std_logic_vector(5 downto 0);
signal VN1528_sign_out : std_logic_vector(5 downto 0);
signal VN1529_data_out : std_logic_vector(5 downto 0);
signal VN1529_sign_out : std_logic_vector(5 downto 0);
signal VN1530_data_out : std_logic_vector(5 downto 0);
signal VN1530_sign_out : std_logic_vector(5 downto 0);
signal VN1531_data_out : std_logic_vector(5 downto 0);
signal VN1531_sign_out : std_logic_vector(5 downto 0);
signal VN1532_data_out : std_logic_vector(5 downto 0);
signal VN1532_sign_out : std_logic_vector(5 downto 0);
signal VN1533_data_out : std_logic_vector(5 downto 0);
signal VN1533_sign_out : std_logic_vector(5 downto 0);
signal VN1534_data_out : std_logic_vector(5 downto 0);
signal VN1534_sign_out : std_logic_vector(5 downto 0);
signal VN1535_data_out : std_logic_vector(5 downto 0);
signal VN1535_sign_out : std_logic_vector(5 downto 0);
signal VN1536_data_out : std_logic_vector(5 downto 0);
signal VN1536_sign_out : std_logic_vector(5 downto 0);
signal VN1537_data_out : std_logic_vector(5 downto 0);
signal VN1537_sign_out : std_logic_vector(5 downto 0);
signal VN1538_data_out : std_logic_vector(5 downto 0);
signal VN1538_sign_out : std_logic_vector(5 downto 0);
signal VN1539_data_out : std_logic_vector(5 downto 0);
signal VN1539_sign_out : std_logic_vector(5 downto 0);
signal VN1540_data_out : std_logic_vector(5 downto 0);
signal VN1540_sign_out : std_logic_vector(5 downto 0);
signal VN1541_data_out : std_logic_vector(5 downto 0);
signal VN1541_sign_out : std_logic_vector(5 downto 0);
signal VN1542_data_out : std_logic_vector(5 downto 0);
signal VN1542_sign_out : std_logic_vector(5 downto 0);
signal VN1543_data_out : std_logic_vector(5 downto 0);
signal VN1543_sign_out : std_logic_vector(5 downto 0);
signal VN1544_data_out : std_logic_vector(5 downto 0);
signal VN1544_sign_out : std_logic_vector(5 downto 0);
signal VN1545_data_out : std_logic_vector(5 downto 0);
signal VN1545_sign_out : std_logic_vector(5 downto 0);
signal VN1546_data_out : std_logic_vector(5 downto 0);
signal VN1546_sign_out : std_logic_vector(5 downto 0);
signal VN1547_data_out : std_logic_vector(5 downto 0);
signal VN1547_sign_out : std_logic_vector(5 downto 0);
signal VN1548_data_out : std_logic_vector(5 downto 0);
signal VN1548_sign_out : std_logic_vector(5 downto 0);
signal VN1549_data_out : std_logic_vector(5 downto 0);
signal VN1549_sign_out : std_logic_vector(5 downto 0);
signal VN1550_data_out : std_logic_vector(5 downto 0);
signal VN1550_sign_out : std_logic_vector(5 downto 0);
signal VN1551_data_out : std_logic_vector(5 downto 0);
signal VN1551_sign_out : std_logic_vector(5 downto 0);
signal VN1552_data_out : std_logic_vector(5 downto 0);
signal VN1552_sign_out : std_logic_vector(5 downto 0);
signal VN1553_data_out : std_logic_vector(5 downto 0);
signal VN1553_sign_out : std_logic_vector(5 downto 0);
signal VN1554_data_out : std_logic_vector(5 downto 0);
signal VN1554_sign_out : std_logic_vector(5 downto 0);
signal VN1555_data_out : std_logic_vector(5 downto 0);
signal VN1555_sign_out : std_logic_vector(5 downto 0);
signal VN1556_data_out : std_logic_vector(5 downto 0);
signal VN1556_sign_out : std_logic_vector(5 downto 0);
signal VN1557_data_out : std_logic_vector(5 downto 0);
signal VN1557_sign_out : std_logic_vector(5 downto 0);
signal VN1558_data_out : std_logic_vector(5 downto 0);
signal VN1558_sign_out : std_logic_vector(5 downto 0);
signal VN1559_data_out : std_logic_vector(5 downto 0);
signal VN1559_sign_out : std_logic_vector(5 downto 0);
signal VN1560_data_out : std_logic_vector(5 downto 0);
signal VN1560_sign_out : std_logic_vector(5 downto 0);
signal VN1561_data_out : std_logic_vector(5 downto 0);
signal VN1561_sign_out : std_logic_vector(5 downto 0);
signal VN1562_data_out : std_logic_vector(5 downto 0);
signal VN1562_sign_out : std_logic_vector(5 downto 0);
signal VN1563_data_out : std_logic_vector(5 downto 0);
signal VN1563_sign_out : std_logic_vector(5 downto 0);
signal VN1564_data_out : std_logic_vector(5 downto 0);
signal VN1564_sign_out : std_logic_vector(5 downto 0);
signal VN1565_data_out : std_logic_vector(5 downto 0);
signal VN1565_sign_out : std_logic_vector(5 downto 0);
signal VN1566_data_out : std_logic_vector(5 downto 0);
signal VN1566_sign_out : std_logic_vector(5 downto 0);
signal VN1567_data_out : std_logic_vector(5 downto 0);
signal VN1567_sign_out : std_logic_vector(5 downto 0);
signal VN1568_data_out : std_logic_vector(5 downto 0);
signal VN1568_sign_out : std_logic_vector(5 downto 0);
signal VN1569_data_out : std_logic_vector(5 downto 0);
signal VN1569_sign_out : std_logic_vector(5 downto 0);
signal VN1570_data_out : std_logic_vector(5 downto 0);
signal VN1570_sign_out : std_logic_vector(5 downto 0);
signal VN1571_data_out : std_logic_vector(5 downto 0);
signal VN1571_sign_out : std_logic_vector(5 downto 0);
signal VN1572_data_out : std_logic_vector(5 downto 0);
signal VN1572_sign_out : std_logic_vector(5 downto 0);
signal VN1573_data_out : std_logic_vector(5 downto 0);
signal VN1573_sign_out : std_logic_vector(5 downto 0);
signal VN1574_data_out : std_logic_vector(5 downto 0);
signal VN1574_sign_out : std_logic_vector(5 downto 0);
signal VN1575_data_out : std_logic_vector(5 downto 0);
signal VN1575_sign_out : std_logic_vector(5 downto 0);
signal VN1576_data_out : std_logic_vector(5 downto 0);
signal VN1576_sign_out : std_logic_vector(5 downto 0);
signal VN1577_data_out : std_logic_vector(5 downto 0);
signal VN1577_sign_out : std_logic_vector(5 downto 0);
signal VN1578_data_out : std_logic_vector(5 downto 0);
signal VN1578_sign_out : std_logic_vector(5 downto 0);
signal VN1579_data_out : std_logic_vector(5 downto 0);
signal VN1579_sign_out : std_logic_vector(5 downto 0);
signal VN1580_data_out : std_logic_vector(5 downto 0);
signal VN1580_sign_out : std_logic_vector(5 downto 0);
signal VN1581_data_out : std_logic_vector(5 downto 0);
signal VN1581_sign_out : std_logic_vector(5 downto 0);
signal VN1582_data_out : std_logic_vector(5 downto 0);
signal VN1582_sign_out : std_logic_vector(5 downto 0);
signal VN1583_data_out : std_logic_vector(5 downto 0);
signal VN1583_sign_out : std_logic_vector(5 downto 0);
signal VN1584_data_out : std_logic_vector(5 downto 0);
signal VN1584_sign_out : std_logic_vector(5 downto 0);
signal VN1585_data_out : std_logic_vector(5 downto 0);
signal VN1585_sign_out : std_logic_vector(5 downto 0);
signal VN1586_data_out : std_logic_vector(5 downto 0);
signal VN1586_sign_out : std_logic_vector(5 downto 0);
signal VN1587_data_out : std_logic_vector(5 downto 0);
signal VN1587_sign_out : std_logic_vector(5 downto 0);
signal VN1588_data_out : std_logic_vector(5 downto 0);
signal VN1588_sign_out : std_logic_vector(5 downto 0);
signal VN1589_data_out : std_logic_vector(5 downto 0);
signal VN1589_sign_out : std_logic_vector(5 downto 0);
signal VN1590_data_out : std_logic_vector(5 downto 0);
signal VN1590_sign_out : std_logic_vector(5 downto 0);
signal VN1591_data_out : std_logic_vector(5 downto 0);
signal VN1591_sign_out : std_logic_vector(5 downto 0);
signal VN1592_data_out : std_logic_vector(5 downto 0);
signal VN1592_sign_out : std_logic_vector(5 downto 0);
signal VN1593_data_out : std_logic_vector(5 downto 0);
signal VN1593_sign_out : std_logic_vector(5 downto 0);
signal VN1594_data_out : std_logic_vector(5 downto 0);
signal VN1594_sign_out : std_logic_vector(5 downto 0);
signal VN1595_data_out : std_logic_vector(5 downto 0);
signal VN1595_sign_out : std_logic_vector(5 downto 0);
signal VN1596_data_out : std_logic_vector(5 downto 0);
signal VN1596_sign_out : std_logic_vector(5 downto 0);
signal VN1597_data_out : std_logic_vector(5 downto 0);
signal VN1597_sign_out : std_logic_vector(5 downto 0);
signal VN1598_data_out : std_logic_vector(5 downto 0);
signal VN1598_sign_out : std_logic_vector(5 downto 0);
signal VN1599_data_out : std_logic_vector(5 downto 0);
signal VN1599_sign_out : std_logic_vector(5 downto 0);
signal VN1600_data_out : std_logic_vector(5 downto 0);
signal VN1600_sign_out : std_logic_vector(5 downto 0);
signal VN1601_data_out : std_logic_vector(5 downto 0);
signal VN1601_sign_out : std_logic_vector(5 downto 0);
signal VN1602_data_out : std_logic_vector(5 downto 0);
signal VN1602_sign_out : std_logic_vector(5 downto 0);
signal VN1603_data_out : std_logic_vector(5 downto 0);
signal VN1603_sign_out : std_logic_vector(5 downto 0);
signal VN1604_data_out : std_logic_vector(5 downto 0);
signal VN1604_sign_out : std_logic_vector(5 downto 0);
signal VN1605_data_out : std_logic_vector(5 downto 0);
signal VN1605_sign_out : std_logic_vector(5 downto 0);
signal VN1606_data_out : std_logic_vector(5 downto 0);
signal VN1606_sign_out : std_logic_vector(5 downto 0);
signal VN1607_data_out : std_logic_vector(5 downto 0);
signal VN1607_sign_out : std_logic_vector(5 downto 0);
signal VN1608_data_out : std_logic_vector(5 downto 0);
signal VN1608_sign_out : std_logic_vector(5 downto 0);
signal VN1609_data_out : std_logic_vector(5 downto 0);
signal VN1609_sign_out : std_logic_vector(5 downto 0);
signal VN1610_data_out : std_logic_vector(5 downto 0);
signal VN1610_sign_out : std_logic_vector(5 downto 0);
signal VN1611_data_out : std_logic_vector(5 downto 0);
signal VN1611_sign_out : std_logic_vector(5 downto 0);
signal VN1612_data_out : std_logic_vector(5 downto 0);
signal VN1612_sign_out : std_logic_vector(5 downto 0);
signal VN1613_data_out : std_logic_vector(5 downto 0);
signal VN1613_sign_out : std_logic_vector(5 downto 0);
signal VN1614_data_out : std_logic_vector(5 downto 0);
signal VN1614_sign_out : std_logic_vector(5 downto 0);
signal VN1615_data_out : std_logic_vector(5 downto 0);
signal VN1615_sign_out : std_logic_vector(5 downto 0);
signal VN1616_data_out : std_logic_vector(5 downto 0);
signal VN1616_sign_out : std_logic_vector(5 downto 0);
signal VN1617_data_out : std_logic_vector(5 downto 0);
signal VN1617_sign_out : std_logic_vector(5 downto 0);
signal VN1618_data_out : std_logic_vector(5 downto 0);
signal VN1618_sign_out : std_logic_vector(5 downto 0);
signal VN1619_data_out : std_logic_vector(5 downto 0);
signal VN1619_sign_out : std_logic_vector(5 downto 0);
signal VN1620_data_out : std_logic_vector(5 downto 0);
signal VN1620_sign_out : std_logic_vector(5 downto 0);
signal VN1621_data_out : std_logic_vector(5 downto 0);
signal VN1621_sign_out : std_logic_vector(5 downto 0);
signal VN1622_data_out : std_logic_vector(5 downto 0);
signal VN1622_sign_out : std_logic_vector(5 downto 0);
signal VN1623_data_out : std_logic_vector(5 downto 0);
signal VN1623_sign_out : std_logic_vector(5 downto 0);
signal VN1624_data_out : std_logic_vector(5 downto 0);
signal VN1624_sign_out : std_logic_vector(5 downto 0);
signal VN1625_data_out : std_logic_vector(5 downto 0);
signal VN1625_sign_out : std_logic_vector(5 downto 0);
signal VN1626_data_out : std_logic_vector(5 downto 0);
signal VN1626_sign_out : std_logic_vector(5 downto 0);
signal VN1627_data_out : std_logic_vector(5 downto 0);
signal VN1627_sign_out : std_logic_vector(5 downto 0);
signal VN1628_data_out : std_logic_vector(5 downto 0);
signal VN1628_sign_out : std_logic_vector(5 downto 0);
signal VN1629_data_out : std_logic_vector(5 downto 0);
signal VN1629_sign_out : std_logic_vector(5 downto 0);
signal VN1630_data_out : std_logic_vector(5 downto 0);
signal VN1630_sign_out : std_logic_vector(5 downto 0);
signal VN1631_data_out : std_logic_vector(5 downto 0);
signal VN1631_sign_out : std_logic_vector(5 downto 0);
signal VN1632_data_out : std_logic_vector(5 downto 0);
signal VN1632_sign_out : std_logic_vector(5 downto 0);
signal VN1633_data_out : std_logic_vector(5 downto 0);
signal VN1633_sign_out : std_logic_vector(5 downto 0);
signal VN1634_data_out : std_logic_vector(5 downto 0);
signal VN1634_sign_out : std_logic_vector(5 downto 0);
signal VN1635_data_out : std_logic_vector(5 downto 0);
signal VN1635_sign_out : std_logic_vector(5 downto 0);
signal VN1636_data_out : std_logic_vector(5 downto 0);
signal VN1636_sign_out : std_logic_vector(5 downto 0);
signal VN1637_data_out : std_logic_vector(5 downto 0);
signal VN1637_sign_out : std_logic_vector(5 downto 0);
signal VN1638_data_out : std_logic_vector(5 downto 0);
signal VN1638_sign_out : std_logic_vector(5 downto 0);
signal VN1639_data_out : std_logic_vector(5 downto 0);
signal VN1639_sign_out : std_logic_vector(5 downto 0);
signal VN1640_data_out : std_logic_vector(5 downto 0);
signal VN1640_sign_out : std_logic_vector(5 downto 0);
signal VN1641_data_out : std_logic_vector(5 downto 0);
signal VN1641_sign_out : std_logic_vector(5 downto 0);
signal VN1642_data_out : std_logic_vector(5 downto 0);
signal VN1642_sign_out : std_logic_vector(5 downto 0);
signal VN1643_data_out : std_logic_vector(5 downto 0);
signal VN1643_sign_out : std_logic_vector(5 downto 0);
signal VN1644_data_out : std_logic_vector(5 downto 0);
signal VN1644_sign_out : std_logic_vector(5 downto 0);
signal VN1645_data_out : std_logic_vector(5 downto 0);
signal VN1645_sign_out : std_logic_vector(5 downto 0);
signal VN1646_data_out : std_logic_vector(5 downto 0);
signal VN1646_sign_out : std_logic_vector(5 downto 0);
signal VN1647_data_out : std_logic_vector(5 downto 0);
signal VN1647_sign_out : std_logic_vector(5 downto 0);
signal VN1648_data_out : std_logic_vector(5 downto 0);
signal VN1648_sign_out : std_logic_vector(5 downto 0);
signal VN1649_data_out : std_logic_vector(5 downto 0);
signal VN1649_sign_out : std_logic_vector(5 downto 0);
signal VN1650_data_out : std_logic_vector(5 downto 0);
signal VN1650_sign_out : std_logic_vector(5 downto 0);
signal VN1651_data_out : std_logic_vector(5 downto 0);
signal VN1651_sign_out : std_logic_vector(5 downto 0);
signal VN1652_data_out : std_logic_vector(5 downto 0);
signal VN1652_sign_out : std_logic_vector(5 downto 0);
signal VN1653_data_out : std_logic_vector(5 downto 0);
signal VN1653_sign_out : std_logic_vector(5 downto 0);
signal VN1654_data_out : std_logic_vector(5 downto 0);
signal VN1654_sign_out : std_logic_vector(5 downto 0);
signal VN1655_data_out : std_logic_vector(5 downto 0);
signal VN1655_sign_out : std_logic_vector(5 downto 0);
signal VN1656_data_out : std_logic_vector(5 downto 0);
signal VN1656_sign_out : std_logic_vector(5 downto 0);
signal VN1657_data_out : std_logic_vector(5 downto 0);
signal VN1657_sign_out : std_logic_vector(5 downto 0);
signal VN1658_data_out : std_logic_vector(5 downto 0);
signal VN1658_sign_out : std_logic_vector(5 downto 0);
signal VN1659_data_out : std_logic_vector(5 downto 0);
signal VN1659_sign_out : std_logic_vector(5 downto 0);
signal VN1660_data_out : std_logic_vector(5 downto 0);
signal VN1660_sign_out : std_logic_vector(5 downto 0);
signal VN1661_data_out : std_logic_vector(5 downto 0);
signal VN1661_sign_out : std_logic_vector(5 downto 0);
signal VN1662_data_out : std_logic_vector(5 downto 0);
signal VN1662_sign_out : std_logic_vector(5 downto 0);
signal VN1663_data_out : std_logic_vector(5 downto 0);
signal VN1663_sign_out : std_logic_vector(5 downto 0);
signal VN1664_data_out : std_logic_vector(5 downto 0);
signal VN1664_sign_out : std_logic_vector(5 downto 0);
signal VN1665_data_out : std_logic_vector(5 downto 0);
signal VN1665_sign_out : std_logic_vector(5 downto 0);
signal VN1666_data_out : std_logic_vector(5 downto 0);
signal VN1666_sign_out : std_logic_vector(5 downto 0);
signal VN1667_data_out : std_logic_vector(5 downto 0);
signal VN1667_sign_out : std_logic_vector(5 downto 0);
signal VN1668_data_out : std_logic_vector(5 downto 0);
signal VN1668_sign_out : std_logic_vector(5 downto 0);
signal VN1669_data_out : std_logic_vector(5 downto 0);
signal VN1669_sign_out : std_logic_vector(5 downto 0);
signal VN1670_data_out : std_logic_vector(5 downto 0);
signal VN1670_sign_out : std_logic_vector(5 downto 0);
signal VN1671_data_out : std_logic_vector(5 downto 0);
signal VN1671_sign_out : std_logic_vector(5 downto 0);
signal VN1672_data_out : std_logic_vector(5 downto 0);
signal VN1672_sign_out : std_logic_vector(5 downto 0);
signal VN1673_data_out : std_logic_vector(5 downto 0);
signal VN1673_sign_out : std_logic_vector(5 downto 0);
signal VN1674_data_out : std_logic_vector(5 downto 0);
signal VN1674_sign_out : std_logic_vector(5 downto 0);
signal VN1675_data_out : std_logic_vector(5 downto 0);
signal VN1675_sign_out : std_logic_vector(5 downto 0);
signal VN1676_data_out : std_logic_vector(5 downto 0);
signal VN1676_sign_out : std_logic_vector(5 downto 0);
signal VN1677_data_out : std_logic_vector(5 downto 0);
signal VN1677_sign_out : std_logic_vector(5 downto 0);
signal VN1678_data_out : std_logic_vector(5 downto 0);
signal VN1678_sign_out : std_logic_vector(5 downto 0);
signal VN1679_data_out : std_logic_vector(5 downto 0);
signal VN1679_sign_out : std_logic_vector(5 downto 0);
signal VN1680_data_out : std_logic_vector(5 downto 0);
signal VN1680_sign_out : std_logic_vector(5 downto 0);
signal VN1681_data_out : std_logic_vector(5 downto 0);
signal VN1681_sign_out : std_logic_vector(5 downto 0);
signal VN1682_data_out : std_logic_vector(5 downto 0);
signal VN1682_sign_out : std_logic_vector(5 downto 0);
signal VN1683_data_out : std_logic_vector(5 downto 0);
signal VN1683_sign_out : std_logic_vector(5 downto 0);
signal VN1684_data_out : std_logic_vector(5 downto 0);
signal VN1684_sign_out : std_logic_vector(5 downto 0);
signal VN1685_data_out : std_logic_vector(5 downto 0);
signal VN1685_sign_out : std_logic_vector(5 downto 0);
signal VN1686_data_out : std_logic_vector(5 downto 0);
signal VN1686_sign_out : std_logic_vector(5 downto 0);
signal VN1687_data_out : std_logic_vector(5 downto 0);
signal VN1687_sign_out : std_logic_vector(5 downto 0);
signal VN1688_data_out : std_logic_vector(5 downto 0);
signal VN1688_sign_out : std_logic_vector(5 downto 0);
signal VN1689_data_out : std_logic_vector(5 downto 0);
signal VN1689_sign_out : std_logic_vector(5 downto 0);
signal VN1690_data_out : std_logic_vector(5 downto 0);
signal VN1690_sign_out : std_logic_vector(5 downto 0);
signal VN1691_data_out : std_logic_vector(5 downto 0);
signal VN1691_sign_out : std_logic_vector(5 downto 0);
signal VN1692_data_out : std_logic_vector(5 downto 0);
signal VN1692_sign_out : std_logic_vector(5 downto 0);
signal VN1693_data_out : std_logic_vector(5 downto 0);
signal VN1693_sign_out : std_logic_vector(5 downto 0);
signal VN1694_data_out : std_logic_vector(5 downto 0);
signal VN1694_sign_out : std_logic_vector(5 downto 0);
signal VN1695_data_out : std_logic_vector(5 downto 0);
signal VN1695_sign_out : std_logic_vector(5 downto 0);
signal VN1696_data_out : std_logic_vector(5 downto 0);
signal VN1696_sign_out : std_logic_vector(5 downto 0);
signal VN1697_data_out : std_logic_vector(5 downto 0);
signal VN1697_sign_out : std_logic_vector(5 downto 0);
signal VN1698_data_out : std_logic_vector(5 downto 0);
signal VN1698_sign_out : std_logic_vector(5 downto 0);
signal VN1699_data_out : std_logic_vector(5 downto 0);
signal VN1699_sign_out : std_logic_vector(5 downto 0);
signal VN1700_data_out : std_logic_vector(5 downto 0);
signal VN1700_sign_out : std_logic_vector(5 downto 0);
signal VN1701_data_out : std_logic_vector(5 downto 0);
signal VN1701_sign_out : std_logic_vector(5 downto 0);
signal VN1702_data_out : std_logic_vector(5 downto 0);
signal VN1702_sign_out : std_logic_vector(5 downto 0);
signal VN1703_data_out : std_logic_vector(5 downto 0);
signal VN1703_sign_out : std_logic_vector(5 downto 0);
signal VN1704_data_out : std_logic_vector(5 downto 0);
signal VN1704_sign_out : std_logic_vector(5 downto 0);
signal VN1705_data_out : std_logic_vector(5 downto 0);
signal VN1705_sign_out : std_logic_vector(5 downto 0);
signal VN1706_data_out : std_logic_vector(5 downto 0);
signal VN1706_sign_out : std_logic_vector(5 downto 0);
signal VN1707_data_out : std_logic_vector(5 downto 0);
signal VN1707_sign_out : std_logic_vector(5 downto 0);
signal VN1708_data_out : std_logic_vector(5 downto 0);
signal VN1708_sign_out : std_logic_vector(5 downto 0);
signal VN1709_data_out : std_logic_vector(5 downto 0);
signal VN1709_sign_out : std_logic_vector(5 downto 0);
signal VN1710_data_out : std_logic_vector(5 downto 0);
signal VN1710_sign_out : std_logic_vector(5 downto 0);
signal VN1711_data_out : std_logic_vector(5 downto 0);
signal VN1711_sign_out : std_logic_vector(5 downto 0);
signal VN1712_data_out : std_logic_vector(5 downto 0);
signal VN1712_sign_out : std_logic_vector(5 downto 0);
signal VN1713_data_out : std_logic_vector(5 downto 0);
signal VN1713_sign_out : std_logic_vector(5 downto 0);
signal VN1714_data_out : std_logic_vector(5 downto 0);
signal VN1714_sign_out : std_logic_vector(5 downto 0);
signal VN1715_data_out : std_logic_vector(5 downto 0);
signal VN1715_sign_out : std_logic_vector(5 downto 0);
signal VN1716_data_out : std_logic_vector(5 downto 0);
signal VN1716_sign_out : std_logic_vector(5 downto 0);
signal VN1717_data_out : std_logic_vector(5 downto 0);
signal VN1717_sign_out : std_logic_vector(5 downto 0);
signal VN1718_data_out : std_logic_vector(5 downto 0);
signal VN1718_sign_out : std_logic_vector(5 downto 0);
signal VN1719_data_out : std_logic_vector(5 downto 0);
signal VN1719_sign_out : std_logic_vector(5 downto 0);
signal VN1720_data_out : std_logic_vector(5 downto 0);
signal VN1720_sign_out : std_logic_vector(5 downto 0);
signal VN1721_data_out : std_logic_vector(5 downto 0);
signal VN1721_sign_out : std_logic_vector(5 downto 0);
signal VN1722_data_out : std_logic_vector(5 downto 0);
signal VN1722_sign_out : std_logic_vector(5 downto 0);
signal VN1723_data_out : std_logic_vector(5 downto 0);
signal VN1723_sign_out : std_logic_vector(5 downto 0);
signal VN1724_data_out : std_logic_vector(5 downto 0);
signal VN1724_sign_out : std_logic_vector(5 downto 0);
signal VN1725_data_out : std_logic_vector(5 downto 0);
signal VN1725_sign_out : std_logic_vector(5 downto 0);
signal VN1726_data_out : std_logic_vector(5 downto 0);
signal VN1726_sign_out : std_logic_vector(5 downto 0);
signal VN1727_data_out : std_logic_vector(5 downto 0);
signal VN1727_sign_out : std_logic_vector(5 downto 0);
signal VN1728_data_out : std_logic_vector(5 downto 0);
signal VN1728_sign_out : std_logic_vector(5 downto 0);
signal VN1729_data_out : std_logic_vector(5 downto 0);
signal VN1729_sign_out : std_logic_vector(5 downto 0);
signal VN1730_data_out : std_logic_vector(5 downto 0);
signal VN1730_sign_out : std_logic_vector(5 downto 0);
signal VN1731_data_out : std_logic_vector(5 downto 0);
signal VN1731_sign_out : std_logic_vector(5 downto 0);
signal VN1732_data_out : std_logic_vector(5 downto 0);
signal VN1732_sign_out : std_logic_vector(5 downto 0);
signal VN1733_data_out : std_logic_vector(5 downto 0);
signal VN1733_sign_out : std_logic_vector(5 downto 0);
signal VN1734_data_out : std_logic_vector(5 downto 0);
signal VN1734_sign_out : std_logic_vector(5 downto 0);
signal VN1735_data_out : std_logic_vector(5 downto 0);
signal VN1735_sign_out : std_logic_vector(5 downto 0);
signal VN1736_data_out : std_logic_vector(5 downto 0);
signal VN1736_sign_out : std_logic_vector(5 downto 0);
signal VN1737_data_out : std_logic_vector(5 downto 0);
signal VN1737_sign_out : std_logic_vector(5 downto 0);
signal VN1738_data_out : std_logic_vector(5 downto 0);
signal VN1738_sign_out : std_logic_vector(5 downto 0);
signal VN1739_data_out : std_logic_vector(5 downto 0);
signal VN1739_sign_out : std_logic_vector(5 downto 0);
signal VN1740_data_out : std_logic_vector(5 downto 0);
signal VN1740_sign_out : std_logic_vector(5 downto 0);
signal VN1741_data_out : std_logic_vector(5 downto 0);
signal VN1741_sign_out : std_logic_vector(5 downto 0);
signal VN1742_data_out : std_logic_vector(5 downto 0);
signal VN1742_sign_out : std_logic_vector(5 downto 0);
signal VN1743_data_out : std_logic_vector(5 downto 0);
signal VN1743_sign_out : std_logic_vector(5 downto 0);
signal VN1744_data_out : std_logic_vector(5 downto 0);
signal VN1744_sign_out : std_logic_vector(5 downto 0);
signal VN1745_data_out : std_logic_vector(5 downto 0);
signal VN1745_sign_out : std_logic_vector(5 downto 0);
signal VN1746_data_out : std_logic_vector(5 downto 0);
signal VN1746_sign_out : std_logic_vector(5 downto 0);
signal VN1747_data_out : std_logic_vector(5 downto 0);
signal VN1747_sign_out : std_logic_vector(5 downto 0);
signal VN1748_data_out : std_logic_vector(5 downto 0);
signal VN1748_sign_out : std_logic_vector(5 downto 0);
signal VN1749_data_out : std_logic_vector(5 downto 0);
signal VN1749_sign_out : std_logic_vector(5 downto 0);
signal VN1750_data_out : std_logic_vector(5 downto 0);
signal VN1750_sign_out : std_logic_vector(5 downto 0);
signal VN1751_data_out : std_logic_vector(5 downto 0);
signal VN1751_sign_out : std_logic_vector(5 downto 0);
signal VN1752_data_out : std_logic_vector(5 downto 0);
signal VN1752_sign_out : std_logic_vector(5 downto 0);
signal VN1753_data_out : std_logic_vector(5 downto 0);
signal VN1753_sign_out : std_logic_vector(5 downto 0);
signal VN1754_data_out : std_logic_vector(5 downto 0);
signal VN1754_sign_out : std_logic_vector(5 downto 0);
signal VN1755_data_out : std_logic_vector(5 downto 0);
signal VN1755_sign_out : std_logic_vector(5 downto 0);
signal VN1756_data_out : std_logic_vector(5 downto 0);
signal VN1756_sign_out : std_logic_vector(5 downto 0);
signal VN1757_data_out : std_logic_vector(5 downto 0);
signal VN1757_sign_out : std_logic_vector(5 downto 0);
signal VN1758_data_out : std_logic_vector(5 downto 0);
signal VN1758_sign_out : std_logic_vector(5 downto 0);
signal VN1759_data_out : std_logic_vector(5 downto 0);
signal VN1759_sign_out : std_logic_vector(5 downto 0);
signal VN1760_data_out : std_logic_vector(5 downto 0);
signal VN1760_sign_out : std_logic_vector(5 downto 0);
signal VN1761_data_out : std_logic_vector(5 downto 0);
signal VN1761_sign_out : std_logic_vector(5 downto 0);
signal VN1762_data_out : std_logic_vector(5 downto 0);
signal VN1762_sign_out : std_logic_vector(5 downto 0);
signal VN1763_data_out : std_logic_vector(5 downto 0);
signal VN1763_sign_out : std_logic_vector(5 downto 0);
signal VN1764_data_out : std_logic_vector(5 downto 0);
signal VN1764_sign_out : std_logic_vector(5 downto 0);
signal VN1765_data_out : std_logic_vector(5 downto 0);
signal VN1765_sign_out : std_logic_vector(5 downto 0);
signal VN1766_data_out : std_logic_vector(5 downto 0);
signal VN1766_sign_out : std_logic_vector(5 downto 0);
signal VN1767_data_out : std_logic_vector(5 downto 0);
signal VN1767_sign_out : std_logic_vector(5 downto 0);
signal VN1768_data_out : std_logic_vector(5 downto 0);
signal VN1768_sign_out : std_logic_vector(5 downto 0);
signal VN1769_data_out : std_logic_vector(5 downto 0);
signal VN1769_sign_out : std_logic_vector(5 downto 0);
signal VN1770_data_out : std_logic_vector(5 downto 0);
signal VN1770_sign_out : std_logic_vector(5 downto 0);
signal VN1771_data_out : std_logic_vector(5 downto 0);
signal VN1771_sign_out : std_logic_vector(5 downto 0);
signal VN1772_data_out : std_logic_vector(5 downto 0);
signal VN1772_sign_out : std_logic_vector(5 downto 0);
signal VN1773_data_out : std_logic_vector(5 downto 0);
signal VN1773_sign_out : std_logic_vector(5 downto 0);
signal VN1774_data_out : std_logic_vector(5 downto 0);
signal VN1774_sign_out : std_logic_vector(5 downto 0);
signal VN1775_data_out : std_logic_vector(5 downto 0);
signal VN1775_sign_out : std_logic_vector(5 downto 0);
signal VN1776_data_out : std_logic_vector(5 downto 0);
signal VN1776_sign_out : std_logic_vector(5 downto 0);
signal VN1777_data_out : std_logic_vector(5 downto 0);
signal VN1777_sign_out : std_logic_vector(5 downto 0);
signal VN1778_data_out : std_logic_vector(5 downto 0);
signal VN1778_sign_out : std_logic_vector(5 downto 0);
signal VN1779_data_out : std_logic_vector(5 downto 0);
signal VN1779_sign_out : std_logic_vector(5 downto 0);
signal VN1780_data_out : std_logic_vector(5 downto 0);
signal VN1780_sign_out : std_logic_vector(5 downto 0);
signal VN1781_data_out : std_logic_vector(5 downto 0);
signal VN1781_sign_out : std_logic_vector(5 downto 0);
signal VN1782_data_out : std_logic_vector(5 downto 0);
signal VN1782_sign_out : std_logic_vector(5 downto 0);
signal VN1783_data_out : std_logic_vector(5 downto 0);
signal VN1783_sign_out : std_logic_vector(5 downto 0);
signal VN1784_data_out : std_logic_vector(5 downto 0);
signal VN1784_sign_out : std_logic_vector(5 downto 0);
signal VN1785_data_out : std_logic_vector(5 downto 0);
signal VN1785_sign_out : std_logic_vector(5 downto 0);
signal VN1786_data_out : std_logic_vector(5 downto 0);
signal VN1786_sign_out : std_logic_vector(5 downto 0);
signal VN1787_data_out : std_logic_vector(5 downto 0);
signal VN1787_sign_out : std_logic_vector(5 downto 0);
signal VN1788_data_out : std_logic_vector(5 downto 0);
signal VN1788_sign_out : std_logic_vector(5 downto 0);
signal VN1789_data_out : std_logic_vector(5 downto 0);
signal VN1789_sign_out : std_logic_vector(5 downto 0);
signal VN1790_data_out : std_logic_vector(5 downto 0);
signal VN1790_sign_out : std_logic_vector(5 downto 0);
signal VN1791_data_out : std_logic_vector(5 downto 0);
signal VN1791_sign_out : std_logic_vector(5 downto 0);
signal VN1792_data_out : std_logic_vector(5 downto 0);
signal VN1792_sign_out : std_logic_vector(5 downto 0);
signal VN1793_data_out : std_logic_vector(5 downto 0);
signal VN1793_sign_out : std_logic_vector(5 downto 0);
signal VN1794_data_out : std_logic_vector(5 downto 0);
signal VN1794_sign_out : std_logic_vector(5 downto 0);
signal VN1795_data_out : std_logic_vector(5 downto 0);
signal VN1795_sign_out : std_logic_vector(5 downto 0);
signal VN1796_data_out : std_logic_vector(5 downto 0);
signal VN1796_sign_out : std_logic_vector(5 downto 0);
signal VN1797_data_out : std_logic_vector(5 downto 0);
signal VN1797_sign_out : std_logic_vector(5 downto 0);
signal VN1798_data_out : std_logic_vector(5 downto 0);
signal VN1798_sign_out : std_logic_vector(5 downto 0);
signal VN1799_data_out : std_logic_vector(5 downto 0);
signal VN1799_sign_out : std_logic_vector(5 downto 0);
signal VN1800_data_out : std_logic_vector(5 downto 0);
signal VN1800_sign_out : std_logic_vector(5 downto 0);
signal VN1801_data_out : std_logic_vector(5 downto 0);
signal VN1801_sign_out : std_logic_vector(5 downto 0);
signal VN1802_data_out : std_logic_vector(5 downto 0);
signal VN1802_sign_out : std_logic_vector(5 downto 0);
signal VN1803_data_out : std_logic_vector(5 downto 0);
signal VN1803_sign_out : std_logic_vector(5 downto 0);
signal VN1804_data_out : std_logic_vector(5 downto 0);
signal VN1804_sign_out : std_logic_vector(5 downto 0);
signal VN1805_data_out : std_logic_vector(5 downto 0);
signal VN1805_sign_out : std_logic_vector(5 downto 0);
signal VN1806_data_out : std_logic_vector(5 downto 0);
signal VN1806_sign_out : std_logic_vector(5 downto 0);
signal VN1807_data_out : std_logic_vector(5 downto 0);
signal VN1807_sign_out : std_logic_vector(5 downto 0);
signal VN1808_data_out : std_logic_vector(5 downto 0);
signal VN1808_sign_out : std_logic_vector(5 downto 0);
signal VN1809_data_out : std_logic_vector(5 downto 0);
signal VN1809_sign_out : std_logic_vector(5 downto 0);
signal VN1810_data_out : std_logic_vector(5 downto 0);
signal VN1810_sign_out : std_logic_vector(5 downto 0);
signal VN1811_data_out : std_logic_vector(5 downto 0);
signal VN1811_sign_out : std_logic_vector(5 downto 0);
signal VN1812_data_out : std_logic_vector(5 downto 0);
signal VN1812_sign_out : std_logic_vector(5 downto 0);
signal VN1813_data_out : std_logic_vector(5 downto 0);
signal VN1813_sign_out : std_logic_vector(5 downto 0);
signal VN1814_data_out : std_logic_vector(5 downto 0);
signal VN1814_sign_out : std_logic_vector(5 downto 0);
signal VN1815_data_out : std_logic_vector(5 downto 0);
signal VN1815_sign_out : std_logic_vector(5 downto 0);
signal VN1816_data_out : std_logic_vector(5 downto 0);
signal VN1816_sign_out : std_logic_vector(5 downto 0);
signal VN1817_data_out : std_logic_vector(5 downto 0);
signal VN1817_sign_out : std_logic_vector(5 downto 0);
signal VN1818_data_out : std_logic_vector(5 downto 0);
signal VN1818_sign_out : std_logic_vector(5 downto 0);
signal VN1819_data_out : std_logic_vector(5 downto 0);
signal VN1819_sign_out : std_logic_vector(5 downto 0);
signal VN1820_data_out : std_logic_vector(5 downto 0);
signal VN1820_sign_out : std_logic_vector(5 downto 0);
signal VN1821_data_out : std_logic_vector(5 downto 0);
signal VN1821_sign_out : std_logic_vector(5 downto 0);
signal VN1822_data_out : std_logic_vector(5 downto 0);
signal VN1822_sign_out : std_logic_vector(5 downto 0);
signal VN1823_data_out : std_logic_vector(5 downto 0);
signal VN1823_sign_out : std_logic_vector(5 downto 0);
signal VN1824_data_out : std_logic_vector(5 downto 0);
signal VN1824_sign_out : std_logic_vector(5 downto 0);
signal VN1825_data_out : std_logic_vector(5 downto 0);
signal VN1825_sign_out : std_logic_vector(5 downto 0);
signal VN1826_data_out : std_logic_vector(5 downto 0);
signal VN1826_sign_out : std_logic_vector(5 downto 0);
signal VN1827_data_out : std_logic_vector(5 downto 0);
signal VN1827_sign_out : std_logic_vector(5 downto 0);
signal VN1828_data_out : std_logic_vector(5 downto 0);
signal VN1828_sign_out : std_logic_vector(5 downto 0);
signal VN1829_data_out : std_logic_vector(5 downto 0);
signal VN1829_sign_out : std_logic_vector(5 downto 0);
signal VN1830_data_out : std_logic_vector(5 downto 0);
signal VN1830_sign_out : std_logic_vector(5 downto 0);
signal VN1831_data_out : std_logic_vector(5 downto 0);
signal VN1831_sign_out : std_logic_vector(5 downto 0);
signal VN1832_data_out : std_logic_vector(5 downto 0);
signal VN1832_sign_out : std_logic_vector(5 downto 0);
signal VN1833_data_out : std_logic_vector(5 downto 0);
signal VN1833_sign_out : std_logic_vector(5 downto 0);
signal VN1834_data_out : std_logic_vector(5 downto 0);
signal VN1834_sign_out : std_logic_vector(5 downto 0);
signal VN1835_data_out : std_logic_vector(5 downto 0);
signal VN1835_sign_out : std_logic_vector(5 downto 0);
signal VN1836_data_out : std_logic_vector(5 downto 0);
signal VN1836_sign_out : std_logic_vector(5 downto 0);
signal VN1837_data_out : std_logic_vector(5 downto 0);
signal VN1837_sign_out : std_logic_vector(5 downto 0);
signal VN1838_data_out : std_logic_vector(5 downto 0);
signal VN1838_sign_out : std_logic_vector(5 downto 0);
signal VN1839_data_out : std_logic_vector(5 downto 0);
signal VN1839_sign_out : std_logic_vector(5 downto 0);
signal VN1840_data_out : std_logic_vector(5 downto 0);
signal VN1840_sign_out : std_logic_vector(5 downto 0);
signal VN1841_data_out : std_logic_vector(5 downto 0);
signal VN1841_sign_out : std_logic_vector(5 downto 0);
signal VN1842_data_out : std_logic_vector(5 downto 0);
signal VN1842_sign_out : std_logic_vector(5 downto 0);
signal VN1843_data_out : std_logic_vector(5 downto 0);
signal VN1843_sign_out : std_logic_vector(5 downto 0);
signal VN1844_data_out : std_logic_vector(5 downto 0);
signal VN1844_sign_out : std_logic_vector(5 downto 0);
signal VN1845_data_out : std_logic_vector(5 downto 0);
signal VN1845_sign_out : std_logic_vector(5 downto 0);
signal VN1846_data_out : std_logic_vector(5 downto 0);
signal VN1846_sign_out : std_logic_vector(5 downto 0);
signal VN1847_data_out : std_logic_vector(5 downto 0);
signal VN1847_sign_out : std_logic_vector(5 downto 0);
signal VN1848_data_out : std_logic_vector(5 downto 0);
signal VN1848_sign_out : std_logic_vector(5 downto 0);
signal VN1849_data_out : std_logic_vector(5 downto 0);
signal VN1849_sign_out : std_logic_vector(5 downto 0);
signal VN1850_data_out : std_logic_vector(5 downto 0);
signal VN1850_sign_out : std_logic_vector(5 downto 0);
signal VN1851_data_out : std_logic_vector(5 downto 0);
signal VN1851_sign_out : std_logic_vector(5 downto 0);
signal VN1852_data_out : std_logic_vector(5 downto 0);
signal VN1852_sign_out : std_logic_vector(5 downto 0);
signal VN1853_data_out : std_logic_vector(5 downto 0);
signal VN1853_sign_out : std_logic_vector(5 downto 0);
signal VN1854_data_out : std_logic_vector(5 downto 0);
signal VN1854_sign_out : std_logic_vector(5 downto 0);
signal VN1855_data_out : std_logic_vector(5 downto 0);
signal VN1855_sign_out : std_logic_vector(5 downto 0);
signal VN1856_data_out : std_logic_vector(5 downto 0);
signal VN1856_sign_out : std_logic_vector(5 downto 0);
signal VN1857_data_out : std_logic_vector(5 downto 0);
signal VN1857_sign_out : std_logic_vector(5 downto 0);
signal VN1858_data_out : std_logic_vector(5 downto 0);
signal VN1858_sign_out : std_logic_vector(5 downto 0);
signal VN1859_data_out : std_logic_vector(5 downto 0);
signal VN1859_sign_out : std_logic_vector(5 downto 0);
signal VN1860_data_out : std_logic_vector(5 downto 0);
signal VN1860_sign_out : std_logic_vector(5 downto 0);
signal VN1861_data_out : std_logic_vector(5 downto 0);
signal VN1861_sign_out : std_logic_vector(5 downto 0);
signal VN1862_data_out : std_logic_vector(5 downto 0);
signal VN1862_sign_out : std_logic_vector(5 downto 0);
signal VN1863_data_out : std_logic_vector(5 downto 0);
signal VN1863_sign_out : std_logic_vector(5 downto 0);
signal VN1864_data_out : std_logic_vector(5 downto 0);
signal VN1864_sign_out : std_logic_vector(5 downto 0);
signal VN1865_data_out : std_logic_vector(5 downto 0);
signal VN1865_sign_out : std_logic_vector(5 downto 0);
signal VN1866_data_out : std_logic_vector(5 downto 0);
signal VN1866_sign_out : std_logic_vector(5 downto 0);
signal VN1867_data_out : std_logic_vector(5 downto 0);
signal VN1867_sign_out : std_logic_vector(5 downto 0);
signal VN1868_data_out : std_logic_vector(5 downto 0);
signal VN1868_sign_out : std_logic_vector(5 downto 0);
signal VN1869_data_out : std_logic_vector(5 downto 0);
signal VN1869_sign_out : std_logic_vector(5 downto 0);
signal VN1870_data_out : std_logic_vector(5 downto 0);
signal VN1870_sign_out : std_logic_vector(5 downto 0);
signal VN1871_data_out : std_logic_vector(5 downto 0);
signal VN1871_sign_out : std_logic_vector(5 downto 0);
signal VN1872_data_out : std_logic_vector(5 downto 0);
signal VN1872_sign_out : std_logic_vector(5 downto 0);
signal VN1873_data_out : std_logic_vector(5 downto 0);
signal VN1873_sign_out : std_logic_vector(5 downto 0);
signal VN1874_data_out : std_logic_vector(5 downto 0);
signal VN1874_sign_out : std_logic_vector(5 downto 0);
signal VN1875_data_out : std_logic_vector(5 downto 0);
signal VN1875_sign_out : std_logic_vector(5 downto 0);
signal VN1876_data_out : std_logic_vector(5 downto 0);
signal VN1876_sign_out : std_logic_vector(5 downto 0);
signal VN1877_data_out : std_logic_vector(5 downto 0);
signal VN1877_sign_out : std_logic_vector(5 downto 0);
signal VN1878_data_out : std_logic_vector(5 downto 0);
signal VN1878_sign_out : std_logic_vector(5 downto 0);
signal VN1879_data_out : std_logic_vector(5 downto 0);
signal VN1879_sign_out : std_logic_vector(5 downto 0);
signal VN1880_data_out : std_logic_vector(5 downto 0);
signal VN1880_sign_out : std_logic_vector(5 downto 0);
signal VN1881_data_out : std_logic_vector(5 downto 0);
signal VN1881_sign_out : std_logic_vector(5 downto 0);
signal VN1882_data_out : std_logic_vector(5 downto 0);
signal VN1882_sign_out : std_logic_vector(5 downto 0);
signal VN1883_data_out : std_logic_vector(5 downto 0);
signal VN1883_sign_out : std_logic_vector(5 downto 0);
signal VN1884_data_out : std_logic_vector(5 downto 0);
signal VN1884_sign_out : std_logic_vector(5 downto 0);
signal VN1885_data_out : std_logic_vector(5 downto 0);
signal VN1885_sign_out : std_logic_vector(5 downto 0);
signal VN1886_data_out : std_logic_vector(5 downto 0);
signal VN1886_sign_out : std_logic_vector(5 downto 0);
signal VN1887_data_out : std_logic_vector(5 downto 0);
signal VN1887_sign_out : std_logic_vector(5 downto 0);
signal VN1888_data_out : std_logic_vector(5 downto 0);
signal VN1888_sign_out : std_logic_vector(5 downto 0);
signal VN1889_data_out : std_logic_vector(5 downto 0);
signal VN1889_sign_out : std_logic_vector(5 downto 0);
signal VN1890_data_out : std_logic_vector(5 downto 0);
signal VN1890_sign_out : std_logic_vector(5 downto 0);
signal VN1891_data_out : std_logic_vector(5 downto 0);
signal VN1891_sign_out : std_logic_vector(5 downto 0);
signal VN1892_data_out : std_logic_vector(5 downto 0);
signal VN1892_sign_out : std_logic_vector(5 downto 0);
signal VN1893_data_out : std_logic_vector(5 downto 0);
signal VN1893_sign_out : std_logic_vector(5 downto 0);
signal VN1894_data_out : std_logic_vector(5 downto 0);
signal VN1894_sign_out : std_logic_vector(5 downto 0);
signal VN1895_data_out : std_logic_vector(5 downto 0);
signal VN1895_sign_out : std_logic_vector(5 downto 0);
signal VN1896_data_out : std_logic_vector(5 downto 0);
signal VN1896_sign_out : std_logic_vector(5 downto 0);
signal VN1897_data_out : std_logic_vector(5 downto 0);
signal VN1897_sign_out : std_logic_vector(5 downto 0);
signal VN1898_data_out : std_logic_vector(5 downto 0);
signal VN1898_sign_out : std_logic_vector(5 downto 0);
signal VN1899_data_out : std_logic_vector(5 downto 0);
signal VN1899_sign_out : std_logic_vector(5 downto 0);
signal VN1900_data_out : std_logic_vector(5 downto 0);
signal VN1900_sign_out : std_logic_vector(5 downto 0);
signal VN1901_data_out : std_logic_vector(5 downto 0);
signal VN1901_sign_out : std_logic_vector(5 downto 0);
signal VN1902_data_out : std_logic_vector(5 downto 0);
signal VN1902_sign_out : std_logic_vector(5 downto 0);
signal VN1903_data_out : std_logic_vector(5 downto 0);
signal VN1903_sign_out : std_logic_vector(5 downto 0);
signal VN1904_data_out : std_logic_vector(5 downto 0);
signal VN1904_sign_out : std_logic_vector(5 downto 0);
signal VN1905_data_out : std_logic_vector(5 downto 0);
signal VN1905_sign_out : std_logic_vector(5 downto 0);
signal VN1906_data_out : std_logic_vector(5 downto 0);
signal VN1906_sign_out : std_logic_vector(5 downto 0);
signal VN1907_data_out : std_logic_vector(5 downto 0);
signal VN1907_sign_out : std_logic_vector(5 downto 0);
signal VN1908_data_out : std_logic_vector(5 downto 0);
signal VN1908_sign_out : std_logic_vector(5 downto 0);
signal VN1909_data_out : std_logic_vector(5 downto 0);
signal VN1909_sign_out : std_logic_vector(5 downto 0);
signal VN1910_data_out : std_logic_vector(5 downto 0);
signal VN1910_sign_out : std_logic_vector(5 downto 0);
signal VN1911_data_out : std_logic_vector(5 downto 0);
signal VN1911_sign_out : std_logic_vector(5 downto 0);
signal VN1912_data_out : std_logic_vector(5 downto 0);
signal VN1912_sign_out : std_logic_vector(5 downto 0);
signal VN1913_data_out : std_logic_vector(5 downto 0);
signal VN1913_sign_out : std_logic_vector(5 downto 0);
signal VN1914_data_out : std_logic_vector(5 downto 0);
signal VN1914_sign_out : std_logic_vector(5 downto 0);
signal VN1915_data_out : std_logic_vector(5 downto 0);
signal VN1915_sign_out : std_logic_vector(5 downto 0);
signal VN1916_data_out : std_logic_vector(5 downto 0);
signal VN1916_sign_out : std_logic_vector(5 downto 0);
signal VN1917_data_out : std_logic_vector(5 downto 0);
signal VN1917_sign_out : std_logic_vector(5 downto 0);
signal VN1918_data_out : std_logic_vector(5 downto 0);
signal VN1918_sign_out : std_logic_vector(5 downto 0);
signal VN1919_data_out : std_logic_vector(5 downto 0);
signal VN1919_sign_out : std_logic_vector(5 downto 0);
signal VN1920_data_out : std_logic_vector(5 downto 0);
signal VN1920_sign_out : std_logic_vector(5 downto 0);
signal VN1921_data_out : std_logic_vector(5 downto 0);
signal VN1921_sign_out : std_logic_vector(5 downto 0);
signal VN1922_data_out : std_logic_vector(5 downto 0);
signal VN1922_sign_out : std_logic_vector(5 downto 0);
signal VN1923_data_out : std_logic_vector(5 downto 0);
signal VN1923_sign_out : std_logic_vector(5 downto 0);
signal VN1924_data_out : std_logic_vector(5 downto 0);
signal VN1924_sign_out : std_logic_vector(5 downto 0);
signal VN1925_data_out : std_logic_vector(5 downto 0);
signal VN1925_sign_out : std_logic_vector(5 downto 0);
signal VN1926_data_out : std_logic_vector(5 downto 0);
signal VN1926_sign_out : std_logic_vector(5 downto 0);
signal VN1927_data_out : std_logic_vector(5 downto 0);
signal VN1927_sign_out : std_logic_vector(5 downto 0);
signal VN1928_data_out : std_logic_vector(5 downto 0);
signal VN1928_sign_out : std_logic_vector(5 downto 0);
signal VN1929_data_out : std_logic_vector(5 downto 0);
signal VN1929_sign_out : std_logic_vector(5 downto 0);
signal VN1930_data_out : std_logic_vector(5 downto 0);
signal VN1930_sign_out : std_logic_vector(5 downto 0);
signal VN1931_data_out : std_logic_vector(5 downto 0);
signal VN1931_sign_out : std_logic_vector(5 downto 0);
signal VN1932_data_out : std_logic_vector(5 downto 0);
signal VN1932_sign_out : std_logic_vector(5 downto 0);
signal VN1933_data_out : std_logic_vector(5 downto 0);
signal VN1933_sign_out : std_logic_vector(5 downto 0);
signal VN1934_data_out : std_logic_vector(5 downto 0);
signal VN1934_sign_out : std_logic_vector(5 downto 0);
signal VN1935_data_out : std_logic_vector(5 downto 0);
signal VN1935_sign_out : std_logic_vector(5 downto 0);
signal VN1936_data_out : std_logic_vector(5 downto 0);
signal VN1936_sign_out : std_logic_vector(5 downto 0);
signal VN1937_data_out : std_logic_vector(5 downto 0);
signal VN1937_sign_out : std_logic_vector(5 downto 0);
signal VN1938_data_out : std_logic_vector(5 downto 0);
signal VN1938_sign_out : std_logic_vector(5 downto 0);
signal VN1939_data_out : std_logic_vector(5 downto 0);
signal VN1939_sign_out : std_logic_vector(5 downto 0);
signal VN1940_data_out : std_logic_vector(5 downto 0);
signal VN1940_sign_out : std_logic_vector(5 downto 0);
signal VN1941_data_out : std_logic_vector(5 downto 0);
signal VN1941_sign_out : std_logic_vector(5 downto 0);
signal VN1942_data_out : std_logic_vector(5 downto 0);
signal VN1942_sign_out : std_logic_vector(5 downto 0);
signal VN1943_data_out : std_logic_vector(5 downto 0);
signal VN1943_sign_out : std_logic_vector(5 downto 0);
signal VN1944_data_out : std_logic_vector(5 downto 0);
signal VN1944_sign_out : std_logic_vector(5 downto 0);
signal VN1945_data_out : std_logic_vector(5 downto 0);
signal VN1945_sign_out : std_logic_vector(5 downto 0);
signal VN1946_data_out : std_logic_vector(5 downto 0);
signal VN1946_sign_out : std_logic_vector(5 downto 0);
signal VN1947_data_out : std_logic_vector(5 downto 0);
signal VN1947_sign_out : std_logic_vector(5 downto 0);
signal VN1948_data_out : std_logic_vector(5 downto 0);
signal VN1948_sign_out : std_logic_vector(5 downto 0);
signal VN1949_data_out : std_logic_vector(5 downto 0);
signal VN1949_sign_out : std_logic_vector(5 downto 0);
signal VN1950_data_out : std_logic_vector(5 downto 0);
signal VN1950_sign_out : std_logic_vector(5 downto 0);
signal VN1951_data_out : std_logic_vector(5 downto 0);
signal VN1951_sign_out : std_logic_vector(5 downto 0);
signal VN1952_data_out : std_logic_vector(5 downto 0);
signal VN1952_sign_out : std_logic_vector(5 downto 0);
signal VN1953_data_out : std_logic_vector(5 downto 0);
signal VN1953_sign_out : std_logic_vector(5 downto 0);
signal VN1954_data_out : std_logic_vector(5 downto 0);
signal VN1954_sign_out : std_logic_vector(5 downto 0);
signal VN1955_data_out : std_logic_vector(5 downto 0);
signal VN1955_sign_out : std_logic_vector(5 downto 0);
signal VN1956_data_out : std_logic_vector(5 downto 0);
signal VN1956_sign_out : std_logic_vector(5 downto 0);
signal VN1957_data_out : std_logic_vector(5 downto 0);
signal VN1957_sign_out : std_logic_vector(5 downto 0);
signal VN1958_data_out : std_logic_vector(5 downto 0);
signal VN1958_sign_out : std_logic_vector(5 downto 0);
signal VN1959_data_out : std_logic_vector(5 downto 0);
signal VN1959_sign_out : std_logic_vector(5 downto 0);
signal VN1960_data_out : std_logic_vector(5 downto 0);
signal VN1960_sign_out : std_logic_vector(5 downto 0);
signal VN1961_data_out : std_logic_vector(5 downto 0);
signal VN1961_sign_out : std_logic_vector(5 downto 0);
signal VN1962_data_out : std_logic_vector(5 downto 0);
signal VN1962_sign_out : std_logic_vector(5 downto 0);
signal VN1963_data_out : std_logic_vector(5 downto 0);
signal VN1963_sign_out : std_logic_vector(5 downto 0);
signal VN1964_data_out : std_logic_vector(5 downto 0);
signal VN1964_sign_out : std_logic_vector(5 downto 0);
signal VN1965_data_out : std_logic_vector(5 downto 0);
signal VN1965_sign_out : std_logic_vector(5 downto 0);
signal VN1966_data_out : std_logic_vector(5 downto 0);
signal VN1966_sign_out : std_logic_vector(5 downto 0);
signal VN1967_data_out : std_logic_vector(5 downto 0);
signal VN1967_sign_out : std_logic_vector(5 downto 0);
signal VN1968_data_out : std_logic_vector(5 downto 0);
signal VN1968_sign_out : std_logic_vector(5 downto 0);
signal VN1969_data_out : std_logic_vector(5 downto 0);
signal VN1969_sign_out : std_logic_vector(5 downto 0);
signal VN1970_data_out : std_logic_vector(5 downto 0);
signal VN1970_sign_out : std_logic_vector(5 downto 0);
signal VN1971_data_out : std_logic_vector(5 downto 0);
signal VN1971_sign_out : std_logic_vector(5 downto 0);
signal VN1972_data_out : std_logic_vector(5 downto 0);
signal VN1972_sign_out : std_logic_vector(5 downto 0);
signal VN1973_data_out : std_logic_vector(5 downto 0);
signal VN1973_sign_out : std_logic_vector(5 downto 0);
signal VN1974_data_out : std_logic_vector(5 downto 0);
signal VN1974_sign_out : std_logic_vector(5 downto 0);
signal VN1975_data_out : std_logic_vector(5 downto 0);
signal VN1975_sign_out : std_logic_vector(5 downto 0);
signal VN1976_data_out : std_logic_vector(5 downto 0);
signal VN1976_sign_out : std_logic_vector(5 downto 0);
signal VN1977_data_out : std_logic_vector(5 downto 0);
signal VN1977_sign_out : std_logic_vector(5 downto 0);
signal VN1978_data_out : std_logic_vector(5 downto 0);
signal VN1978_sign_out : std_logic_vector(5 downto 0);
signal VN1979_data_out : std_logic_vector(5 downto 0);
signal VN1979_sign_out : std_logic_vector(5 downto 0);
signal VN1980_data_out : std_logic_vector(5 downto 0);
signal VN1980_sign_out : std_logic_vector(5 downto 0);
signal VN1981_data_out : std_logic_vector(5 downto 0);
signal VN1981_sign_out : std_logic_vector(5 downto 0);
signal VN1982_data_out : std_logic_vector(5 downto 0);
signal VN1982_sign_out : std_logic_vector(5 downto 0);
signal VN1983_data_out : std_logic_vector(5 downto 0);
signal VN1983_sign_out : std_logic_vector(5 downto 0);
signal VN1984_data_out : std_logic_vector(5 downto 0);
signal VN1984_sign_out : std_logic_vector(5 downto 0);
signal VN1985_data_out : std_logic_vector(5 downto 0);
signal VN1985_sign_out : std_logic_vector(5 downto 0);
signal VN1986_data_out : std_logic_vector(5 downto 0);
signal VN1986_sign_out : std_logic_vector(5 downto 0);
signal VN1987_data_out : std_logic_vector(5 downto 0);
signal VN1987_sign_out : std_logic_vector(5 downto 0);
signal VN1988_data_out : std_logic_vector(5 downto 0);
signal VN1988_sign_out : std_logic_vector(5 downto 0);
signal VN1989_data_out : std_logic_vector(5 downto 0);
signal VN1989_sign_out : std_logic_vector(5 downto 0);
signal VN1990_data_out : std_logic_vector(5 downto 0);
signal VN1990_sign_out : std_logic_vector(5 downto 0);
signal VN1991_data_out : std_logic_vector(5 downto 0);
signal VN1991_sign_out : std_logic_vector(5 downto 0);
signal VN1992_data_out : std_logic_vector(5 downto 0);
signal VN1992_sign_out : std_logic_vector(5 downto 0);
signal VN1993_data_out : std_logic_vector(5 downto 0);
signal VN1993_sign_out : std_logic_vector(5 downto 0);
signal VN1994_data_out : std_logic_vector(5 downto 0);
signal VN1994_sign_out : std_logic_vector(5 downto 0);
signal VN1995_data_out : std_logic_vector(5 downto 0);
signal VN1995_sign_out : std_logic_vector(5 downto 0);
signal VN1996_data_out : std_logic_vector(5 downto 0);
signal VN1996_sign_out : std_logic_vector(5 downto 0);
signal VN1997_data_out : std_logic_vector(5 downto 0);
signal VN1997_sign_out : std_logic_vector(5 downto 0);
signal VN1998_data_out : std_logic_vector(5 downto 0);
signal VN1998_sign_out : std_logic_vector(5 downto 0);
signal VN1999_data_out : std_logic_vector(5 downto 0);
signal VN1999_sign_out : std_logic_vector(5 downto 0);
signal VN2000_data_out : std_logic_vector(5 downto 0);
signal VN2000_sign_out : std_logic_vector(5 downto 0);
signal VN2001_data_out : std_logic_vector(5 downto 0);
signal VN2001_sign_out : std_logic_vector(5 downto 0);
signal VN2002_data_out : std_logic_vector(5 downto 0);
signal VN2002_sign_out : std_logic_vector(5 downto 0);
signal VN2003_data_out : std_logic_vector(5 downto 0);
signal VN2003_sign_out : std_logic_vector(5 downto 0);
signal VN2004_data_out : std_logic_vector(5 downto 0);
signal VN2004_sign_out : std_logic_vector(5 downto 0);
signal VN2005_data_out : std_logic_vector(5 downto 0);
signal VN2005_sign_out : std_logic_vector(5 downto 0);
signal VN2006_data_out : std_logic_vector(5 downto 0);
signal VN2006_sign_out : std_logic_vector(5 downto 0);
signal VN2007_data_out : std_logic_vector(5 downto 0);
signal VN2007_sign_out : std_logic_vector(5 downto 0);
signal VN2008_data_out : std_logic_vector(5 downto 0);
signal VN2008_sign_out : std_logic_vector(5 downto 0);
signal VN2009_data_out : std_logic_vector(5 downto 0);
signal VN2009_sign_out : std_logic_vector(5 downto 0);
signal VN2010_data_out : std_logic_vector(5 downto 0);
signal VN2010_sign_out : std_logic_vector(5 downto 0);
signal VN2011_data_out : std_logic_vector(5 downto 0);
signal VN2011_sign_out : std_logic_vector(5 downto 0);
signal VN2012_data_out : std_logic_vector(5 downto 0);
signal VN2012_sign_out : std_logic_vector(5 downto 0);
signal VN2013_data_out : std_logic_vector(5 downto 0);
signal VN2013_sign_out : std_logic_vector(5 downto 0);
signal VN2014_data_out : std_logic_vector(5 downto 0);
signal VN2014_sign_out : std_logic_vector(5 downto 0);
signal VN2015_data_out : std_logic_vector(5 downto 0);
signal VN2015_sign_out : std_logic_vector(5 downto 0);
signal VN2016_data_out : std_logic_vector(5 downto 0);
signal VN2016_sign_out : std_logic_vector(5 downto 0);
signal VN2017_data_out : std_logic_vector(5 downto 0);
signal VN2017_sign_out : std_logic_vector(5 downto 0);
signal VN2018_data_out : std_logic_vector(5 downto 0);
signal VN2018_sign_out : std_logic_vector(5 downto 0);
signal VN2019_data_out : std_logic_vector(5 downto 0);
signal VN2019_sign_out : std_logic_vector(5 downto 0);
signal VN2020_data_out : std_logic_vector(5 downto 0);
signal VN2020_sign_out : std_logic_vector(5 downto 0);
signal VN2021_data_out : std_logic_vector(5 downto 0);
signal VN2021_sign_out : std_logic_vector(5 downto 0);
signal VN2022_data_out : std_logic_vector(5 downto 0);
signal VN2022_sign_out : std_logic_vector(5 downto 0);
signal VN2023_data_out : std_logic_vector(5 downto 0);
signal VN2023_sign_out : std_logic_vector(5 downto 0);
signal VN2024_data_out : std_logic_vector(5 downto 0);
signal VN2024_sign_out : std_logic_vector(5 downto 0);
signal VN2025_data_out : std_logic_vector(5 downto 0);
signal VN2025_sign_out : std_logic_vector(5 downto 0);
signal VN2026_data_out : std_logic_vector(5 downto 0);
signal VN2026_sign_out : std_logic_vector(5 downto 0);
signal VN2027_data_out : std_logic_vector(5 downto 0);
signal VN2027_sign_out : std_logic_vector(5 downto 0);
signal VN2028_data_out : std_logic_vector(5 downto 0);
signal VN2028_sign_out : std_logic_vector(5 downto 0);
signal VN2029_data_out : std_logic_vector(5 downto 0);
signal VN2029_sign_out : std_logic_vector(5 downto 0);
signal VN2030_data_out : std_logic_vector(5 downto 0);
signal VN2030_sign_out : std_logic_vector(5 downto 0);
signal VN2031_data_out : std_logic_vector(5 downto 0);
signal VN2031_sign_out : std_logic_vector(5 downto 0);
signal VN2032_data_out : std_logic_vector(5 downto 0);
signal VN2032_sign_out : std_logic_vector(5 downto 0);
signal VN2033_data_out : std_logic_vector(5 downto 0);
signal VN2033_sign_out : std_logic_vector(5 downto 0);
signal VN2034_data_out : std_logic_vector(5 downto 0);
signal VN2034_sign_out : std_logic_vector(5 downto 0);
signal VN2035_data_out : std_logic_vector(5 downto 0);
signal VN2035_sign_out : std_logic_vector(5 downto 0);
signal VN2036_data_out : std_logic_vector(5 downto 0);
signal VN2036_sign_out : std_logic_vector(5 downto 0);
signal VN2037_data_out : std_logic_vector(5 downto 0);
signal VN2037_sign_out : std_logic_vector(5 downto 0);
signal VN2038_data_out : std_logic_vector(5 downto 0);
signal VN2038_sign_out : std_logic_vector(5 downto 0);
signal VN2039_data_out : std_logic_vector(5 downto 0);
signal VN2039_sign_out : std_logic_vector(5 downto 0);
signal VN2040_data_out : std_logic_vector(5 downto 0);
signal VN2040_sign_out : std_logic_vector(5 downto 0);
signal VN2041_data_out : std_logic_vector(5 downto 0);
signal VN2041_sign_out : std_logic_vector(5 downto 0);
signal VN2042_data_out : std_logic_vector(5 downto 0);
signal VN2042_sign_out : std_logic_vector(5 downto 0);
signal VN2043_data_out : std_logic_vector(5 downto 0);
signal VN2043_sign_out : std_logic_vector(5 downto 0);
signal VN2044_data_out : std_logic_vector(5 downto 0);
signal VN2044_sign_out : std_logic_vector(5 downto 0);
signal VN2045_data_out : std_logic_vector(5 downto 0);
signal VN2045_sign_out : std_logic_vector(5 downto 0);
signal VN2046_data_out : std_logic_vector(5 downto 0);
signal VN2046_sign_out : std_logic_vector(5 downto 0);
signal VN2047_data_out : std_logic_vector(5 downto 0);
signal VN2047_sign_out : std_logic_vector(5 downto 0);
begin

    CN_data_in( 31 downto 0) <= CN0_data_in;
    CN_sign_in( 31 downto 0) <= CN0_sign_in;
    CN_data_in( 63 downto 32) <= CN1_data_in;
    CN_sign_in( 63 downto 32) <= CN1_sign_in;
    CN_data_in( 95 downto 64) <= CN2_data_in;
    CN_sign_in( 95 downto 64) <= CN2_sign_in;
    CN_data_in( 127 downto 96) <= CN3_data_in;
    CN_sign_in( 127 downto 96) <= CN3_sign_in;
    CN_data_in( 159 downto 128) <= CN4_data_in;
    CN_sign_in( 159 downto 128) <= CN4_sign_in;
    CN_data_in( 191 downto 160) <= CN5_data_in;
    CN_sign_in( 191 downto 160) <= CN5_sign_in;
    CN_data_in( 223 downto 192) <= CN6_data_in;
    CN_sign_in( 223 downto 192) <= CN6_sign_in;
    CN_data_in( 255 downto 224) <= CN7_data_in;
    CN_sign_in( 255 downto 224) <= CN7_sign_in;
    CN_data_in( 287 downto 256) <= CN8_data_in;
    CN_sign_in( 287 downto 256) <= CN8_sign_in;
    CN_data_in( 319 downto 288) <= CN9_data_in;
    CN_sign_in( 319 downto 288) <= CN9_sign_in;
    CN_data_in( 351 downto 320) <= CN10_data_in;
    CN_sign_in( 351 downto 320) <= CN10_sign_in;
    CN_data_in( 383 downto 352) <= CN11_data_in;
    CN_sign_in( 383 downto 352) <= CN11_sign_in;
    CN_data_in( 415 downto 384) <= CN12_data_in;
    CN_sign_in( 415 downto 384) <= CN12_sign_in;
    CN_data_in( 447 downto 416) <= CN13_data_in;
    CN_sign_in( 447 downto 416) <= CN13_sign_in;
    CN_data_in( 479 downto 448) <= CN14_data_in;
    CN_sign_in( 479 downto 448) <= CN14_sign_in;
    CN_data_in( 511 downto 480) <= CN15_data_in;
    CN_sign_in( 511 downto 480) <= CN15_sign_in;
    CN_data_in( 543 downto 512) <= CN16_data_in;
    CN_sign_in( 543 downto 512) <= CN16_sign_in;
    CN_data_in( 575 downto 544) <= CN17_data_in;
    CN_sign_in( 575 downto 544) <= CN17_sign_in;
    CN_data_in( 607 downto 576) <= CN18_data_in;
    CN_sign_in( 607 downto 576) <= CN18_sign_in;
    CN_data_in( 639 downto 608) <= CN19_data_in;
    CN_sign_in( 639 downto 608) <= CN19_sign_in;
    CN_data_in( 671 downto 640) <= CN20_data_in;
    CN_sign_in( 671 downto 640) <= CN20_sign_in;
    CN_data_in( 703 downto 672) <= CN21_data_in;
    CN_sign_in( 703 downto 672) <= CN21_sign_in;
    CN_data_in( 735 downto 704) <= CN22_data_in;
    CN_sign_in( 735 downto 704) <= CN22_sign_in;
    CN_data_in( 767 downto 736) <= CN23_data_in;
    CN_sign_in( 767 downto 736) <= CN23_sign_in;
    CN_data_in( 799 downto 768) <= CN24_data_in;
    CN_sign_in( 799 downto 768) <= CN24_sign_in;
    CN_data_in( 831 downto 800) <= CN25_data_in;
    CN_sign_in( 831 downto 800) <= CN25_sign_in;
    CN_data_in( 863 downto 832) <= CN26_data_in;
    CN_sign_in( 863 downto 832) <= CN26_sign_in;
    CN_data_in( 895 downto 864) <= CN27_data_in;
    CN_sign_in( 895 downto 864) <= CN27_sign_in;
    CN_data_in( 927 downto 896) <= CN28_data_in;
    CN_sign_in( 927 downto 896) <= CN28_sign_in;
    CN_data_in( 959 downto 928) <= CN29_data_in;
    CN_sign_in( 959 downto 928) <= CN29_sign_in;
    CN_data_in( 991 downto 960) <= CN30_data_in;
    CN_sign_in( 991 downto 960) <= CN30_sign_in;
    CN_data_in( 1023 downto 992) <= CN31_data_in;
    CN_sign_in( 1023 downto 992) <= CN31_sign_in;
    CN_data_in( 1055 downto 1024) <= CN32_data_in;
    CN_sign_in( 1055 downto 1024) <= CN32_sign_in;
    CN_data_in( 1087 downto 1056) <= CN33_data_in;
    CN_sign_in( 1087 downto 1056) <= CN33_sign_in;
    CN_data_in( 1119 downto 1088) <= CN34_data_in;
    CN_sign_in( 1119 downto 1088) <= CN34_sign_in;
    CN_data_in( 1151 downto 1120) <= CN35_data_in;
    CN_sign_in( 1151 downto 1120) <= CN35_sign_in;
    CN_data_in( 1183 downto 1152) <= CN36_data_in;
    CN_sign_in( 1183 downto 1152) <= CN36_sign_in;
    CN_data_in( 1215 downto 1184) <= CN37_data_in;
    CN_sign_in( 1215 downto 1184) <= CN37_sign_in;
    CN_data_in( 1247 downto 1216) <= CN38_data_in;
    CN_sign_in( 1247 downto 1216) <= CN38_sign_in;
    CN_data_in( 1279 downto 1248) <= CN39_data_in;
    CN_sign_in( 1279 downto 1248) <= CN39_sign_in;
    CN_data_in( 1311 downto 1280) <= CN40_data_in;
    CN_sign_in( 1311 downto 1280) <= CN40_sign_in;
    CN_data_in( 1343 downto 1312) <= CN41_data_in;
    CN_sign_in( 1343 downto 1312) <= CN41_sign_in;
    CN_data_in( 1375 downto 1344) <= CN42_data_in;
    CN_sign_in( 1375 downto 1344) <= CN42_sign_in;
    CN_data_in( 1407 downto 1376) <= CN43_data_in;
    CN_sign_in( 1407 downto 1376) <= CN43_sign_in;
    CN_data_in( 1439 downto 1408) <= CN44_data_in;
    CN_sign_in( 1439 downto 1408) <= CN44_sign_in;
    CN_data_in( 1471 downto 1440) <= CN45_data_in;
    CN_sign_in( 1471 downto 1440) <= CN45_sign_in;
    CN_data_in( 1503 downto 1472) <= CN46_data_in;
    CN_sign_in( 1503 downto 1472) <= CN46_sign_in;
    CN_data_in( 1535 downto 1504) <= CN47_data_in;
    CN_sign_in( 1535 downto 1504) <= CN47_sign_in;
    CN_data_in( 1567 downto 1536) <= CN48_data_in;
    CN_sign_in( 1567 downto 1536) <= CN48_sign_in;
    CN_data_in( 1599 downto 1568) <= CN49_data_in;
    CN_sign_in( 1599 downto 1568) <= CN49_sign_in;
    CN_data_in( 1631 downto 1600) <= CN50_data_in;
    CN_sign_in( 1631 downto 1600) <= CN50_sign_in;
    CN_data_in( 1663 downto 1632) <= CN51_data_in;
    CN_sign_in( 1663 downto 1632) <= CN51_sign_in;
    CN_data_in( 1695 downto 1664) <= CN52_data_in;
    CN_sign_in( 1695 downto 1664) <= CN52_sign_in;
    CN_data_in( 1727 downto 1696) <= CN53_data_in;
    CN_sign_in( 1727 downto 1696) <= CN53_sign_in;
    CN_data_in( 1759 downto 1728) <= CN54_data_in;
    CN_sign_in( 1759 downto 1728) <= CN54_sign_in;
    CN_data_in( 1791 downto 1760) <= CN55_data_in;
    CN_sign_in( 1791 downto 1760) <= CN55_sign_in;
    CN_data_in( 1823 downto 1792) <= CN56_data_in;
    CN_sign_in( 1823 downto 1792) <= CN56_sign_in;
    CN_data_in( 1855 downto 1824) <= CN57_data_in;
    CN_sign_in( 1855 downto 1824) <= CN57_sign_in;
    CN_data_in( 1887 downto 1856) <= CN58_data_in;
    CN_sign_in( 1887 downto 1856) <= CN58_sign_in;
    CN_data_in( 1919 downto 1888) <= CN59_data_in;
    CN_sign_in( 1919 downto 1888) <= CN59_sign_in;
    CN_data_in( 1951 downto 1920) <= CN60_data_in;
    CN_sign_in( 1951 downto 1920) <= CN60_sign_in;
    CN_data_in( 1983 downto 1952) <= CN61_data_in;
    CN_sign_in( 1983 downto 1952) <= CN61_sign_in;
    CN_data_in( 2015 downto 1984) <= CN62_data_in;
    CN_sign_in( 2015 downto 1984) <= CN62_sign_in;
    CN_data_in( 2047 downto 2016) <= CN63_data_in;
    CN_sign_in( 2047 downto 2016) <= CN63_sign_in;
    CN_data_in( 2079 downto 2048) <= CN64_data_in;
    CN_sign_in( 2079 downto 2048) <= CN64_sign_in;
    CN_data_in( 2111 downto 2080) <= CN65_data_in;
    CN_sign_in( 2111 downto 2080) <= CN65_sign_in;
    CN_data_in( 2143 downto 2112) <= CN66_data_in;
    CN_sign_in( 2143 downto 2112) <= CN66_sign_in;
    CN_data_in( 2175 downto 2144) <= CN67_data_in;
    CN_sign_in( 2175 downto 2144) <= CN67_sign_in;
    CN_data_in( 2207 downto 2176) <= CN68_data_in;
    CN_sign_in( 2207 downto 2176) <= CN68_sign_in;
    CN_data_in( 2239 downto 2208) <= CN69_data_in;
    CN_sign_in( 2239 downto 2208) <= CN69_sign_in;
    CN_data_in( 2271 downto 2240) <= CN70_data_in;
    CN_sign_in( 2271 downto 2240) <= CN70_sign_in;
    CN_data_in( 2303 downto 2272) <= CN71_data_in;
    CN_sign_in( 2303 downto 2272) <= CN71_sign_in;
    CN_data_in( 2335 downto 2304) <= CN72_data_in;
    CN_sign_in( 2335 downto 2304) <= CN72_sign_in;
    CN_data_in( 2367 downto 2336) <= CN73_data_in;
    CN_sign_in( 2367 downto 2336) <= CN73_sign_in;
    CN_data_in( 2399 downto 2368) <= CN74_data_in;
    CN_sign_in( 2399 downto 2368) <= CN74_sign_in;
    CN_data_in( 2431 downto 2400) <= CN75_data_in;
    CN_sign_in( 2431 downto 2400) <= CN75_sign_in;
    CN_data_in( 2463 downto 2432) <= CN76_data_in;
    CN_sign_in( 2463 downto 2432) <= CN76_sign_in;
    CN_data_in( 2495 downto 2464) <= CN77_data_in;
    CN_sign_in( 2495 downto 2464) <= CN77_sign_in;
    CN_data_in( 2527 downto 2496) <= CN78_data_in;
    CN_sign_in( 2527 downto 2496) <= CN78_sign_in;
    CN_data_in( 2559 downto 2528) <= CN79_data_in;
    CN_sign_in( 2559 downto 2528) <= CN79_sign_in;
    CN_data_in( 2591 downto 2560) <= CN80_data_in;
    CN_sign_in( 2591 downto 2560) <= CN80_sign_in;
    CN_data_in( 2623 downto 2592) <= CN81_data_in;
    CN_sign_in( 2623 downto 2592) <= CN81_sign_in;
    CN_data_in( 2655 downto 2624) <= CN82_data_in;
    CN_sign_in( 2655 downto 2624) <= CN82_sign_in;
    CN_data_in( 2687 downto 2656) <= CN83_data_in;
    CN_sign_in( 2687 downto 2656) <= CN83_sign_in;
    CN_data_in( 2719 downto 2688) <= CN84_data_in;
    CN_sign_in( 2719 downto 2688) <= CN84_sign_in;
    CN_data_in( 2751 downto 2720) <= CN85_data_in;
    CN_sign_in( 2751 downto 2720) <= CN85_sign_in;
    CN_data_in( 2783 downto 2752) <= CN86_data_in;
    CN_sign_in( 2783 downto 2752) <= CN86_sign_in;
    CN_data_in( 2815 downto 2784) <= CN87_data_in;
    CN_sign_in( 2815 downto 2784) <= CN87_sign_in;
    CN_data_in( 2847 downto 2816) <= CN88_data_in;
    CN_sign_in( 2847 downto 2816) <= CN88_sign_in;
    CN_data_in( 2879 downto 2848) <= CN89_data_in;
    CN_sign_in( 2879 downto 2848) <= CN89_sign_in;
    CN_data_in( 2911 downto 2880) <= CN90_data_in;
    CN_sign_in( 2911 downto 2880) <= CN90_sign_in;
    CN_data_in( 2943 downto 2912) <= CN91_data_in;
    CN_sign_in( 2943 downto 2912) <= CN91_sign_in;
    CN_data_in( 2975 downto 2944) <= CN92_data_in;
    CN_sign_in( 2975 downto 2944) <= CN92_sign_in;
    CN_data_in( 3007 downto 2976) <= CN93_data_in;
    CN_sign_in( 3007 downto 2976) <= CN93_sign_in;
    CN_data_in( 3039 downto 3008) <= CN94_data_in;
    CN_sign_in( 3039 downto 3008) <= CN94_sign_in;
    CN_data_in( 3071 downto 3040) <= CN95_data_in;
    CN_sign_in( 3071 downto 3040) <= CN95_sign_in;
    CN_data_in( 3103 downto 3072) <= CN96_data_in;
    CN_sign_in( 3103 downto 3072) <= CN96_sign_in;
    CN_data_in( 3135 downto 3104) <= CN97_data_in;
    CN_sign_in( 3135 downto 3104) <= CN97_sign_in;
    CN_data_in( 3167 downto 3136) <= CN98_data_in;
    CN_sign_in( 3167 downto 3136) <= CN98_sign_in;
    CN_data_in( 3199 downto 3168) <= CN99_data_in;
    CN_sign_in( 3199 downto 3168) <= CN99_sign_in;
    CN_data_in( 3231 downto 3200) <= CN100_data_in;
    CN_sign_in( 3231 downto 3200) <= CN100_sign_in;
    CN_data_in( 3263 downto 3232) <= CN101_data_in;
    CN_sign_in( 3263 downto 3232) <= CN101_sign_in;
    CN_data_in( 3295 downto 3264) <= CN102_data_in;
    CN_sign_in( 3295 downto 3264) <= CN102_sign_in;
    CN_data_in( 3327 downto 3296) <= CN103_data_in;
    CN_sign_in( 3327 downto 3296) <= CN103_sign_in;
    CN_data_in( 3359 downto 3328) <= CN104_data_in;
    CN_sign_in( 3359 downto 3328) <= CN104_sign_in;
    CN_data_in( 3391 downto 3360) <= CN105_data_in;
    CN_sign_in( 3391 downto 3360) <= CN105_sign_in;
    CN_data_in( 3423 downto 3392) <= CN106_data_in;
    CN_sign_in( 3423 downto 3392) <= CN106_sign_in;
    CN_data_in( 3455 downto 3424) <= CN107_data_in;
    CN_sign_in( 3455 downto 3424) <= CN107_sign_in;
    CN_data_in( 3487 downto 3456) <= CN108_data_in;
    CN_sign_in( 3487 downto 3456) <= CN108_sign_in;
    CN_data_in( 3519 downto 3488) <= CN109_data_in;
    CN_sign_in( 3519 downto 3488) <= CN109_sign_in;
    CN_data_in( 3551 downto 3520) <= CN110_data_in;
    CN_sign_in( 3551 downto 3520) <= CN110_sign_in;
    CN_data_in( 3583 downto 3552) <= CN111_data_in;
    CN_sign_in( 3583 downto 3552) <= CN111_sign_in;
    CN_data_in( 3615 downto 3584) <= CN112_data_in;
    CN_sign_in( 3615 downto 3584) <= CN112_sign_in;
    CN_data_in( 3647 downto 3616) <= CN113_data_in;
    CN_sign_in( 3647 downto 3616) <= CN113_sign_in;
    CN_data_in( 3679 downto 3648) <= CN114_data_in;
    CN_sign_in( 3679 downto 3648) <= CN114_sign_in;
    CN_data_in( 3711 downto 3680) <= CN115_data_in;
    CN_sign_in( 3711 downto 3680) <= CN115_sign_in;
    CN_data_in( 3743 downto 3712) <= CN116_data_in;
    CN_sign_in( 3743 downto 3712) <= CN116_sign_in;
    CN_data_in( 3775 downto 3744) <= CN117_data_in;
    CN_sign_in( 3775 downto 3744) <= CN117_sign_in;
    CN_data_in( 3807 downto 3776) <= CN118_data_in;
    CN_sign_in( 3807 downto 3776) <= CN118_sign_in;
    CN_data_in( 3839 downto 3808) <= CN119_data_in;
    CN_sign_in( 3839 downto 3808) <= CN119_sign_in;
    CN_data_in( 3871 downto 3840) <= CN120_data_in;
    CN_sign_in( 3871 downto 3840) <= CN120_sign_in;
    CN_data_in( 3903 downto 3872) <= CN121_data_in;
    CN_sign_in( 3903 downto 3872) <= CN121_sign_in;
    CN_data_in( 3935 downto 3904) <= CN122_data_in;
    CN_sign_in( 3935 downto 3904) <= CN122_sign_in;
    CN_data_in( 3967 downto 3936) <= CN123_data_in;
    CN_sign_in( 3967 downto 3936) <= CN123_sign_in;
    CN_data_in( 3999 downto 3968) <= CN124_data_in;
    CN_sign_in( 3999 downto 3968) <= CN124_sign_in;
    CN_data_in( 4031 downto 4000) <= CN125_data_in;
    CN_sign_in( 4031 downto 4000) <= CN125_sign_in;
    CN_data_in( 4063 downto 4032) <= CN126_data_in;
    CN_sign_in( 4063 downto 4032) <= CN126_sign_in;
    CN_data_in( 4095 downto 4064) <= CN127_data_in;
    CN_sign_in( 4095 downto 4064) <= CN127_sign_in;
    CN_data_in( 4127 downto 4096) <= CN128_data_in;
    CN_sign_in( 4127 downto 4096) <= CN128_sign_in;
    CN_data_in( 4159 downto 4128) <= CN129_data_in;
    CN_sign_in( 4159 downto 4128) <= CN129_sign_in;
    CN_data_in( 4191 downto 4160) <= CN130_data_in;
    CN_sign_in( 4191 downto 4160) <= CN130_sign_in;
    CN_data_in( 4223 downto 4192) <= CN131_data_in;
    CN_sign_in( 4223 downto 4192) <= CN131_sign_in;
    CN_data_in( 4255 downto 4224) <= CN132_data_in;
    CN_sign_in( 4255 downto 4224) <= CN132_sign_in;
    CN_data_in( 4287 downto 4256) <= CN133_data_in;
    CN_sign_in( 4287 downto 4256) <= CN133_sign_in;
    CN_data_in( 4319 downto 4288) <= CN134_data_in;
    CN_sign_in( 4319 downto 4288) <= CN134_sign_in;
    CN_data_in( 4351 downto 4320) <= CN135_data_in;
    CN_sign_in( 4351 downto 4320) <= CN135_sign_in;
    CN_data_in( 4383 downto 4352) <= CN136_data_in;
    CN_sign_in( 4383 downto 4352) <= CN136_sign_in;
    CN_data_in( 4415 downto 4384) <= CN137_data_in;
    CN_sign_in( 4415 downto 4384) <= CN137_sign_in;
    CN_data_in( 4447 downto 4416) <= CN138_data_in;
    CN_sign_in( 4447 downto 4416) <= CN138_sign_in;
    CN_data_in( 4479 downto 4448) <= CN139_data_in;
    CN_sign_in( 4479 downto 4448) <= CN139_sign_in;
    CN_data_in( 4511 downto 4480) <= CN140_data_in;
    CN_sign_in( 4511 downto 4480) <= CN140_sign_in;
    CN_data_in( 4543 downto 4512) <= CN141_data_in;
    CN_sign_in( 4543 downto 4512) <= CN141_sign_in;
    CN_data_in( 4575 downto 4544) <= CN142_data_in;
    CN_sign_in( 4575 downto 4544) <= CN142_sign_in;
    CN_data_in( 4607 downto 4576) <= CN143_data_in;
    CN_sign_in( 4607 downto 4576) <= CN143_sign_in;
    CN_data_in( 4639 downto 4608) <= CN144_data_in;
    CN_sign_in( 4639 downto 4608) <= CN144_sign_in;
    CN_data_in( 4671 downto 4640) <= CN145_data_in;
    CN_sign_in( 4671 downto 4640) <= CN145_sign_in;
    CN_data_in( 4703 downto 4672) <= CN146_data_in;
    CN_sign_in( 4703 downto 4672) <= CN146_sign_in;
    CN_data_in( 4735 downto 4704) <= CN147_data_in;
    CN_sign_in( 4735 downto 4704) <= CN147_sign_in;
    CN_data_in( 4767 downto 4736) <= CN148_data_in;
    CN_sign_in( 4767 downto 4736) <= CN148_sign_in;
    CN_data_in( 4799 downto 4768) <= CN149_data_in;
    CN_sign_in( 4799 downto 4768) <= CN149_sign_in;
    CN_data_in( 4831 downto 4800) <= CN150_data_in;
    CN_sign_in( 4831 downto 4800) <= CN150_sign_in;
    CN_data_in( 4863 downto 4832) <= CN151_data_in;
    CN_sign_in( 4863 downto 4832) <= CN151_sign_in;
    CN_data_in( 4895 downto 4864) <= CN152_data_in;
    CN_sign_in( 4895 downto 4864) <= CN152_sign_in;
    CN_data_in( 4927 downto 4896) <= CN153_data_in;
    CN_sign_in( 4927 downto 4896) <= CN153_sign_in;
    CN_data_in( 4959 downto 4928) <= CN154_data_in;
    CN_sign_in( 4959 downto 4928) <= CN154_sign_in;
    CN_data_in( 4991 downto 4960) <= CN155_data_in;
    CN_sign_in( 4991 downto 4960) <= CN155_sign_in;
    CN_data_in( 5023 downto 4992) <= CN156_data_in;
    CN_sign_in( 5023 downto 4992) <= CN156_sign_in;
    CN_data_in( 5055 downto 5024) <= CN157_data_in;
    CN_sign_in( 5055 downto 5024) <= CN157_sign_in;
    CN_data_in( 5087 downto 5056) <= CN158_data_in;
    CN_sign_in( 5087 downto 5056) <= CN158_sign_in;
    CN_data_in( 5119 downto 5088) <= CN159_data_in;
    CN_sign_in( 5119 downto 5088) <= CN159_sign_in;
    CN_data_in( 5151 downto 5120) <= CN160_data_in;
    CN_sign_in( 5151 downto 5120) <= CN160_sign_in;
    CN_data_in( 5183 downto 5152) <= CN161_data_in;
    CN_sign_in( 5183 downto 5152) <= CN161_sign_in;
    CN_data_in( 5215 downto 5184) <= CN162_data_in;
    CN_sign_in( 5215 downto 5184) <= CN162_sign_in;
    CN_data_in( 5247 downto 5216) <= CN163_data_in;
    CN_sign_in( 5247 downto 5216) <= CN163_sign_in;
    CN_data_in( 5279 downto 5248) <= CN164_data_in;
    CN_sign_in( 5279 downto 5248) <= CN164_sign_in;
    CN_data_in( 5311 downto 5280) <= CN165_data_in;
    CN_sign_in( 5311 downto 5280) <= CN165_sign_in;
    CN_data_in( 5343 downto 5312) <= CN166_data_in;
    CN_sign_in( 5343 downto 5312) <= CN166_sign_in;
    CN_data_in( 5375 downto 5344) <= CN167_data_in;
    CN_sign_in( 5375 downto 5344) <= CN167_sign_in;
    CN_data_in( 5407 downto 5376) <= CN168_data_in;
    CN_sign_in( 5407 downto 5376) <= CN168_sign_in;
    CN_data_in( 5439 downto 5408) <= CN169_data_in;
    CN_sign_in( 5439 downto 5408) <= CN169_sign_in;
    CN_data_in( 5471 downto 5440) <= CN170_data_in;
    CN_sign_in( 5471 downto 5440) <= CN170_sign_in;
    CN_data_in( 5503 downto 5472) <= CN171_data_in;
    CN_sign_in( 5503 downto 5472) <= CN171_sign_in;
    CN_data_in( 5535 downto 5504) <= CN172_data_in;
    CN_sign_in( 5535 downto 5504) <= CN172_sign_in;
    CN_data_in( 5567 downto 5536) <= CN173_data_in;
    CN_sign_in( 5567 downto 5536) <= CN173_sign_in;
    CN_data_in( 5599 downto 5568) <= CN174_data_in;
    CN_sign_in( 5599 downto 5568) <= CN174_sign_in;
    CN_data_in( 5631 downto 5600) <= CN175_data_in;
    CN_sign_in( 5631 downto 5600) <= CN175_sign_in;
    CN_data_in( 5663 downto 5632) <= CN176_data_in;
    CN_sign_in( 5663 downto 5632) <= CN176_sign_in;
    CN_data_in( 5695 downto 5664) <= CN177_data_in;
    CN_sign_in( 5695 downto 5664) <= CN177_sign_in;
    CN_data_in( 5727 downto 5696) <= CN178_data_in;
    CN_sign_in( 5727 downto 5696) <= CN178_sign_in;
    CN_data_in( 5759 downto 5728) <= CN179_data_in;
    CN_sign_in( 5759 downto 5728) <= CN179_sign_in;
    CN_data_in( 5791 downto 5760) <= CN180_data_in;
    CN_sign_in( 5791 downto 5760) <= CN180_sign_in;
    CN_data_in( 5823 downto 5792) <= CN181_data_in;
    CN_sign_in( 5823 downto 5792) <= CN181_sign_in;
    CN_data_in( 5855 downto 5824) <= CN182_data_in;
    CN_sign_in( 5855 downto 5824) <= CN182_sign_in;
    CN_data_in( 5887 downto 5856) <= CN183_data_in;
    CN_sign_in( 5887 downto 5856) <= CN183_sign_in;
    CN_data_in( 5919 downto 5888) <= CN184_data_in;
    CN_sign_in( 5919 downto 5888) <= CN184_sign_in;
    CN_data_in( 5951 downto 5920) <= CN185_data_in;
    CN_sign_in( 5951 downto 5920) <= CN185_sign_in;
    CN_data_in( 5983 downto 5952) <= CN186_data_in;
    CN_sign_in( 5983 downto 5952) <= CN186_sign_in;
    CN_data_in( 6015 downto 5984) <= CN187_data_in;
    CN_sign_in( 6015 downto 5984) <= CN187_sign_in;
    CN_data_in( 6047 downto 6016) <= CN188_data_in;
    CN_sign_in( 6047 downto 6016) <= CN188_sign_in;
    CN_data_in( 6079 downto 6048) <= CN189_data_in;
    CN_sign_in( 6079 downto 6048) <= CN189_sign_in;
    CN_data_in( 6111 downto 6080) <= CN190_data_in;
    CN_sign_in( 6111 downto 6080) <= CN190_sign_in;
    CN_data_in( 6143 downto 6112) <= CN191_data_in;
    CN_sign_in( 6143 downto 6112) <= CN191_sign_in;
    CN_data_in( 6175 downto 6144) <= CN192_data_in;
    CN_sign_in( 6175 downto 6144) <= CN192_sign_in;
    CN_data_in( 6207 downto 6176) <= CN193_data_in;
    CN_sign_in( 6207 downto 6176) <= CN193_sign_in;
    CN_data_in( 6239 downto 6208) <= CN194_data_in;
    CN_sign_in( 6239 downto 6208) <= CN194_sign_in;
    CN_data_in( 6271 downto 6240) <= CN195_data_in;
    CN_sign_in( 6271 downto 6240) <= CN195_sign_in;
    CN_data_in( 6303 downto 6272) <= CN196_data_in;
    CN_sign_in( 6303 downto 6272) <= CN196_sign_in;
    CN_data_in( 6335 downto 6304) <= CN197_data_in;
    CN_sign_in( 6335 downto 6304) <= CN197_sign_in;
    CN_data_in( 6367 downto 6336) <= CN198_data_in;
    CN_sign_in( 6367 downto 6336) <= CN198_sign_in;
    CN_data_in( 6399 downto 6368) <= CN199_data_in;
    CN_sign_in( 6399 downto 6368) <= CN199_sign_in;
    CN_data_in( 6431 downto 6400) <= CN200_data_in;
    CN_sign_in( 6431 downto 6400) <= CN200_sign_in;
    CN_data_in( 6463 downto 6432) <= CN201_data_in;
    CN_sign_in( 6463 downto 6432) <= CN201_sign_in;
    CN_data_in( 6495 downto 6464) <= CN202_data_in;
    CN_sign_in( 6495 downto 6464) <= CN202_sign_in;
    CN_data_in( 6527 downto 6496) <= CN203_data_in;
    CN_sign_in( 6527 downto 6496) <= CN203_sign_in;
    CN_data_in( 6559 downto 6528) <= CN204_data_in;
    CN_sign_in( 6559 downto 6528) <= CN204_sign_in;
    CN_data_in( 6591 downto 6560) <= CN205_data_in;
    CN_sign_in( 6591 downto 6560) <= CN205_sign_in;
    CN_data_in( 6623 downto 6592) <= CN206_data_in;
    CN_sign_in( 6623 downto 6592) <= CN206_sign_in;
    CN_data_in( 6655 downto 6624) <= CN207_data_in;
    CN_sign_in( 6655 downto 6624) <= CN207_sign_in;
    CN_data_in( 6687 downto 6656) <= CN208_data_in;
    CN_sign_in( 6687 downto 6656) <= CN208_sign_in;
    CN_data_in( 6719 downto 6688) <= CN209_data_in;
    CN_sign_in( 6719 downto 6688) <= CN209_sign_in;
    CN_data_in( 6751 downto 6720) <= CN210_data_in;
    CN_sign_in( 6751 downto 6720) <= CN210_sign_in;
    CN_data_in( 6783 downto 6752) <= CN211_data_in;
    CN_sign_in( 6783 downto 6752) <= CN211_sign_in;
    CN_data_in( 6815 downto 6784) <= CN212_data_in;
    CN_sign_in( 6815 downto 6784) <= CN212_sign_in;
    CN_data_in( 6847 downto 6816) <= CN213_data_in;
    CN_sign_in( 6847 downto 6816) <= CN213_sign_in;
    CN_data_in( 6879 downto 6848) <= CN214_data_in;
    CN_sign_in( 6879 downto 6848) <= CN214_sign_in;
    CN_data_in( 6911 downto 6880) <= CN215_data_in;
    CN_sign_in( 6911 downto 6880) <= CN215_sign_in;
    CN_data_in( 6943 downto 6912) <= CN216_data_in;
    CN_sign_in( 6943 downto 6912) <= CN216_sign_in;
    CN_data_in( 6975 downto 6944) <= CN217_data_in;
    CN_sign_in( 6975 downto 6944) <= CN217_sign_in;
    CN_data_in( 7007 downto 6976) <= CN218_data_in;
    CN_sign_in( 7007 downto 6976) <= CN218_sign_in;
    CN_data_in( 7039 downto 7008) <= CN219_data_in;
    CN_sign_in( 7039 downto 7008) <= CN219_sign_in;
    CN_data_in( 7071 downto 7040) <= CN220_data_in;
    CN_sign_in( 7071 downto 7040) <= CN220_sign_in;
    CN_data_in( 7103 downto 7072) <= CN221_data_in;
    CN_sign_in( 7103 downto 7072) <= CN221_sign_in;
    CN_data_in( 7135 downto 7104) <= CN222_data_in;
    CN_sign_in( 7135 downto 7104) <= CN222_sign_in;
    CN_data_in( 7167 downto 7136) <= CN223_data_in;
    CN_sign_in( 7167 downto 7136) <= CN223_sign_in;
    CN_data_in( 7199 downto 7168) <= CN224_data_in;
    CN_sign_in( 7199 downto 7168) <= CN224_sign_in;
    CN_data_in( 7231 downto 7200) <= CN225_data_in;
    CN_sign_in( 7231 downto 7200) <= CN225_sign_in;
    CN_data_in( 7263 downto 7232) <= CN226_data_in;
    CN_sign_in( 7263 downto 7232) <= CN226_sign_in;
    CN_data_in( 7295 downto 7264) <= CN227_data_in;
    CN_sign_in( 7295 downto 7264) <= CN227_sign_in;
    CN_data_in( 7327 downto 7296) <= CN228_data_in;
    CN_sign_in( 7327 downto 7296) <= CN228_sign_in;
    CN_data_in( 7359 downto 7328) <= CN229_data_in;
    CN_sign_in( 7359 downto 7328) <= CN229_sign_in;
    CN_data_in( 7391 downto 7360) <= CN230_data_in;
    CN_sign_in( 7391 downto 7360) <= CN230_sign_in;
    CN_data_in( 7423 downto 7392) <= CN231_data_in;
    CN_sign_in( 7423 downto 7392) <= CN231_sign_in;
    CN_data_in( 7455 downto 7424) <= CN232_data_in;
    CN_sign_in( 7455 downto 7424) <= CN232_sign_in;
    CN_data_in( 7487 downto 7456) <= CN233_data_in;
    CN_sign_in( 7487 downto 7456) <= CN233_sign_in;
    CN_data_in( 7519 downto 7488) <= CN234_data_in;
    CN_sign_in( 7519 downto 7488) <= CN234_sign_in;
    CN_data_in( 7551 downto 7520) <= CN235_data_in;
    CN_sign_in( 7551 downto 7520) <= CN235_sign_in;
    CN_data_in( 7583 downto 7552) <= CN236_data_in;
    CN_sign_in( 7583 downto 7552) <= CN236_sign_in;
    CN_data_in( 7615 downto 7584) <= CN237_data_in;
    CN_sign_in( 7615 downto 7584) <= CN237_sign_in;
    CN_data_in( 7647 downto 7616) <= CN238_data_in;
    CN_sign_in( 7647 downto 7616) <= CN238_sign_in;
    CN_data_in( 7679 downto 7648) <= CN239_data_in;
    CN_sign_in( 7679 downto 7648) <= CN239_sign_in;
    CN_data_in( 7711 downto 7680) <= CN240_data_in;
    CN_sign_in( 7711 downto 7680) <= CN240_sign_in;
    CN_data_in( 7743 downto 7712) <= CN241_data_in;
    CN_sign_in( 7743 downto 7712) <= CN241_sign_in;
    CN_data_in( 7775 downto 7744) <= CN242_data_in;
    CN_sign_in( 7775 downto 7744) <= CN242_sign_in;
    CN_data_in( 7807 downto 7776) <= CN243_data_in;
    CN_sign_in( 7807 downto 7776) <= CN243_sign_in;
    CN_data_in( 7839 downto 7808) <= CN244_data_in;
    CN_sign_in( 7839 downto 7808) <= CN244_sign_in;
    CN_data_in( 7871 downto 7840) <= CN245_data_in;
    CN_sign_in( 7871 downto 7840) <= CN245_sign_in;
    CN_data_in( 7903 downto 7872) <= CN246_data_in;
    CN_sign_in( 7903 downto 7872) <= CN246_sign_in;
    CN_data_in( 7935 downto 7904) <= CN247_data_in;
    CN_sign_in( 7935 downto 7904) <= CN247_sign_in;
    CN_data_in( 7967 downto 7936) <= CN248_data_in;
    CN_sign_in( 7967 downto 7936) <= CN248_sign_in;
    CN_data_in( 7999 downto 7968) <= CN249_data_in;
    CN_sign_in( 7999 downto 7968) <= CN249_sign_in;
    CN_data_in( 8031 downto 8000) <= CN250_data_in;
    CN_sign_in( 8031 downto 8000) <= CN250_sign_in;
    CN_data_in( 8063 downto 8032) <= CN251_data_in;
    CN_sign_in( 8063 downto 8032) <= CN251_sign_in;
    CN_data_in( 8095 downto 8064) <= CN252_data_in;
    CN_sign_in( 8095 downto 8064) <= CN252_sign_in;
    CN_data_in( 8127 downto 8096) <= CN253_data_in;
    CN_sign_in( 8127 downto 8096) <= CN253_sign_in;
    CN_data_in( 8159 downto 8128) <= CN254_data_in;
    CN_sign_in( 8159 downto 8128) <= CN254_sign_in;
    CN_data_in( 8191 downto 8160) <= CN255_data_in;
    CN_sign_in( 8191 downto 8160) <= CN255_sign_in;
    CN_data_in( 8223 downto 8192) <= CN256_data_in;
    CN_sign_in( 8223 downto 8192) <= CN256_sign_in;
    CN_data_in( 8255 downto 8224) <= CN257_data_in;
    CN_sign_in( 8255 downto 8224) <= CN257_sign_in;
    CN_data_in( 8287 downto 8256) <= CN258_data_in;
    CN_sign_in( 8287 downto 8256) <= CN258_sign_in;
    CN_data_in( 8319 downto 8288) <= CN259_data_in;
    CN_sign_in( 8319 downto 8288) <= CN259_sign_in;
    CN_data_in( 8351 downto 8320) <= CN260_data_in;
    CN_sign_in( 8351 downto 8320) <= CN260_sign_in;
    CN_data_in( 8383 downto 8352) <= CN261_data_in;
    CN_sign_in( 8383 downto 8352) <= CN261_sign_in;
    CN_data_in( 8415 downto 8384) <= CN262_data_in;
    CN_sign_in( 8415 downto 8384) <= CN262_sign_in;
    CN_data_in( 8447 downto 8416) <= CN263_data_in;
    CN_sign_in( 8447 downto 8416) <= CN263_sign_in;
    CN_data_in( 8479 downto 8448) <= CN264_data_in;
    CN_sign_in( 8479 downto 8448) <= CN264_sign_in;
    CN_data_in( 8511 downto 8480) <= CN265_data_in;
    CN_sign_in( 8511 downto 8480) <= CN265_sign_in;
    CN_data_in( 8543 downto 8512) <= CN266_data_in;
    CN_sign_in( 8543 downto 8512) <= CN266_sign_in;
    CN_data_in( 8575 downto 8544) <= CN267_data_in;
    CN_sign_in( 8575 downto 8544) <= CN267_sign_in;
    CN_data_in( 8607 downto 8576) <= CN268_data_in;
    CN_sign_in( 8607 downto 8576) <= CN268_sign_in;
    CN_data_in( 8639 downto 8608) <= CN269_data_in;
    CN_sign_in( 8639 downto 8608) <= CN269_sign_in;
    CN_data_in( 8671 downto 8640) <= CN270_data_in;
    CN_sign_in( 8671 downto 8640) <= CN270_sign_in;
    CN_data_in( 8703 downto 8672) <= CN271_data_in;
    CN_sign_in( 8703 downto 8672) <= CN271_sign_in;
    CN_data_in( 8735 downto 8704) <= CN272_data_in;
    CN_sign_in( 8735 downto 8704) <= CN272_sign_in;
    CN_data_in( 8767 downto 8736) <= CN273_data_in;
    CN_sign_in( 8767 downto 8736) <= CN273_sign_in;
    CN_data_in( 8799 downto 8768) <= CN274_data_in;
    CN_sign_in( 8799 downto 8768) <= CN274_sign_in;
    CN_data_in( 8831 downto 8800) <= CN275_data_in;
    CN_sign_in( 8831 downto 8800) <= CN275_sign_in;
    CN_data_in( 8863 downto 8832) <= CN276_data_in;
    CN_sign_in( 8863 downto 8832) <= CN276_sign_in;
    CN_data_in( 8895 downto 8864) <= CN277_data_in;
    CN_sign_in( 8895 downto 8864) <= CN277_sign_in;
    CN_data_in( 8927 downto 8896) <= CN278_data_in;
    CN_sign_in( 8927 downto 8896) <= CN278_sign_in;
    CN_data_in( 8959 downto 8928) <= CN279_data_in;
    CN_sign_in( 8959 downto 8928) <= CN279_sign_in;
    CN_data_in( 8991 downto 8960) <= CN280_data_in;
    CN_sign_in( 8991 downto 8960) <= CN280_sign_in;
    CN_data_in( 9023 downto 8992) <= CN281_data_in;
    CN_sign_in( 9023 downto 8992) <= CN281_sign_in;
    CN_data_in( 9055 downto 9024) <= CN282_data_in;
    CN_sign_in( 9055 downto 9024) <= CN282_sign_in;
    CN_data_in( 9087 downto 9056) <= CN283_data_in;
    CN_sign_in( 9087 downto 9056) <= CN283_sign_in;
    CN_data_in( 9119 downto 9088) <= CN284_data_in;
    CN_sign_in( 9119 downto 9088) <= CN284_sign_in;
    CN_data_in( 9151 downto 9120) <= CN285_data_in;
    CN_sign_in( 9151 downto 9120) <= CN285_sign_in;
    CN_data_in( 9183 downto 9152) <= CN286_data_in;
    CN_sign_in( 9183 downto 9152) <= CN286_sign_in;
    CN_data_in( 9215 downto 9184) <= CN287_data_in;
    CN_sign_in( 9215 downto 9184) <= CN287_sign_in;
    CN_data_in( 9247 downto 9216) <= CN288_data_in;
    CN_sign_in( 9247 downto 9216) <= CN288_sign_in;
    CN_data_in( 9279 downto 9248) <= CN289_data_in;
    CN_sign_in( 9279 downto 9248) <= CN289_sign_in;
    CN_data_in( 9311 downto 9280) <= CN290_data_in;
    CN_sign_in( 9311 downto 9280) <= CN290_sign_in;
    CN_data_in( 9343 downto 9312) <= CN291_data_in;
    CN_sign_in( 9343 downto 9312) <= CN291_sign_in;
    CN_data_in( 9375 downto 9344) <= CN292_data_in;
    CN_sign_in( 9375 downto 9344) <= CN292_sign_in;
    CN_data_in( 9407 downto 9376) <= CN293_data_in;
    CN_sign_in( 9407 downto 9376) <= CN293_sign_in;
    CN_data_in( 9439 downto 9408) <= CN294_data_in;
    CN_sign_in( 9439 downto 9408) <= CN294_sign_in;
    CN_data_in( 9471 downto 9440) <= CN295_data_in;
    CN_sign_in( 9471 downto 9440) <= CN295_sign_in;
    CN_data_in( 9503 downto 9472) <= CN296_data_in;
    CN_sign_in( 9503 downto 9472) <= CN296_sign_in;
    CN_data_in( 9535 downto 9504) <= CN297_data_in;
    CN_sign_in( 9535 downto 9504) <= CN297_sign_in;
    CN_data_in( 9567 downto 9536) <= CN298_data_in;
    CN_sign_in( 9567 downto 9536) <= CN298_sign_in;
    CN_data_in( 9599 downto 9568) <= CN299_data_in;
    CN_sign_in( 9599 downto 9568) <= CN299_sign_in;
    CN_data_in( 9631 downto 9600) <= CN300_data_in;
    CN_sign_in( 9631 downto 9600) <= CN300_sign_in;
    CN_data_in( 9663 downto 9632) <= CN301_data_in;
    CN_sign_in( 9663 downto 9632) <= CN301_sign_in;
    CN_data_in( 9695 downto 9664) <= CN302_data_in;
    CN_sign_in( 9695 downto 9664) <= CN302_sign_in;
    CN_data_in( 9727 downto 9696) <= CN303_data_in;
    CN_sign_in( 9727 downto 9696) <= CN303_sign_in;
    CN_data_in( 9759 downto 9728) <= CN304_data_in;
    CN_sign_in( 9759 downto 9728) <= CN304_sign_in;
    CN_data_in( 9791 downto 9760) <= CN305_data_in;
    CN_sign_in( 9791 downto 9760) <= CN305_sign_in;
    CN_data_in( 9823 downto 9792) <= CN306_data_in;
    CN_sign_in( 9823 downto 9792) <= CN306_sign_in;
    CN_data_in( 9855 downto 9824) <= CN307_data_in;
    CN_sign_in( 9855 downto 9824) <= CN307_sign_in;
    CN_data_in( 9887 downto 9856) <= CN308_data_in;
    CN_sign_in( 9887 downto 9856) <= CN308_sign_in;
    CN_data_in( 9919 downto 9888) <= CN309_data_in;
    CN_sign_in( 9919 downto 9888) <= CN309_sign_in;
    CN_data_in( 9951 downto 9920) <= CN310_data_in;
    CN_sign_in( 9951 downto 9920) <= CN310_sign_in;
    CN_data_in( 9983 downto 9952) <= CN311_data_in;
    CN_sign_in( 9983 downto 9952) <= CN311_sign_in;
    CN_data_in( 10015 downto 9984) <= CN312_data_in;
    CN_sign_in( 10015 downto 9984) <= CN312_sign_in;
    CN_data_in( 10047 downto 10016) <= CN313_data_in;
    CN_sign_in( 10047 downto 10016) <= CN313_sign_in;
    CN_data_in( 10079 downto 10048) <= CN314_data_in;
    CN_sign_in( 10079 downto 10048) <= CN314_sign_in;
    CN_data_in( 10111 downto 10080) <= CN315_data_in;
    CN_sign_in( 10111 downto 10080) <= CN315_sign_in;
    CN_data_in( 10143 downto 10112) <= CN316_data_in;
    CN_sign_in( 10143 downto 10112) <= CN316_sign_in;
    CN_data_in( 10175 downto 10144) <= CN317_data_in;
    CN_sign_in( 10175 downto 10144) <= CN317_sign_in;
    CN_data_in( 10207 downto 10176) <= CN318_data_in;
    CN_sign_in( 10207 downto 10176) <= CN318_sign_in;
    CN_data_in( 10239 downto 10208) <= CN319_data_in;
    CN_sign_in( 10239 downto 10208) <= CN319_sign_in;
    CN_data_in( 10271 downto 10240) <= CN320_data_in;
    CN_sign_in( 10271 downto 10240) <= CN320_sign_in;
    CN_data_in( 10303 downto 10272) <= CN321_data_in;
    CN_sign_in( 10303 downto 10272) <= CN321_sign_in;
    CN_data_in( 10335 downto 10304) <= CN322_data_in;
    CN_sign_in( 10335 downto 10304) <= CN322_sign_in;
    CN_data_in( 10367 downto 10336) <= CN323_data_in;
    CN_sign_in( 10367 downto 10336) <= CN323_sign_in;
    CN_data_in( 10399 downto 10368) <= CN324_data_in;
    CN_sign_in( 10399 downto 10368) <= CN324_sign_in;
    CN_data_in( 10431 downto 10400) <= CN325_data_in;
    CN_sign_in( 10431 downto 10400) <= CN325_sign_in;
    CN_data_in( 10463 downto 10432) <= CN326_data_in;
    CN_sign_in( 10463 downto 10432) <= CN326_sign_in;
    CN_data_in( 10495 downto 10464) <= CN327_data_in;
    CN_sign_in( 10495 downto 10464) <= CN327_sign_in;
    CN_data_in( 10527 downto 10496) <= CN328_data_in;
    CN_sign_in( 10527 downto 10496) <= CN328_sign_in;
    CN_data_in( 10559 downto 10528) <= CN329_data_in;
    CN_sign_in( 10559 downto 10528) <= CN329_sign_in;
    CN_data_in( 10591 downto 10560) <= CN330_data_in;
    CN_sign_in( 10591 downto 10560) <= CN330_sign_in;
    CN_data_in( 10623 downto 10592) <= CN331_data_in;
    CN_sign_in( 10623 downto 10592) <= CN331_sign_in;
    CN_data_in( 10655 downto 10624) <= CN332_data_in;
    CN_sign_in( 10655 downto 10624) <= CN332_sign_in;
    CN_data_in( 10687 downto 10656) <= CN333_data_in;
    CN_sign_in( 10687 downto 10656) <= CN333_sign_in;
    CN_data_in( 10719 downto 10688) <= CN334_data_in;
    CN_sign_in( 10719 downto 10688) <= CN334_sign_in;
    CN_data_in( 10751 downto 10720) <= CN335_data_in;
    CN_sign_in( 10751 downto 10720) <= CN335_sign_in;
    CN_data_in( 10783 downto 10752) <= CN336_data_in;
    CN_sign_in( 10783 downto 10752) <= CN336_sign_in;
    CN_data_in( 10815 downto 10784) <= CN337_data_in;
    CN_sign_in( 10815 downto 10784) <= CN337_sign_in;
    CN_data_in( 10847 downto 10816) <= CN338_data_in;
    CN_sign_in( 10847 downto 10816) <= CN338_sign_in;
    CN_data_in( 10879 downto 10848) <= CN339_data_in;
    CN_sign_in( 10879 downto 10848) <= CN339_sign_in;
    CN_data_in( 10911 downto 10880) <= CN340_data_in;
    CN_sign_in( 10911 downto 10880) <= CN340_sign_in;
    CN_data_in( 10943 downto 10912) <= CN341_data_in;
    CN_sign_in( 10943 downto 10912) <= CN341_sign_in;
    CN_data_in( 10975 downto 10944) <= CN342_data_in;
    CN_sign_in( 10975 downto 10944) <= CN342_sign_in;
    CN_data_in( 11007 downto 10976) <= CN343_data_in;
    CN_sign_in( 11007 downto 10976) <= CN343_sign_in;
    CN_data_in( 11039 downto 11008) <= CN344_data_in;
    CN_sign_in( 11039 downto 11008) <= CN344_sign_in;
    CN_data_in( 11071 downto 11040) <= CN345_data_in;
    CN_sign_in( 11071 downto 11040) <= CN345_sign_in;
    CN_data_in( 11103 downto 11072) <= CN346_data_in;
    CN_sign_in( 11103 downto 11072) <= CN346_sign_in;
    CN_data_in( 11135 downto 11104) <= CN347_data_in;
    CN_sign_in( 11135 downto 11104) <= CN347_sign_in;
    CN_data_in( 11167 downto 11136) <= CN348_data_in;
    CN_sign_in( 11167 downto 11136) <= CN348_sign_in;
    CN_data_in( 11199 downto 11168) <= CN349_data_in;
    CN_sign_in( 11199 downto 11168) <= CN349_sign_in;
    CN_data_in( 11231 downto 11200) <= CN350_data_in;
    CN_sign_in( 11231 downto 11200) <= CN350_sign_in;
    CN_data_in( 11263 downto 11232) <= CN351_data_in;
    CN_sign_in( 11263 downto 11232) <= CN351_sign_in;
    CN_data_in( 11295 downto 11264) <= CN352_data_in;
    CN_sign_in( 11295 downto 11264) <= CN352_sign_in;
    CN_data_in( 11327 downto 11296) <= CN353_data_in;
    CN_sign_in( 11327 downto 11296) <= CN353_sign_in;
    CN_data_in( 11359 downto 11328) <= CN354_data_in;
    CN_sign_in( 11359 downto 11328) <= CN354_sign_in;
    CN_data_in( 11391 downto 11360) <= CN355_data_in;
    CN_sign_in( 11391 downto 11360) <= CN355_sign_in;
    CN_data_in( 11423 downto 11392) <= CN356_data_in;
    CN_sign_in( 11423 downto 11392) <= CN356_sign_in;
    CN_data_in( 11455 downto 11424) <= CN357_data_in;
    CN_sign_in( 11455 downto 11424) <= CN357_sign_in;
    CN_data_in( 11487 downto 11456) <= CN358_data_in;
    CN_sign_in( 11487 downto 11456) <= CN358_sign_in;
    CN_data_in( 11519 downto 11488) <= CN359_data_in;
    CN_sign_in( 11519 downto 11488) <= CN359_sign_in;
    CN_data_in( 11551 downto 11520) <= CN360_data_in;
    CN_sign_in( 11551 downto 11520) <= CN360_sign_in;
    CN_data_in( 11583 downto 11552) <= CN361_data_in;
    CN_sign_in( 11583 downto 11552) <= CN361_sign_in;
    CN_data_in( 11615 downto 11584) <= CN362_data_in;
    CN_sign_in( 11615 downto 11584) <= CN362_sign_in;
    CN_data_in( 11647 downto 11616) <= CN363_data_in;
    CN_sign_in( 11647 downto 11616) <= CN363_sign_in;
    CN_data_in( 11679 downto 11648) <= CN364_data_in;
    CN_sign_in( 11679 downto 11648) <= CN364_sign_in;
    CN_data_in( 11711 downto 11680) <= CN365_data_in;
    CN_sign_in( 11711 downto 11680) <= CN365_sign_in;
    CN_data_in( 11743 downto 11712) <= CN366_data_in;
    CN_sign_in( 11743 downto 11712) <= CN366_sign_in;
    CN_data_in( 11775 downto 11744) <= CN367_data_in;
    CN_sign_in( 11775 downto 11744) <= CN367_sign_in;
    CN_data_in( 11807 downto 11776) <= CN368_data_in;
    CN_sign_in( 11807 downto 11776) <= CN368_sign_in;
    CN_data_in( 11839 downto 11808) <= CN369_data_in;
    CN_sign_in( 11839 downto 11808) <= CN369_sign_in;
    CN_data_in( 11871 downto 11840) <= CN370_data_in;
    CN_sign_in( 11871 downto 11840) <= CN370_sign_in;
    CN_data_in( 11903 downto 11872) <= CN371_data_in;
    CN_sign_in( 11903 downto 11872) <= CN371_sign_in;
    CN_data_in( 11935 downto 11904) <= CN372_data_in;
    CN_sign_in( 11935 downto 11904) <= CN372_sign_in;
    CN_data_in( 11967 downto 11936) <= CN373_data_in;
    CN_sign_in( 11967 downto 11936) <= CN373_sign_in;
    CN_data_in( 11999 downto 11968) <= CN374_data_in;
    CN_sign_in( 11999 downto 11968) <= CN374_sign_in;
    CN_data_in( 12031 downto 12000) <= CN375_data_in;
    CN_sign_in( 12031 downto 12000) <= CN375_sign_in;
    CN_data_in( 12063 downto 12032) <= CN376_data_in;
    CN_sign_in( 12063 downto 12032) <= CN376_sign_in;
    CN_data_in( 12095 downto 12064) <= CN377_data_in;
    CN_sign_in( 12095 downto 12064) <= CN377_sign_in;
    CN_data_in( 12127 downto 12096) <= CN378_data_in;
    CN_sign_in( 12127 downto 12096) <= CN378_sign_in;
    CN_data_in( 12159 downto 12128) <= CN379_data_in;
    CN_sign_in( 12159 downto 12128) <= CN379_sign_in;
    CN_data_in( 12191 downto 12160) <= CN380_data_in;
    CN_sign_in( 12191 downto 12160) <= CN380_sign_in;
    CN_data_in( 12223 downto 12192) <= CN381_data_in;
    CN_sign_in( 12223 downto 12192) <= CN381_sign_in;
    CN_data_in( 12255 downto 12224) <= CN382_data_in;
    CN_sign_in( 12255 downto 12224) <= CN382_sign_in;
    CN_data_in( 12287 downto 12256) <= CN383_data_in;
    CN_sign_in( 12287 downto 12256) <= CN383_sign_in;
    VN0_data_out <= VN_data_out( 5 downto 0 );
    VN0_sign_out <= VN_sign_out( 5 downto 0 );
    VN1_data_out <= VN_data_out( 11 downto 6 );
    VN1_sign_out <= VN_sign_out( 11 downto 6 );
    VN2_data_out <= VN_data_out( 17 downto 12 );
    VN2_sign_out <= VN_sign_out( 17 downto 12 );
    VN3_data_out <= VN_data_out( 23 downto 18 );
    VN3_sign_out <= VN_sign_out( 23 downto 18 );
    VN4_data_out <= VN_data_out( 29 downto 24 );
    VN4_sign_out <= VN_sign_out( 29 downto 24 );
    VN5_data_out <= VN_data_out( 35 downto 30 );
    VN5_sign_out <= VN_sign_out( 35 downto 30 );
    VN6_data_out <= VN_data_out( 41 downto 36 );
    VN6_sign_out <= VN_sign_out( 41 downto 36 );
    VN7_data_out <= VN_data_out( 47 downto 42 );
    VN7_sign_out <= VN_sign_out( 47 downto 42 );
    VN8_data_out <= VN_data_out( 53 downto 48 );
    VN8_sign_out <= VN_sign_out( 53 downto 48 );
    VN9_data_out <= VN_data_out( 59 downto 54 );
    VN9_sign_out <= VN_sign_out( 59 downto 54 );
    VN10_data_out <= VN_data_out( 65 downto 60 );
    VN10_sign_out <= VN_sign_out( 65 downto 60 );
    VN11_data_out <= VN_data_out( 71 downto 66 );
    VN11_sign_out <= VN_sign_out( 71 downto 66 );
    VN12_data_out <= VN_data_out( 77 downto 72 );
    VN12_sign_out <= VN_sign_out( 77 downto 72 );
    VN13_data_out <= VN_data_out( 83 downto 78 );
    VN13_sign_out <= VN_sign_out( 83 downto 78 );
    VN14_data_out <= VN_data_out( 89 downto 84 );
    VN14_sign_out <= VN_sign_out( 89 downto 84 );
    VN15_data_out <= VN_data_out( 95 downto 90 );
    VN15_sign_out <= VN_sign_out( 95 downto 90 );
    VN16_data_out <= VN_data_out( 101 downto 96 );
    VN16_sign_out <= VN_sign_out( 101 downto 96 );
    VN17_data_out <= VN_data_out( 107 downto 102 );
    VN17_sign_out <= VN_sign_out( 107 downto 102 );
    VN18_data_out <= VN_data_out( 113 downto 108 );
    VN18_sign_out <= VN_sign_out( 113 downto 108 );
    VN19_data_out <= VN_data_out( 119 downto 114 );
    VN19_sign_out <= VN_sign_out( 119 downto 114 );
    VN20_data_out <= VN_data_out( 125 downto 120 );
    VN20_sign_out <= VN_sign_out( 125 downto 120 );
    VN21_data_out <= VN_data_out( 131 downto 126 );
    VN21_sign_out <= VN_sign_out( 131 downto 126 );
    VN22_data_out <= VN_data_out( 137 downto 132 );
    VN22_sign_out <= VN_sign_out( 137 downto 132 );
    VN23_data_out <= VN_data_out( 143 downto 138 );
    VN23_sign_out <= VN_sign_out( 143 downto 138 );
    VN24_data_out <= VN_data_out( 149 downto 144 );
    VN24_sign_out <= VN_sign_out( 149 downto 144 );
    VN25_data_out <= VN_data_out( 155 downto 150 );
    VN25_sign_out <= VN_sign_out( 155 downto 150 );
    VN26_data_out <= VN_data_out( 161 downto 156 );
    VN26_sign_out <= VN_sign_out( 161 downto 156 );
    VN27_data_out <= VN_data_out( 167 downto 162 );
    VN27_sign_out <= VN_sign_out( 167 downto 162 );
    VN28_data_out <= VN_data_out( 173 downto 168 );
    VN28_sign_out <= VN_sign_out( 173 downto 168 );
    VN29_data_out <= VN_data_out( 179 downto 174 );
    VN29_sign_out <= VN_sign_out( 179 downto 174 );
    VN30_data_out <= VN_data_out( 185 downto 180 );
    VN30_sign_out <= VN_sign_out( 185 downto 180 );
    VN31_data_out <= VN_data_out( 191 downto 186 );
    VN31_sign_out <= VN_sign_out( 191 downto 186 );
    VN32_data_out <= VN_data_out( 197 downto 192 );
    VN32_sign_out <= VN_sign_out( 197 downto 192 );
    VN33_data_out <= VN_data_out( 203 downto 198 );
    VN33_sign_out <= VN_sign_out( 203 downto 198 );
    VN34_data_out <= VN_data_out( 209 downto 204 );
    VN34_sign_out <= VN_sign_out( 209 downto 204 );
    VN35_data_out <= VN_data_out( 215 downto 210 );
    VN35_sign_out <= VN_sign_out( 215 downto 210 );
    VN36_data_out <= VN_data_out( 221 downto 216 );
    VN36_sign_out <= VN_sign_out( 221 downto 216 );
    VN37_data_out <= VN_data_out( 227 downto 222 );
    VN37_sign_out <= VN_sign_out( 227 downto 222 );
    VN38_data_out <= VN_data_out( 233 downto 228 );
    VN38_sign_out <= VN_sign_out( 233 downto 228 );
    VN39_data_out <= VN_data_out( 239 downto 234 );
    VN39_sign_out <= VN_sign_out( 239 downto 234 );
    VN40_data_out <= VN_data_out( 245 downto 240 );
    VN40_sign_out <= VN_sign_out( 245 downto 240 );
    VN41_data_out <= VN_data_out( 251 downto 246 );
    VN41_sign_out <= VN_sign_out( 251 downto 246 );
    VN42_data_out <= VN_data_out( 257 downto 252 );
    VN42_sign_out <= VN_sign_out( 257 downto 252 );
    VN43_data_out <= VN_data_out( 263 downto 258 );
    VN43_sign_out <= VN_sign_out( 263 downto 258 );
    VN44_data_out <= VN_data_out( 269 downto 264 );
    VN44_sign_out <= VN_sign_out( 269 downto 264 );
    VN45_data_out <= VN_data_out( 275 downto 270 );
    VN45_sign_out <= VN_sign_out( 275 downto 270 );
    VN46_data_out <= VN_data_out( 281 downto 276 );
    VN46_sign_out <= VN_sign_out( 281 downto 276 );
    VN47_data_out <= VN_data_out( 287 downto 282 );
    VN47_sign_out <= VN_sign_out( 287 downto 282 );
    VN48_data_out <= VN_data_out( 293 downto 288 );
    VN48_sign_out <= VN_sign_out( 293 downto 288 );
    VN49_data_out <= VN_data_out( 299 downto 294 );
    VN49_sign_out <= VN_sign_out( 299 downto 294 );
    VN50_data_out <= VN_data_out( 305 downto 300 );
    VN50_sign_out <= VN_sign_out( 305 downto 300 );
    VN51_data_out <= VN_data_out( 311 downto 306 );
    VN51_sign_out <= VN_sign_out( 311 downto 306 );
    VN52_data_out <= VN_data_out( 317 downto 312 );
    VN52_sign_out <= VN_sign_out( 317 downto 312 );
    VN53_data_out <= VN_data_out( 323 downto 318 );
    VN53_sign_out <= VN_sign_out( 323 downto 318 );
    VN54_data_out <= VN_data_out( 329 downto 324 );
    VN54_sign_out <= VN_sign_out( 329 downto 324 );
    VN55_data_out <= VN_data_out( 335 downto 330 );
    VN55_sign_out <= VN_sign_out( 335 downto 330 );
    VN56_data_out <= VN_data_out( 341 downto 336 );
    VN56_sign_out <= VN_sign_out( 341 downto 336 );
    VN57_data_out <= VN_data_out( 347 downto 342 );
    VN57_sign_out <= VN_sign_out( 347 downto 342 );
    VN58_data_out <= VN_data_out( 353 downto 348 );
    VN58_sign_out <= VN_sign_out( 353 downto 348 );
    VN59_data_out <= VN_data_out( 359 downto 354 );
    VN59_sign_out <= VN_sign_out( 359 downto 354 );
    VN60_data_out <= VN_data_out( 365 downto 360 );
    VN60_sign_out <= VN_sign_out( 365 downto 360 );
    VN61_data_out <= VN_data_out( 371 downto 366 );
    VN61_sign_out <= VN_sign_out( 371 downto 366 );
    VN62_data_out <= VN_data_out( 377 downto 372 );
    VN62_sign_out <= VN_sign_out( 377 downto 372 );
    VN63_data_out <= VN_data_out( 383 downto 378 );
    VN63_sign_out <= VN_sign_out( 383 downto 378 );
    VN64_data_out <= VN_data_out( 389 downto 384 );
    VN64_sign_out <= VN_sign_out( 389 downto 384 );
    VN65_data_out <= VN_data_out( 395 downto 390 );
    VN65_sign_out <= VN_sign_out( 395 downto 390 );
    VN66_data_out <= VN_data_out( 401 downto 396 );
    VN66_sign_out <= VN_sign_out( 401 downto 396 );
    VN67_data_out <= VN_data_out( 407 downto 402 );
    VN67_sign_out <= VN_sign_out( 407 downto 402 );
    VN68_data_out <= VN_data_out( 413 downto 408 );
    VN68_sign_out <= VN_sign_out( 413 downto 408 );
    VN69_data_out <= VN_data_out( 419 downto 414 );
    VN69_sign_out <= VN_sign_out( 419 downto 414 );
    VN70_data_out <= VN_data_out( 425 downto 420 );
    VN70_sign_out <= VN_sign_out( 425 downto 420 );
    VN71_data_out <= VN_data_out( 431 downto 426 );
    VN71_sign_out <= VN_sign_out( 431 downto 426 );
    VN72_data_out <= VN_data_out( 437 downto 432 );
    VN72_sign_out <= VN_sign_out( 437 downto 432 );
    VN73_data_out <= VN_data_out( 443 downto 438 );
    VN73_sign_out <= VN_sign_out( 443 downto 438 );
    VN74_data_out <= VN_data_out( 449 downto 444 );
    VN74_sign_out <= VN_sign_out( 449 downto 444 );
    VN75_data_out <= VN_data_out( 455 downto 450 );
    VN75_sign_out <= VN_sign_out( 455 downto 450 );
    VN76_data_out <= VN_data_out( 461 downto 456 );
    VN76_sign_out <= VN_sign_out( 461 downto 456 );
    VN77_data_out <= VN_data_out( 467 downto 462 );
    VN77_sign_out <= VN_sign_out( 467 downto 462 );
    VN78_data_out <= VN_data_out( 473 downto 468 );
    VN78_sign_out <= VN_sign_out( 473 downto 468 );
    VN79_data_out <= VN_data_out( 479 downto 474 );
    VN79_sign_out <= VN_sign_out( 479 downto 474 );
    VN80_data_out <= VN_data_out( 485 downto 480 );
    VN80_sign_out <= VN_sign_out( 485 downto 480 );
    VN81_data_out <= VN_data_out( 491 downto 486 );
    VN81_sign_out <= VN_sign_out( 491 downto 486 );
    VN82_data_out <= VN_data_out( 497 downto 492 );
    VN82_sign_out <= VN_sign_out( 497 downto 492 );
    VN83_data_out <= VN_data_out( 503 downto 498 );
    VN83_sign_out <= VN_sign_out( 503 downto 498 );
    VN84_data_out <= VN_data_out( 509 downto 504 );
    VN84_sign_out <= VN_sign_out( 509 downto 504 );
    VN85_data_out <= VN_data_out( 515 downto 510 );
    VN85_sign_out <= VN_sign_out( 515 downto 510 );
    VN86_data_out <= VN_data_out( 521 downto 516 );
    VN86_sign_out <= VN_sign_out( 521 downto 516 );
    VN87_data_out <= VN_data_out( 527 downto 522 );
    VN87_sign_out <= VN_sign_out( 527 downto 522 );
    VN88_data_out <= VN_data_out( 533 downto 528 );
    VN88_sign_out <= VN_sign_out( 533 downto 528 );
    VN89_data_out <= VN_data_out( 539 downto 534 );
    VN89_sign_out <= VN_sign_out( 539 downto 534 );
    VN90_data_out <= VN_data_out( 545 downto 540 );
    VN90_sign_out <= VN_sign_out( 545 downto 540 );
    VN91_data_out <= VN_data_out( 551 downto 546 );
    VN91_sign_out <= VN_sign_out( 551 downto 546 );
    VN92_data_out <= VN_data_out( 557 downto 552 );
    VN92_sign_out <= VN_sign_out( 557 downto 552 );
    VN93_data_out <= VN_data_out( 563 downto 558 );
    VN93_sign_out <= VN_sign_out( 563 downto 558 );
    VN94_data_out <= VN_data_out( 569 downto 564 );
    VN94_sign_out <= VN_sign_out( 569 downto 564 );
    VN95_data_out <= VN_data_out( 575 downto 570 );
    VN95_sign_out <= VN_sign_out( 575 downto 570 );
    VN96_data_out <= VN_data_out( 581 downto 576 );
    VN96_sign_out <= VN_sign_out( 581 downto 576 );
    VN97_data_out <= VN_data_out( 587 downto 582 );
    VN97_sign_out <= VN_sign_out( 587 downto 582 );
    VN98_data_out <= VN_data_out( 593 downto 588 );
    VN98_sign_out <= VN_sign_out( 593 downto 588 );
    VN99_data_out <= VN_data_out( 599 downto 594 );
    VN99_sign_out <= VN_sign_out( 599 downto 594 );
    VN100_data_out <= VN_data_out( 605 downto 600 );
    VN100_sign_out <= VN_sign_out( 605 downto 600 );
    VN101_data_out <= VN_data_out( 611 downto 606 );
    VN101_sign_out <= VN_sign_out( 611 downto 606 );
    VN102_data_out <= VN_data_out( 617 downto 612 );
    VN102_sign_out <= VN_sign_out( 617 downto 612 );
    VN103_data_out <= VN_data_out( 623 downto 618 );
    VN103_sign_out <= VN_sign_out( 623 downto 618 );
    VN104_data_out <= VN_data_out( 629 downto 624 );
    VN104_sign_out <= VN_sign_out( 629 downto 624 );
    VN105_data_out <= VN_data_out( 635 downto 630 );
    VN105_sign_out <= VN_sign_out( 635 downto 630 );
    VN106_data_out <= VN_data_out( 641 downto 636 );
    VN106_sign_out <= VN_sign_out( 641 downto 636 );
    VN107_data_out <= VN_data_out( 647 downto 642 );
    VN107_sign_out <= VN_sign_out( 647 downto 642 );
    VN108_data_out <= VN_data_out( 653 downto 648 );
    VN108_sign_out <= VN_sign_out( 653 downto 648 );
    VN109_data_out <= VN_data_out( 659 downto 654 );
    VN109_sign_out <= VN_sign_out( 659 downto 654 );
    VN110_data_out <= VN_data_out( 665 downto 660 );
    VN110_sign_out <= VN_sign_out( 665 downto 660 );
    VN111_data_out <= VN_data_out( 671 downto 666 );
    VN111_sign_out <= VN_sign_out( 671 downto 666 );
    VN112_data_out <= VN_data_out( 677 downto 672 );
    VN112_sign_out <= VN_sign_out( 677 downto 672 );
    VN113_data_out <= VN_data_out( 683 downto 678 );
    VN113_sign_out <= VN_sign_out( 683 downto 678 );
    VN114_data_out <= VN_data_out( 689 downto 684 );
    VN114_sign_out <= VN_sign_out( 689 downto 684 );
    VN115_data_out <= VN_data_out( 695 downto 690 );
    VN115_sign_out <= VN_sign_out( 695 downto 690 );
    VN116_data_out <= VN_data_out( 701 downto 696 );
    VN116_sign_out <= VN_sign_out( 701 downto 696 );
    VN117_data_out <= VN_data_out( 707 downto 702 );
    VN117_sign_out <= VN_sign_out( 707 downto 702 );
    VN118_data_out <= VN_data_out( 713 downto 708 );
    VN118_sign_out <= VN_sign_out( 713 downto 708 );
    VN119_data_out <= VN_data_out( 719 downto 714 );
    VN119_sign_out <= VN_sign_out( 719 downto 714 );
    VN120_data_out <= VN_data_out( 725 downto 720 );
    VN120_sign_out <= VN_sign_out( 725 downto 720 );
    VN121_data_out <= VN_data_out( 731 downto 726 );
    VN121_sign_out <= VN_sign_out( 731 downto 726 );
    VN122_data_out <= VN_data_out( 737 downto 732 );
    VN122_sign_out <= VN_sign_out( 737 downto 732 );
    VN123_data_out <= VN_data_out( 743 downto 738 );
    VN123_sign_out <= VN_sign_out( 743 downto 738 );
    VN124_data_out <= VN_data_out( 749 downto 744 );
    VN124_sign_out <= VN_sign_out( 749 downto 744 );
    VN125_data_out <= VN_data_out( 755 downto 750 );
    VN125_sign_out <= VN_sign_out( 755 downto 750 );
    VN126_data_out <= VN_data_out( 761 downto 756 );
    VN126_sign_out <= VN_sign_out( 761 downto 756 );
    VN127_data_out <= VN_data_out( 767 downto 762 );
    VN127_sign_out <= VN_sign_out( 767 downto 762 );
    VN128_data_out <= VN_data_out( 773 downto 768 );
    VN128_sign_out <= VN_sign_out( 773 downto 768 );
    VN129_data_out <= VN_data_out( 779 downto 774 );
    VN129_sign_out <= VN_sign_out( 779 downto 774 );
    VN130_data_out <= VN_data_out( 785 downto 780 );
    VN130_sign_out <= VN_sign_out( 785 downto 780 );
    VN131_data_out <= VN_data_out( 791 downto 786 );
    VN131_sign_out <= VN_sign_out( 791 downto 786 );
    VN132_data_out <= VN_data_out( 797 downto 792 );
    VN132_sign_out <= VN_sign_out( 797 downto 792 );
    VN133_data_out <= VN_data_out( 803 downto 798 );
    VN133_sign_out <= VN_sign_out( 803 downto 798 );
    VN134_data_out <= VN_data_out( 809 downto 804 );
    VN134_sign_out <= VN_sign_out( 809 downto 804 );
    VN135_data_out <= VN_data_out( 815 downto 810 );
    VN135_sign_out <= VN_sign_out( 815 downto 810 );
    VN136_data_out <= VN_data_out( 821 downto 816 );
    VN136_sign_out <= VN_sign_out( 821 downto 816 );
    VN137_data_out <= VN_data_out( 827 downto 822 );
    VN137_sign_out <= VN_sign_out( 827 downto 822 );
    VN138_data_out <= VN_data_out( 833 downto 828 );
    VN138_sign_out <= VN_sign_out( 833 downto 828 );
    VN139_data_out <= VN_data_out( 839 downto 834 );
    VN139_sign_out <= VN_sign_out( 839 downto 834 );
    VN140_data_out <= VN_data_out( 845 downto 840 );
    VN140_sign_out <= VN_sign_out( 845 downto 840 );
    VN141_data_out <= VN_data_out( 851 downto 846 );
    VN141_sign_out <= VN_sign_out( 851 downto 846 );
    VN142_data_out <= VN_data_out( 857 downto 852 );
    VN142_sign_out <= VN_sign_out( 857 downto 852 );
    VN143_data_out <= VN_data_out( 863 downto 858 );
    VN143_sign_out <= VN_sign_out( 863 downto 858 );
    VN144_data_out <= VN_data_out( 869 downto 864 );
    VN144_sign_out <= VN_sign_out( 869 downto 864 );
    VN145_data_out <= VN_data_out( 875 downto 870 );
    VN145_sign_out <= VN_sign_out( 875 downto 870 );
    VN146_data_out <= VN_data_out( 881 downto 876 );
    VN146_sign_out <= VN_sign_out( 881 downto 876 );
    VN147_data_out <= VN_data_out( 887 downto 882 );
    VN147_sign_out <= VN_sign_out( 887 downto 882 );
    VN148_data_out <= VN_data_out( 893 downto 888 );
    VN148_sign_out <= VN_sign_out( 893 downto 888 );
    VN149_data_out <= VN_data_out( 899 downto 894 );
    VN149_sign_out <= VN_sign_out( 899 downto 894 );
    VN150_data_out <= VN_data_out( 905 downto 900 );
    VN150_sign_out <= VN_sign_out( 905 downto 900 );
    VN151_data_out <= VN_data_out( 911 downto 906 );
    VN151_sign_out <= VN_sign_out( 911 downto 906 );
    VN152_data_out <= VN_data_out( 917 downto 912 );
    VN152_sign_out <= VN_sign_out( 917 downto 912 );
    VN153_data_out <= VN_data_out( 923 downto 918 );
    VN153_sign_out <= VN_sign_out( 923 downto 918 );
    VN154_data_out <= VN_data_out( 929 downto 924 );
    VN154_sign_out <= VN_sign_out( 929 downto 924 );
    VN155_data_out <= VN_data_out( 935 downto 930 );
    VN155_sign_out <= VN_sign_out( 935 downto 930 );
    VN156_data_out <= VN_data_out( 941 downto 936 );
    VN156_sign_out <= VN_sign_out( 941 downto 936 );
    VN157_data_out <= VN_data_out( 947 downto 942 );
    VN157_sign_out <= VN_sign_out( 947 downto 942 );
    VN158_data_out <= VN_data_out( 953 downto 948 );
    VN158_sign_out <= VN_sign_out( 953 downto 948 );
    VN159_data_out <= VN_data_out( 959 downto 954 );
    VN159_sign_out <= VN_sign_out( 959 downto 954 );
    VN160_data_out <= VN_data_out( 965 downto 960 );
    VN160_sign_out <= VN_sign_out( 965 downto 960 );
    VN161_data_out <= VN_data_out( 971 downto 966 );
    VN161_sign_out <= VN_sign_out( 971 downto 966 );
    VN162_data_out <= VN_data_out( 977 downto 972 );
    VN162_sign_out <= VN_sign_out( 977 downto 972 );
    VN163_data_out <= VN_data_out( 983 downto 978 );
    VN163_sign_out <= VN_sign_out( 983 downto 978 );
    VN164_data_out <= VN_data_out( 989 downto 984 );
    VN164_sign_out <= VN_sign_out( 989 downto 984 );
    VN165_data_out <= VN_data_out( 995 downto 990 );
    VN165_sign_out <= VN_sign_out( 995 downto 990 );
    VN166_data_out <= VN_data_out( 1001 downto 996 );
    VN166_sign_out <= VN_sign_out( 1001 downto 996 );
    VN167_data_out <= VN_data_out( 1007 downto 1002 );
    VN167_sign_out <= VN_sign_out( 1007 downto 1002 );
    VN168_data_out <= VN_data_out( 1013 downto 1008 );
    VN168_sign_out <= VN_sign_out( 1013 downto 1008 );
    VN169_data_out <= VN_data_out( 1019 downto 1014 );
    VN169_sign_out <= VN_sign_out( 1019 downto 1014 );
    VN170_data_out <= VN_data_out( 1025 downto 1020 );
    VN170_sign_out <= VN_sign_out( 1025 downto 1020 );
    VN171_data_out <= VN_data_out( 1031 downto 1026 );
    VN171_sign_out <= VN_sign_out( 1031 downto 1026 );
    VN172_data_out <= VN_data_out( 1037 downto 1032 );
    VN172_sign_out <= VN_sign_out( 1037 downto 1032 );
    VN173_data_out <= VN_data_out( 1043 downto 1038 );
    VN173_sign_out <= VN_sign_out( 1043 downto 1038 );
    VN174_data_out <= VN_data_out( 1049 downto 1044 );
    VN174_sign_out <= VN_sign_out( 1049 downto 1044 );
    VN175_data_out <= VN_data_out( 1055 downto 1050 );
    VN175_sign_out <= VN_sign_out( 1055 downto 1050 );
    VN176_data_out <= VN_data_out( 1061 downto 1056 );
    VN176_sign_out <= VN_sign_out( 1061 downto 1056 );
    VN177_data_out <= VN_data_out( 1067 downto 1062 );
    VN177_sign_out <= VN_sign_out( 1067 downto 1062 );
    VN178_data_out <= VN_data_out( 1073 downto 1068 );
    VN178_sign_out <= VN_sign_out( 1073 downto 1068 );
    VN179_data_out <= VN_data_out( 1079 downto 1074 );
    VN179_sign_out <= VN_sign_out( 1079 downto 1074 );
    VN180_data_out <= VN_data_out( 1085 downto 1080 );
    VN180_sign_out <= VN_sign_out( 1085 downto 1080 );
    VN181_data_out <= VN_data_out( 1091 downto 1086 );
    VN181_sign_out <= VN_sign_out( 1091 downto 1086 );
    VN182_data_out <= VN_data_out( 1097 downto 1092 );
    VN182_sign_out <= VN_sign_out( 1097 downto 1092 );
    VN183_data_out <= VN_data_out( 1103 downto 1098 );
    VN183_sign_out <= VN_sign_out( 1103 downto 1098 );
    VN184_data_out <= VN_data_out( 1109 downto 1104 );
    VN184_sign_out <= VN_sign_out( 1109 downto 1104 );
    VN185_data_out <= VN_data_out( 1115 downto 1110 );
    VN185_sign_out <= VN_sign_out( 1115 downto 1110 );
    VN186_data_out <= VN_data_out( 1121 downto 1116 );
    VN186_sign_out <= VN_sign_out( 1121 downto 1116 );
    VN187_data_out <= VN_data_out( 1127 downto 1122 );
    VN187_sign_out <= VN_sign_out( 1127 downto 1122 );
    VN188_data_out <= VN_data_out( 1133 downto 1128 );
    VN188_sign_out <= VN_sign_out( 1133 downto 1128 );
    VN189_data_out <= VN_data_out( 1139 downto 1134 );
    VN189_sign_out <= VN_sign_out( 1139 downto 1134 );
    VN190_data_out <= VN_data_out( 1145 downto 1140 );
    VN190_sign_out <= VN_sign_out( 1145 downto 1140 );
    VN191_data_out <= VN_data_out( 1151 downto 1146 );
    VN191_sign_out <= VN_sign_out( 1151 downto 1146 );
    VN192_data_out <= VN_data_out( 1157 downto 1152 );
    VN192_sign_out <= VN_sign_out( 1157 downto 1152 );
    VN193_data_out <= VN_data_out( 1163 downto 1158 );
    VN193_sign_out <= VN_sign_out( 1163 downto 1158 );
    VN194_data_out <= VN_data_out( 1169 downto 1164 );
    VN194_sign_out <= VN_sign_out( 1169 downto 1164 );
    VN195_data_out <= VN_data_out( 1175 downto 1170 );
    VN195_sign_out <= VN_sign_out( 1175 downto 1170 );
    VN196_data_out <= VN_data_out( 1181 downto 1176 );
    VN196_sign_out <= VN_sign_out( 1181 downto 1176 );
    VN197_data_out <= VN_data_out( 1187 downto 1182 );
    VN197_sign_out <= VN_sign_out( 1187 downto 1182 );
    VN198_data_out <= VN_data_out( 1193 downto 1188 );
    VN198_sign_out <= VN_sign_out( 1193 downto 1188 );
    VN199_data_out <= VN_data_out( 1199 downto 1194 );
    VN199_sign_out <= VN_sign_out( 1199 downto 1194 );
    VN200_data_out <= VN_data_out( 1205 downto 1200 );
    VN200_sign_out <= VN_sign_out( 1205 downto 1200 );
    VN201_data_out <= VN_data_out( 1211 downto 1206 );
    VN201_sign_out <= VN_sign_out( 1211 downto 1206 );
    VN202_data_out <= VN_data_out( 1217 downto 1212 );
    VN202_sign_out <= VN_sign_out( 1217 downto 1212 );
    VN203_data_out <= VN_data_out( 1223 downto 1218 );
    VN203_sign_out <= VN_sign_out( 1223 downto 1218 );
    VN204_data_out <= VN_data_out( 1229 downto 1224 );
    VN204_sign_out <= VN_sign_out( 1229 downto 1224 );
    VN205_data_out <= VN_data_out( 1235 downto 1230 );
    VN205_sign_out <= VN_sign_out( 1235 downto 1230 );
    VN206_data_out <= VN_data_out( 1241 downto 1236 );
    VN206_sign_out <= VN_sign_out( 1241 downto 1236 );
    VN207_data_out <= VN_data_out( 1247 downto 1242 );
    VN207_sign_out <= VN_sign_out( 1247 downto 1242 );
    VN208_data_out <= VN_data_out( 1253 downto 1248 );
    VN208_sign_out <= VN_sign_out( 1253 downto 1248 );
    VN209_data_out <= VN_data_out( 1259 downto 1254 );
    VN209_sign_out <= VN_sign_out( 1259 downto 1254 );
    VN210_data_out <= VN_data_out( 1265 downto 1260 );
    VN210_sign_out <= VN_sign_out( 1265 downto 1260 );
    VN211_data_out <= VN_data_out( 1271 downto 1266 );
    VN211_sign_out <= VN_sign_out( 1271 downto 1266 );
    VN212_data_out <= VN_data_out( 1277 downto 1272 );
    VN212_sign_out <= VN_sign_out( 1277 downto 1272 );
    VN213_data_out <= VN_data_out( 1283 downto 1278 );
    VN213_sign_out <= VN_sign_out( 1283 downto 1278 );
    VN214_data_out <= VN_data_out( 1289 downto 1284 );
    VN214_sign_out <= VN_sign_out( 1289 downto 1284 );
    VN215_data_out <= VN_data_out( 1295 downto 1290 );
    VN215_sign_out <= VN_sign_out( 1295 downto 1290 );
    VN216_data_out <= VN_data_out( 1301 downto 1296 );
    VN216_sign_out <= VN_sign_out( 1301 downto 1296 );
    VN217_data_out <= VN_data_out( 1307 downto 1302 );
    VN217_sign_out <= VN_sign_out( 1307 downto 1302 );
    VN218_data_out <= VN_data_out( 1313 downto 1308 );
    VN218_sign_out <= VN_sign_out( 1313 downto 1308 );
    VN219_data_out <= VN_data_out( 1319 downto 1314 );
    VN219_sign_out <= VN_sign_out( 1319 downto 1314 );
    VN220_data_out <= VN_data_out( 1325 downto 1320 );
    VN220_sign_out <= VN_sign_out( 1325 downto 1320 );
    VN221_data_out <= VN_data_out( 1331 downto 1326 );
    VN221_sign_out <= VN_sign_out( 1331 downto 1326 );
    VN222_data_out <= VN_data_out( 1337 downto 1332 );
    VN222_sign_out <= VN_sign_out( 1337 downto 1332 );
    VN223_data_out <= VN_data_out( 1343 downto 1338 );
    VN223_sign_out <= VN_sign_out( 1343 downto 1338 );
    VN224_data_out <= VN_data_out( 1349 downto 1344 );
    VN224_sign_out <= VN_sign_out( 1349 downto 1344 );
    VN225_data_out <= VN_data_out( 1355 downto 1350 );
    VN225_sign_out <= VN_sign_out( 1355 downto 1350 );
    VN226_data_out <= VN_data_out( 1361 downto 1356 );
    VN226_sign_out <= VN_sign_out( 1361 downto 1356 );
    VN227_data_out <= VN_data_out( 1367 downto 1362 );
    VN227_sign_out <= VN_sign_out( 1367 downto 1362 );
    VN228_data_out <= VN_data_out( 1373 downto 1368 );
    VN228_sign_out <= VN_sign_out( 1373 downto 1368 );
    VN229_data_out <= VN_data_out( 1379 downto 1374 );
    VN229_sign_out <= VN_sign_out( 1379 downto 1374 );
    VN230_data_out <= VN_data_out( 1385 downto 1380 );
    VN230_sign_out <= VN_sign_out( 1385 downto 1380 );
    VN231_data_out <= VN_data_out( 1391 downto 1386 );
    VN231_sign_out <= VN_sign_out( 1391 downto 1386 );
    VN232_data_out <= VN_data_out( 1397 downto 1392 );
    VN232_sign_out <= VN_sign_out( 1397 downto 1392 );
    VN233_data_out <= VN_data_out( 1403 downto 1398 );
    VN233_sign_out <= VN_sign_out( 1403 downto 1398 );
    VN234_data_out <= VN_data_out( 1409 downto 1404 );
    VN234_sign_out <= VN_sign_out( 1409 downto 1404 );
    VN235_data_out <= VN_data_out( 1415 downto 1410 );
    VN235_sign_out <= VN_sign_out( 1415 downto 1410 );
    VN236_data_out <= VN_data_out( 1421 downto 1416 );
    VN236_sign_out <= VN_sign_out( 1421 downto 1416 );
    VN237_data_out <= VN_data_out( 1427 downto 1422 );
    VN237_sign_out <= VN_sign_out( 1427 downto 1422 );
    VN238_data_out <= VN_data_out( 1433 downto 1428 );
    VN238_sign_out <= VN_sign_out( 1433 downto 1428 );
    VN239_data_out <= VN_data_out( 1439 downto 1434 );
    VN239_sign_out <= VN_sign_out( 1439 downto 1434 );
    VN240_data_out <= VN_data_out( 1445 downto 1440 );
    VN240_sign_out <= VN_sign_out( 1445 downto 1440 );
    VN241_data_out <= VN_data_out( 1451 downto 1446 );
    VN241_sign_out <= VN_sign_out( 1451 downto 1446 );
    VN242_data_out <= VN_data_out( 1457 downto 1452 );
    VN242_sign_out <= VN_sign_out( 1457 downto 1452 );
    VN243_data_out <= VN_data_out( 1463 downto 1458 );
    VN243_sign_out <= VN_sign_out( 1463 downto 1458 );
    VN244_data_out <= VN_data_out( 1469 downto 1464 );
    VN244_sign_out <= VN_sign_out( 1469 downto 1464 );
    VN245_data_out <= VN_data_out( 1475 downto 1470 );
    VN245_sign_out <= VN_sign_out( 1475 downto 1470 );
    VN246_data_out <= VN_data_out( 1481 downto 1476 );
    VN246_sign_out <= VN_sign_out( 1481 downto 1476 );
    VN247_data_out <= VN_data_out( 1487 downto 1482 );
    VN247_sign_out <= VN_sign_out( 1487 downto 1482 );
    VN248_data_out <= VN_data_out( 1493 downto 1488 );
    VN248_sign_out <= VN_sign_out( 1493 downto 1488 );
    VN249_data_out <= VN_data_out( 1499 downto 1494 );
    VN249_sign_out <= VN_sign_out( 1499 downto 1494 );
    VN250_data_out <= VN_data_out( 1505 downto 1500 );
    VN250_sign_out <= VN_sign_out( 1505 downto 1500 );
    VN251_data_out <= VN_data_out( 1511 downto 1506 );
    VN251_sign_out <= VN_sign_out( 1511 downto 1506 );
    VN252_data_out <= VN_data_out( 1517 downto 1512 );
    VN252_sign_out <= VN_sign_out( 1517 downto 1512 );
    VN253_data_out <= VN_data_out( 1523 downto 1518 );
    VN253_sign_out <= VN_sign_out( 1523 downto 1518 );
    VN254_data_out <= VN_data_out( 1529 downto 1524 );
    VN254_sign_out <= VN_sign_out( 1529 downto 1524 );
    VN255_data_out <= VN_data_out( 1535 downto 1530 );
    VN255_sign_out <= VN_sign_out( 1535 downto 1530 );
    VN256_data_out <= VN_data_out( 1541 downto 1536 );
    VN256_sign_out <= VN_sign_out( 1541 downto 1536 );
    VN257_data_out <= VN_data_out( 1547 downto 1542 );
    VN257_sign_out <= VN_sign_out( 1547 downto 1542 );
    VN258_data_out <= VN_data_out( 1553 downto 1548 );
    VN258_sign_out <= VN_sign_out( 1553 downto 1548 );
    VN259_data_out <= VN_data_out( 1559 downto 1554 );
    VN259_sign_out <= VN_sign_out( 1559 downto 1554 );
    VN260_data_out <= VN_data_out( 1565 downto 1560 );
    VN260_sign_out <= VN_sign_out( 1565 downto 1560 );
    VN261_data_out <= VN_data_out( 1571 downto 1566 );
    VN261_sign_out <= VN_sign_out( 1571 downto 1566 );
    VN262_data_out <= VN_data_out( 1577 downto 1572 );
    VN262_sign_out <= VN_sign_out( 1577 downto 1572 );
    VN263_data_out <= VN_data_out( 1583 downto 1578 );
    VN263_sign_out <= VN_sign_out( 1583 downto 1578 );
    VN264_data_out <= VN_data_out( 1589 downto 1584 );
    VN264_sign_out <= VN_sign_out( 1589 downto 1584 );
    VN265_data_out <= VN_data_out( 1595 downto 1590 );
    VN265_sign_out <= VN_sign_out( 1595 downto 1590 );
    VN266_data_out <= VN_data_out( 1601 downto 1596 );
    VN266_sign_out <= VN_sign_out( 1601 downto 1596 );
    VN267_data_out <= VN_data_out( 1607 downto 1602 );
    VN267_sign_out <= VN_sign_out( 1607 downto 1602 );
    VN268_data_out <= VN_data_out( 1613 downto 1608 );
    VN268_sign_out <= VN_sign_out( 1613 downto 1608 );
    VN269_data_out <= VN_data_out( 1619 downto 1614 );
    VN269_sign_out <= VN_sign_out( 1619 downto 1614 );
    VN270_data_out <= VN_data_out( 1625 downto 1620 );
    VN270_sign_out <= VN_sign_out( 1625 downto 1620 );
    VN271_data_out <= VN_data_out( 1631 downto 1626 );
    VN271_sign_out <= VN_sign_out( 1631 downto 1626 );
    VN272_data_out <= VN_data_out( 1637 downto 1632 );
    VN272_sign_out <= VN_sign_out( 1637 downto 1632 );
    VN273_data_out <= VN_data_out( 1643 downto 1638 );
    VN273_sign_out <= VN_sign_out( 1643 downto 1638 );
    VN274_data_out <= VN_data_out( 1649 downto 1644 );
    VN274_sign_out <= VN_sign_out( 1649 downto 1644 );
    VN275_data_out <= VN_data_out( 1655 downto 1650 );
    VN275_sign_out <= VN_sign_out( 1655 downto 1650 );
    VN276_data_out <= VN_data_out( 1661 downto 1656 );
    VN276_sign_out <= VN_sign_out( 1661 downto 1656 );
    VN277_data_out <= VN_data_out( 1667 downto 1662 );
    VN277_sign_out <= VN_sign_out( 1667 downto 1662 );
    VN278_data_out <= VN_data_out( 1673 downto 1668 );
    VN278_sign_out <= VN_sign_out( 1673 downto 1668 );
    VN279_data_out <= VN_data_out( 1679 downto 1674 );
    VN279_sign_out <= VN_sign_out( 1679 downto 1674 );
    VN280_data_out <= VN_data_out( 1685 downto 1680 );
    VN280_sign_out <= VN_sign_out( 1685 downto 1680 );
    VN281_data_out <= VN_data_out( 1691 downto 1686 );
    VN281_sign_out <= VN_sign_out( 1691 downto 1686 );
    VN282_data_out <= VN_data_out( 1697 downto 1692 );
    VN282_sign_out <= VN_sign_out( 1697 downto 1692 );
    VN283_data_out <= VN_data_out( 1703 downto 1698 );
    VN283_sign_out <= VN_sign_out( 1703 downto 1698 );
    VN284_data_out <= VN_data_out( 1709 downto 1704 );
    VN284_sign_out <= VN_sign_out( 1709 downto 1704 );
    VN285_data_out <= VN_data_out( 1715 downto 1710 );
    VN285_sign_out <= VN_sign_out( 1715 downto 1710 );
    VN286_data_out <= VN_data_out( 1721 downto 1716 );
    VN286_sign_out <= VN_sign_out( 1721 downto 1716 );
    VN287_data_out <= VN_data_out( 1727 downto 1722 );
    VN287_sign_out <= VN_sign_out( 1727 downto 1722 );
    VN288_data_out <= VN_data_out( 1733 downto 1728 );
    VN288_sign_out <= VN_sign_out( 1733 downto 1728 );
    VN289_data_out <= VN_data_out( 1739 downto 1734 );
    VN289_sign_out <= VN_sign_out( 1739 downto 1734 );
    VN290_data_out <= VN_data_out( 1745 downto 1740 );
    VN290_sign_out <= VN_sign_out( 1745 downto 1740 );
    VN291_data_out <= VN_data_out( 1751 downto 1746 );
    VN291_sign_out <= VN_sign_out( 1751 downto 1746 );
    VN292_data_out <= VN_data_out( 1757 downto 1752 );
    VN292_sign_out <= VN_sign_out( 1757 downto 1752 );
    VN293_data_out <= VN_data_out( 1763 downto 1758 );
    VN293_sign_out <= VN_sign_out( 1763 downto 1758 );
    VN294_data_out <= VN_data_out( 1769 downto 1764 );
    VN294_sign_out <= VN_sign_out( 1769 downto 1764 );
    VN295_data_out <= VN_data_out( 1775 downto 1770 );
    VN295_sign_out <= VN_sign_out( 1775 downto 1770 );
    VN296_data_out <= VN_data_out( 1781 downto 1776 );
    VN296_sign_out <= VN_sign_out( 1781 downto 1776 );
    VN297_data_out <= VN_data_out( 1787 downto 1782 );
    VN297_sign_out <= VN_sign_out( 1787 downto 1782 );
    VN298_data_out <= VN_data_out( 1793 downto 1788 );
    VN298_sign_out <= VN_sign_out( 1793 downto 1788 );
    VN299_data_out <= VN_data_out( 1799 downto 1794 );
    VN299_sign_out <= VN_sign_out( 1799 downto 1794 );
    VN300_data_out <= VN_data_out( 1805 downto 1800 );
    VN300_sign_out <= VN_sign_out( 1805 downto 1800 );
    VN301_data_out <= VN_data_out( 1811 downto 1806 );
    VN301_sign_out <= VN_sign_out( 1811 downto 1806 );
    VN302_data_out <= VN_data_out( 1817 downto 1812 );
    VN302_sign_out <= VN_sign_out( 1817 downto 1812 );
    VN303_data_out <= VN_data_out( 1823 downto 1818 );
    VN303_sign_out <= VN_sign_out( 1823 downto 1818 );
    VN304_data_out <= VN_data_out( 1829 downto 1824 );
    VN304_sign_out <= VN_sign_out( 1829 downto 1824 );
    VN305_data_out <= VN_data_out( 1835 downto 1830 );
    VN305_sign_out <= VN_sign_out( 1835 downto 1830 );
    VN306_data_out <= VN_data_out( 1841 downto 1836 );
    VN306_sign_out <= VN_sign_out( 1841 downto 1836 );
    VN307_data_out <= VN_data_out( 1847 downto 1842 );
    VN307_sign_out <= VN_sign_out( 1847 downto 1842 );
    VN308_data_out <= VN_data_out( 1853 downto 1848 );
    VN308_sign_out <= VN_sign_out( 1853 downto 1848 );
    VN309_data_out <= VN_data_out( 1859 downto 1854 );
    VN309_sign_out <= VN_sign_out( 1859 downto 1854 );
    VN310_data_out <= VN_data_out( 1865 downto 1860 );
    VN310_sign_out <= VN_sign_out( 1865 downto 1860 );
    VN311_data_out <= VN_data_out( 1871 downto 1866 );
    VN311_sign_out <= VN_sign_out( 1871 downto 1866 );
    VN312_data_out <= VN_data_out( 1877 downto 1872 );
    VN312_sign_out <= VN_sign_out( 1877 downto 1872 );
    VN313_data_out <= VN_data_out( 1883 downto 1878 );
    VN313_sign_out <= VN_sign_out( 1883 downto 1878 );
    VN314_data_out <= VN_data_out( 1889 downto 1884 );
    VN314_sign_out <= VN_sign_out( 1889 downto 1884 );
    VN315_data_out <= VN_data_out( 1895 downto 1890 );
    VN315_sign_out <= VN_sign_out( 1895 downto 1890 );
    VN316_data_out <= VN_data_out( 1901 downto 1896 );
    VN316_sign_out <= VN_sign_out( 1901 downto 1896 );
    VN317_data_out <= VN_data_out( 1907 downto 1902 );
    VN317_sign_out <= VN_sign_out( 1907 downto 1902 );
    VN318_data_out <= VN_data_out( 1913 downto 1908 );
    VN318_sign_out <= VN_sign_out( 1913 downto 1908 );
    VN319_data_out <= VN_data_out( 1919 downto 1914 );
    VN319_sign_out <= VN_sign_out( 1919 downto 1914 );
    VN320_data_out <= VN_data_out( 1925 downto 1920 );
    VN320_sign_out <= VN_sign_out( 1925 downto 1920 );
    VN321_data_out <= VN_data_out( 1931 downto 1926 );
    VN321_sign_out <= VN_sign_out( 1931 downto 1926 );
    VN322_data_out <= VN_data_out( 1937 downto 1932 );
    VN322_sign_out <= VN_sign_out( 1937 downto 1932 );
    VN323_data_out <= VN_data_out( 1943 downto 1938 );
    VN323_sign_out <= VN_sign_out( 1943 downto 1938 );
    VN324_data_out <= VN_data_out( 1949 downto 1944 );
    VN324_sign_out <= VN_sign_out( 1949 downto 1944 );
    VN325_data_out <= VN_data_out( 1955 downto 1950 );
    VN325_sign_out <= VN_sign_out( 1955 downto 1950 );
    VN326_data_out <= VN_data_out( 1961 downto 1956 );
    VN326_sign_out <= VN_sign_out( 1961 downto 1956 );
    VN327_data_out <= VN_data_out( 1967 downto 1962 );
    VN327_sign_out <= VN_sign_out( 1967 downto 1962 );
    VN328_data_out <= VN_data_out( 1973 downto 1968 );
    VN328_sign_out <= VN_sign_out( 1973 downto 1968 );
    VN329_data_out <= VN_data_out( 1979 downto 1974 );
    VN329_sign_out <= VN_sign_out( 1979 downto 1974 );
    VN330_data_out <= VN_data_out( 1985 downto 1980 );
    VN330_sign_out <= VN_sign_out( 1985 downto 1980 );
    VN331_data_out <= VN_data_out( 1991 downto 1986 );
    VN331_sign_out <= VN_sign_out( 1991 downto 1986 );
    VN332_data_out <= VN_data_out( 1997 downto 1992 );
    VN332_sign_out <= VN_sign_out( 1997 downto 1992 );
    VN333_data_out <= VN_data_out( 2003 downto 1998 );
    VN333_sign_out <= VN_sign_out( 2003 downto 1998 );
    VN334_data_out <= VN_data_out( 2009 downto 2004 );
    VN334_sign_out <= VN_sign_out( 2009 downto 2004 );
    VN335_data_out <= VN_data_out( 2015 downto 2010 );
    VN335_sign_out <= VN_sign_out( 2015 downto 2010 );
    VN336_data_out <= VN_data_out( 2021 downto 2016 );
    VN336_sign_out <= VN_sign_out( 2021 downto 2016 );
    VN337_data_out <= VN_data_out( 2027 downto 2022 );
    VN337_sign_out <= VN_sign_out( 2027 downto 2022 );
    VN338_data_out <= VN_data_out( 2033 downto 2028 );
    VN338_sign_out <= VN_sign_out( 2033 downto 2028 );
    VN339_data_out <= VN_data_out( 2039 downto 2034 );
    VN339_sign_out <= VN_sign_out( 2039 downto 2034 );
    VN340_data_out <= VN_data_out( 2045 downto 2040 );
    VN340_sign_out <= VN_sign_out( 2045 downto 2040 );
    VN341_data_out <= VN_data_out( 2051 downto 2046 );
    VN341_sign_out <= VN_sign_out( 2051 downto 2046 );
    VN342_data_out <= VN_data_out( 2057 downto 2052 );
    VN342_sign_out <= VN_sign_out( 2057 downto 2052 );
    VN343_data_out <= VN_data_out( 2063 downto 2058 );
    VN343_sign_out <= VN_sign_out( 2063 downto 2058 );
    VN344_data_out <= VN_data_out( 2069 downto 2064 );
    VN344_sign_out <= VN_sign_out( 2069 downto 2064 );
    VN345_data_out <= VN_data_out( 2075 downto 2070 );
    VN345_sign_out <= VN_sign_out( 2075 downto 2070 );
    VN346_data_out <= VN_data_out( 2081 downto 2076 );
    VN346_sign_out <= VN_sign_out( 2081 downto 2076 );
    VN347_data_out <= VN_data_out( 2087 downto 2082 );
    VN347_sign_out <= VN_sign_out( 2087 downto 2082 );
    VN348_data_out <= VN_data_out( 2093 downto 2088 );
    VN348_sign_out <= VN_sign_out( 2093 downto 2088 );
    VN349_data_out <= VN_data_out( 2099 downto 2094 );
    VN349_sign_out <= VN_sign_out( 2099 downto 2094 );
    VN350_data_out <= VN_data_out( 2105 downto 2100 );
    VN350_sign_out <= VN_sign_out( 2105 downto 2100 );
    VN351_data_out <= VN_data_out( 2111 downto 2106 );
    VN351_sign_out <= VN_sign_out( 2111 downto 2106 );
    VN352_data_out <= VN_data_out( 2117 downto 2112 );
    VN352_sign_out <= VN_sign_out( 2117 downto 2112 );
    VN353_data_out <= VN_data_out( 2123 downto 2118 );
    VN353_sign_out <= VN_sign_out( 2123 downto 2118 );
    VN354_data_out <= VN_data_out( 2129 downto 2124 );
    VN354_sign_out <= VN_sign_out( 2129 downto 2124 );
    VN355_data_out <= VN_data_out( 2135 downto 2130 );
    VN355_sign_out <= VN_sign_out( 2135 downto 2130 );
    VN356_data_out <= VN_data_out( 2141 downto 2136 );
    VN356_sign_out <= VN_sign_out( 2141 downto 2136 );
    VN357_data_out <= VN_data_out( 2147 downto 2142 );
    VN357_sign_out <= VN_sign_out( 2147 downto 2142 );
    VN358_data_out <= VN_data_out( 2153 downto 2148 );
    VN358_sign_out <= VN_sign_out( 2153 downto 2148 );
    VN359_data_out <= VN_data_out( 2159 downto 2154 );
    VN359_sign_out <= VN_sign_out( 2159 downto 2154 );
    VN360_data_out <= VN_data_out( 2165 downto 2160 );
    VN360_sign_out <= VN_sign_out( 2165 downto 2160 );
    VN361_data_out <= VN_data_out( 2171 downto 2166 );
    VN361_sign_out <= VN_sign_out( 2171 downto 2166 );
    VN362_data_out <= VN_data_out( 2177 downto 2172 );
    VN362_sign_out <= VN_sign_out( 2177 downto 2172 );
    VN363_data_out <= VN_data_out( 2183 downto 2178 );
    VN363_sign_out <= VN_sign_out( 2183 downto 2178 );
    VN364_data_out <= VN_data_out( 2189 downto 2184 );
    VN364_sign_out <= VN_sign_out( 2189 downto 2184 );
    VN365_data_out <= VN_data_out( 2195 downto 2190 );
    VN365_sign_out <= VN_sign_out( 2195 downto 2190 );
    VN366_data_out <= VN_data_out( 2201 downto 2196 );
    VN366_sign_out <= VN_sign_out( 2201 downto 2196 );
    VN367_data_out <= VN_data_out( 2207 downto 2202 );
    VN367_sign_out <= VN_sign_out( 2207 downto 2202 );
    VN368_data_out <= VN_data_out( 2213 downto 2208 );
    VN368_sign_out <= VN_sign_out( 2213 downto 2208 );
    VN369_data_out <= VN_data_out( 2219 downto 2214 );
    VN369_sign_out <= VN_sign_out( 2219 downto 2214 );
    VN370_data_out <= VN_data_out( 2225 downto 2220 );
    VN370_sign_out <= VN_sign_out( 2225 downto 2220 );
    VN371_data_out <= VN_data_out( 2231 downto 2226 );
    VN371_sign_out <= VN_sign_out( 2231 downto 2226 );
    VN372_data_out <= VN_data_out( 2237 downto 2232 );
    VN372_sign_out <= VN_sign_out( 2237 downto 2232 );
    VN373_data_out <= VN_data_out( 2243 downto 2238 );
    VN373_sign_out <= VN_sign_out( 2243 downto 2238 );
    VN374_data_out <= VN_data_out( 2249 downto 2244 );
    VN374_sign_out <= VN_sign_out( 2249 downto 2244 );
    VN375_data_out <= VN_data_out( 2255 downto 2250 );
    VN375_sign_out <= VN_sign_out( 2255 downto 2250 );
    VN376_data_out <= VN_data_out( 2261 downto 2256 );
    VN376_sign_out <= VN_sign_out( 2261 downto 2256 );
    VN377_data_out <= VN_data_out( 2267 downto 2262 );
    VN377_sign_out <= VN_sign_out( 2267 downto 2262 );
    VN378_data_out <= VN_data_out( 2273 downto 2268 );
    VN378_sign_out <= VN_sign_out( 2273 downto 2268 );
    VN379_data_out <= VN_data_out( 2279 downto 2274 );
    VN379_sign_out <= VN_sign_out( 2279 downto 2274 );
    VN380_data_out <= VN_data_out( 2285 downto 2280 );
    VN380_sign_out <= VN_sign_out( 2285 downto 2280 );
    VN381_data_out <= VN_data_out( 2291 downto 2286 );
    VN381_sign_out <= VN_sign_out( 2291 downto 2286 );
    VN382_data_out <= VN_data_out( 2297 downto 2292 );
    VN382_sign_out <= VN_sign_out( 2297 downto 2292 );
    VN383_data_out <= VN_data_out( 2303 downto 2298 );
    VN383_sign_out <= VN_sign_out( 2303 downto 2298 );
    VN384_data_out <= VN_data_out( 2309 downto 2304 );
    VN384_sign_out <= VN_sign_out( 2309 downto 2304 );
    VN385_data_out <= VN_data_out( 2315 downto 2310 );
    VN385_sign_out <= VN_sign_out( 2315 downto 2310 );
    VN386_data_out <= VN_data_out( 2321 downto 2316 );
    VN386_sign_out <= VN_sign_out( 2321 downto 2316 );
    VN387_data_out <= VN_data_out( 2327 downto 2322 );
    VN387_sign_out <= VN_sign_out( 2327 downto 2322 );
    VN388_data_out <= VN_data_out( 2333 downto 2328 );
    VN388_sign_out <= VN_sign_out( 2333 downto 2328 );
    VN389_data_out <= VN_data_out( 2339 downto 2334 );
    VN389_sign_out <= VN_sign_out( 2339 downto 2334 );
    VN390_data_out <= VN_data_out( 2345 downto 2340 );
    VN390_sign_out <= VN_sign_out( 2345 downto 2340 );
    VN391_data_out <= VN_data_out( 2351 downto 2346 );
    VN391_sign_out <= VN_sign_out( 2351 downto 2346 );
    VN392_data_out <= VN_data_out( 2357 downto 2352 );
    VN392_sign_out <= VN_sign_out( 2357 downto 2352 );
    VN393_data_out <= VN_data_out( 2363 downto 2358 );
    VN393_sign_out <= VN_sign_out( 2363 downto 2358 );
    VN394_data_out <= VN_data_out( 2369 downto 2364 );
    VN394_sign_out <= VN_sign_out( 2369 downto 2364 );
    VN395_data_out <= VN_data_out( 2375 downto 2370 );
    VN395_sign_out <= VN_sign_out( 2375 downto 2370 );
    VN396_data_out <= VN_data_out( 2381 downto 2376 );
    VN396_sign_out <= VN_sign_out( 2381 downto 2376 );
    VN397_data_out <= VN_data_out( 2387 downto 2382 );
    VN397_sign_out <= VN_sign_out( 2387 downto 2382 );
    VN398_data_out <= VN_data_out( 2393 downto 2388 );
    VN398_sign_out <= VN_sign_out( 2393 downto 2388 );
    VN399_data_out <= VN_data_out( 2399 downto 2394 );
    VN399_sign_out <= VN_sign_out( 2399 downto 2394 );
    VN400_data_out <= VN_data_out( 2405 downto 2400 );
    VN400_sign_out <= VN_sign_out( 2405 downto 2400 );
    VN401_data_out <= VN_data_out( 2411 downto 2406 );
    VN401_sign_out <= VN_sign_out( 2411 downto 2406 );
    VN402_data_out <= VN_data_out( 2417 downto 2412 );
    VN402_sign_out <= VN_sign_out( 2417 downto 2412 );
    VN403_data_out <= VN_data_out( 2423 downto 2418 );
    VN403_sign_out <= VN_sign_out( 2423 downto 2418 );
    VN404_data_out <= VN_data_out( 2429 downto 2424 );
    VN404_sign_out <= VN_sign_out( 2429 downto 2424 );
    VN405_data_out <= VN_data_out( 2435 downto 2430 );
    VN405_sign_out <= VN_sign_out( 2435 downto 2430 );
    VN406_data_out <= VN_data_out( 2441 downto 2436 );
    VN406_sign_out <= VN_sign_out( 2441 downto 2436 );
    VN407_data_out <= VN_data_out( 2447 downto 2442 );
    VN407_sign_out <= VN_sign_out( 2447 downto 2442 );
    VN408_data_out <= VN_data_out( 2453 downto 2448 );
    VN408_sign_out <= VN_sign_out( 2453 downto 2448 );
    VN409_data_out <= VN_data_out( 2459 downto 2454 );
    VN409_sign_out <= VN_sign_out( 2459 downto 2454 );
    VN410_data_out <= VN_data_out( 2465 downto 2460 );
    VN410_sign_out <= VN_sign_out( 2465 downto 2460 );
    VN411_data_out <= VN_data_out( 2471 downto 2466 );
    VN411_sign_out <= VN_sign_out( 2471 downto 2466 );
    VN412_data_out <= VN_data_out( 2477 downto 2472 );
    VN412_sign_out <= VN_sign_out( 2477 downto 2472 );
    VN413_data_out <= VN_data_out( 2483 downto 2478 );
    VN413_sign_out <= VN_sign_out( 2483 downto 2478 );
    VN414_data_out <= VN_data_out( 2489 downto 2484 );
    VN414_sign_out <= VN_sign_out( 2489 downto 2484 );
    VN415_data_out <= VN_data_out( 2495 downto 2490 );
    VN415_sign_out <= VN_sign_out( 2495 downto 2490 );
    VN416_data_out <= VN_data_out( 2501 downto 2496 );
    VN416_sign_out <= VN_sign_out( 2501 downto 2496 );
    VN417_data_out <= VN_data_out( 2507 downto 2502 );
    VN417_sign_out <= VN_sign_out( 2507 downto 2502 );
    VN418_data_out <= VN_data_out( 2513 downto 2508 );
    VN418_sign_out <= VN_sign_out( 2513 downto 2508 );
    VN419_data_out <= VN_data_out( 2519 downto 2514 );
    VN419_sign_out <= VN_sign_out( 2519 downto 2514 );
    VN420_data_out <= VN_data_out( 2525 downto 2520 );
    VN420_sign_out <= VN_sign_out( 2525 downto 2520 );
    VN421_data_out <= VN_data_out( 2531 downto 2526 );
    VN421_sign_out <= VN_sign_out( 2531 downto 2526 );
    VN422_data_out <= VN_data_out( 2537 downto 2532 );
    VN422_sign_out <= VN_sign_out( 2537 downto 2532 );
    VN423_data_out <= VN_data_out( 2543 downto 2538 );
    VN423_sign_out <= VN_sign_out( 2543 downto 2538 );
    VN424_data_out <= VN_data_out( 2549 downto 2544 );
    VN424_sign_out <= VN_sign_out( 2549 downto 2544 );
    VN425_data_out <= VN_data_out( 2555 downto 2550 );
    VN425_sign_out <= VN_sign_out( 2555 downto 2550 );
    VN426_data_out <= VN_data_out( 2561 downto 2556 );
    VN426_sign_out <= VN_sign_out( 2561 downto 2556 );
    VN427_data_out <= VN_data_out( 2567 downto 2562 );
    VN427_sign_out <= VN_sign_out( 2567 downto 2562 );
    VN428_data_out <= VN_data_out( 2573 downto 2568 );
    VN428_sign_out <= VN_sign_out( 2573 downto 2568 );
    VN429_data_out <= VN_data_out( 2579 downto 2574 );
    VN429_sign_out <= VN_sign_out( 2579 downto 2574 );
    VN430_data_out <= VN_data_out( 2585 downto 2580 );
    VN430_sign_out <= VN_sign_out( 2585 downto 2580 );
    VN431_data_out <= VN_data_out( 2591 downto 2586 );
    VN431_sign_out <= VN_sign_out( 2591 downto 2586 );
    VN432_data_out <= VN_data_out( 2597 downto 2592 );
    VN432_sign_out <= VN_sign_out( 2597 downto 2592 );
    VN433_data_out <= VN_data_out( 2603 downto 2598 );
    VN433_sign_out <= VN_sign_out( 2603 downto 2598 );
    VN434_data_out <= VN_data_out( 2609 downto 2604 );
    VN434_sign_out <= VN_sign_out( 2609 downto 2604 );
    VN435_data_out <= VN_data_out( 2615 downto 2610 );
    VN435_sign_out <= VN_sign_out( 2615 downto 2610 );
    VN436_data_out <= VN_data_out( 2621 downto 2616 );
    VN436_sign_out <= VN_sign_out( 2621 downto 2616 );
    VN437_data_out <= VN_data_out( 2627 downto 2622 );
    VN437_sign_out <= VN_sign_out( 2627 downto 2622 );
    VN438_data_out <= VN_data_out( 2633 downto 2628 );
    VN438_sign_out <= VN_sign_out( 2633 downto 2628 );
    VN439_data_out <= VN_data_out( 2639 downto 2634 );
    VN439_sign_out <= VN_sign_out( 2639 downto 2634 );
    VN440_data_out <= VN_data_out( 2645 downto 2640 );
    VN440_sign_out <= VN_sign_out( 2645 downto 2640 );
    VN441_data_out <= VN_data_out( 2651 downto 2646 );
    VN441_sign_out <= VN_sign_out( 2651 downto 2646 );
    VN442_data_out <= VN_data_out( 2657 downto 2652 );
    VN442_sign_out <= VN_sign_out( 2657 downto 2652 );
    VN443_data_out <= VN_data_out( 2663 downto 2658 );
    VN443_sign_out <= VN_sign_out( 2663 downto 2658 );
    VN444_data_out <= VN_data_out( 2669 downto 2664 );
    VN444_sign_out <= VN_sign_out( 2669 downto 2664 );
    VN445_data_out <= VN_data_out( 2675 downto 2670 );
    VN445_sign_out <= VN_sign_out( 2675 downto 2670 );
    VN446_data_out <= VN_data_out( 2681 downto 2676 );
    VN446_sign_out <= VN_sign_out( 2681 downto 2676 );
    VN447_data_out <= VN_data_out( 2687 downto 2682 );
    VN447_sign_out <= VN_sign_out( 2687 downto 2682 );
    VN448_data_out <= VN_data_out( 2693 downto 2688 );
    VN448_sign_out <= VN_sign_out( 2693 downto 2688 );
    VN449_data_out <= VN_data_out( 2699 downto 2694 );
    VN449_sign_out <= VN_sign_out( 2699 downto 2694 );
    VN450_data_out <= VN_data_out( 2705 downto 2700 );
    VN450_sign_out <= VN_sign_out( 2705 downto 2700 );
    VN451_data_out <= VN_data_out( 2711 downto 2706 );
    VN451_sign_out <= VN_sign_out( 2711 downto 2706 );
    VN452_data_out <= VN_data_out( 2717 downto 2712 );
    VN452_sign_out <= VN_sign_out( 2717 downto 2712 );
    VN453_data_out <= VN_data_out( 2723 downto 2718 );
    VN453_sign_out <= VN_sign_out( 2723 downto 2718 );
    VN454_data_out <= VN_data_out( 2729 downto 2724 );
    VN454_sign_out <= VN_sign_out( 2729 downto 2724 );
    VN455_data_out <= VN_data_out( 2735 downto 2730 );
    VN455_sign_out <= VN_sign_out( 2735 downto 2730 );
    VN456_data_out <= VN_data_out( 2741 downto 2736 );
    VN456_sign_out <= VN_sign_out( 2741 downto 2736 );
    VN457_data_out <= VN_data_out( 2747 downto 2742 );
    VN457_sign_out <= VN_sign_out( 2747 downto 2742 );
    VN458_data_out <= VN_data_out( 2753 downto 2748 );
    VN458_sign_out <= VN_sign_out( 2753 downto 2748 );
    VN459_data_out <= VN_data_out( 2759 downto 2754 );
    VN459_sign_out <= VN_sign_out( 2759 downto 2754 );
    VN460_data_out <= VN_data_out( 2765 downto 2760 );
    VN460_sign_out <= VN_sign_out( 2765 downto 2760 );
    VN461_data_out <= VN_data_out( 2771 downto 2766 );
    VN461_sign_out <= VN_sign_out( 2771 downto 2766 );
    VN462_data_out <= VN_data_out( 2777 downto 2772 );
    VN462_sign_out <= VN_sign_out( 2777 downto 2772 );
    VN463_data_out <= VN_data_out( 2783 downto 2778 );
    VN463_sign_out <= VN_sign_out( 2783 downto 2778 );
    VN464_data_out <= VN_data_out( 2789 downto 2784 );
    VN464_sign_out <= VN_sign_out( 2789 downto 2784 );
    VN465_data_out <= VN_data_out( 2795 downto 2790 );
    VN465_sign_out <= VN_sign_out( 2795 downto 2790 );
    VN466_data_out <= VN_data_out( 2801 downto 2796 );
    VN466_sign_out <= VN_sign_out( 2801 downto 2796 );
    VN467_data_out <= VN_data_out( 2807 downto 2802 );
    VN467_sign_out <= VN_sign_out( 2807 downto 2802 );
    VN468_data_out <= VN_data_out( 2813 downto 2808 );
    VN468_sign_out <= VN_sign_out( 2813 downto 2808 );
    VN469_data_out <= VN_data_out( 2819 downto 2814 );
    VN469_sign_out <= VN_sign_out( 2819 downto 2814 );
    VN470_data_out <= VN_data_out( 2825 downto 2820 );
    VN470_sign_out <= VN_sign_out( 2825 downto 2820 );
    VN471_data_out <= VN_data_out( 2831 downto 2826 );
    VN471_sign_out <= VN_sign_out( 2831 downto 2826 );
    VN472_data_out <= VN_data_out( 2837 downto 2832 );
    VN472_sign_out <= VN_sign_out( 2837 downto 2832 );
    VN473_data_out <= VN_data_out( 2843 downto 2838 );
    VN473_sign_out <= VN_sign_out( 2843 downto 2838 );
    VN474_data_out <= VN_data_out( 2849 downto 2844 );
    VN474_sign_out <= VN_sign_out( 2849 downto 2844 );
    VN475_data_out <= VN_data_out( 2855 downto 2850 );
    VN475_sign_out <= VN_sign_out( 2855 downto 2850 );
    VN476_data_out <= VN_data_out( 2861 downto 2856 );
    VN476_sign_out <= VN_sign_out( 2861 downto 2856 );
    VN477_data_out <= VN_data_out( 2867 downto 2862 );
    VN477_sign_out <= VN_sign_out( 2867 downto 2862 );
    VN478_data_out <= VN_data_out( 2873 downto 2868 );
    VN478_sign_out <= VN_sign_out( 2873 downto 2868 );
    VN479_data_out <= VN_data_out( 2879 downto 2874 );
    VN479_sign_out <= VN_sign_out( 2879 downto 2874 );
    VN480_data_out <= VN_data_out( 2885 downto 2880 );
    VN480_sign_out <= VN_sign_out( 2885 downto 2880 );
    VN481_data_out <= VN_data_out( 2891 downto 2886 );
    VN481_sign_out <= VN_sign_out( 2891 downto 2886 );
    VN482_data_out <= VN_data_out( 2897 downto 2892 );
    VN482_sign_out <= VN_sign_out( 2897 downto 2892 );
    VN483_data_out <= VN_data_out( 2903 downto 2898 );
    VN483_sign_out <= VN_sign_out( 2903 downto 2898 );
    VN484_data_out <= VN_data_out( 2909 downto 2904 );
    VN484_sign_out <= VN_sign_out( 2909 downto 2904 );
    VN485_data_out <= VN_data_out( 2915 downto 2910 );
    VN485_sign_out <= VN_sign_out( 2915 downto 2910 );
    VN486_data_out <= VN_data_out( 2921 downto 2916 );
    VN486_sign_out <= VN_sign_out( 2921 downto 2916 );
    VN487_data_out <= VN_data_out( 2927 downto 2922 );
    VN487_sign_out <= VN_sign_out( 2927 downto 2922 );
    VN488_data_out <= VN_data_out( 2933 downto 2928 );
    VN488_sign_out <= VN_sign_out( 2933 downto 2928 );
    VN489_data_out <= VN_data_out( 2939 downto 2934 );
    VN489_sign_out <= VN_sign_out( 2939 downto 2934 );
    VN490_data_out <= VN_data_out( 2945 downto 2940 );
    VN490_sign_out <= VN_sign_out( 2945 downto 2940 );
    VN491_data_out <= VN_data_out( 2951 downto 2946 );
    VN491_sign_out <= VN_sign_out( 2951 downto 2946 );
    VN492_data_out <= VN_data_out( 2957 downto 2952 );
    VN492_sign_out <= VN_sign_out( 2957 downto 2952 );
    VN493_data_out <= VN_data_out( 2963 downto 2958 );
    VN493_sign_out <= VN_sign_out( 2963 downto 2958 );
    VN494_data_out <= VN_data_out( 2969 downto 2964 );
    VN494_sign_out <= VN_sign_out( 2969 downto 2964 );
    VN495_data_out <= VN_data_out( 2975 downto 2970 );
    VN495_sign_out <= VN_sign_out( 2975 downto 2970 );
    VN496_data_out <= VN_data_out( 2981 downto 2976 );
    VN496_sign_out <= VN_sign_out( 2981 downto 2976 );
    VN497_data_out <= VN_data_out( 2987 downto 2982 );
    VN497_sign_out <= VN_sign_out( 2987 downto 2982 );
    VN498_data_out <= VN_data_out( 2993 downto 2988 );
    VN498_sign_out <= VN_sign_out( 2993 downto 2988 );
    VN499_data_out <= VN_data_out( 2999 downto 2994 );
    VN499_sign_out <= VN_sign_out( 2999 downto 2994 );
    VN500_data_out <= VN_data_out( 3005 downto 3000 );
    VN500_sign_out <= VN_sign_out( 3005 downto 3000 );
    VN501_data_out <= VN_data_out( 3011 downto 3006 );
    VN501_sign_out <= VN_sign_out( 3011 downto 3006 );
    VN502_data_out <= VN_data_out( 3017 downto 3012 );
    VN502_sign_out <= VN_sign_out( 3017 downto 3012 );
    VN503_data_out <= VN_data_out( 3023 downto 3018 );
    VN503_sign_out <= VN_sign_out( 3023 downto 3018 );
    VN504_data_out <= VN_data_out( 3029 downto 3024 );
    VN504_sign_out <= VN_sign_out( 3029 downto 3024 );
    VN505_data_out <= VN_data_out( 3035 downto 3030 );
    VN505_sign_out <= VN_sign_out( 3035 downto 3030 );
    VN506_data_out <= VN_data_out( 3041 downto 3036 );
    VN506_sign_out <= VN_sign_out( 3041 downto 3036 );
    VN507_data_out <= VN_data_out( 3047 downto 3042 );
    VN507_sign_out <= VN_sign_out( 3047 downto 3042 );
    VN508_data_out <= VN_data_out( 3053 downto 3048 );
    VN508_sign_out <= VN_sign_out( 3053 downto 3048 );
    VN509_data_out <= VN_data_out( 3059 downto 3054 );
    VN509_sign_out <= VN_sign_out( 3059 downto 3054 );
    VN510_data_out <= VN_data_out( 3065 downto 3060 );
    VN510_sign_out <= VN_sign_out( 3065 downto 3060 );
    VN511_data_out <= VN_data_out( 3071 downto 3066 );
    VN511_sign_out <= VN_sign_out( 3071 downto 3066 );
    VN512_data_out <= VN_data_out( 3077 downto 3072 );
    VN512_sign_out <= VN_sign_out( 3077 downto 3072 );
    VN513_data_out <= VN_data_out( 3083 downto 3078 );
    VN513_sign_out <= VN_sign_out( 3083 downto 3078 );
    VN514_data_out <= VN_data_out( 3089 downto 3084 );
    VN514_sign_out <= VN_sign_out( 3089 downto 3084 );
    VN515_data_out <= VN_data_out( 3095 downto 3090 );
    VN515_sign_out <= VN_sign_out( 3095 downto 3090 );
    VN516_data_out <= VN_data_out( 3101 downto 3096 );
    VN516_sign_out <= VN_sign_out( 3101 downto 3096 );
    VN517_data_out <= VN_data_out( 3107 downto 3102 );
    VN517_sign_out <= VN_sign_out( 3107 downto 3102 );
    VN518_data_out <= VN_data_out( 3113 downto 3108 );
    VN518_sign_out <= VN_sign_out( 3113 downto 3108 );
    VN519_data_out <= VN_data_out( 3119 downto 3114 );
    VN519_sign_out <= VN_sign_out( 3119 downto 3114 );
    VN520_data_out <= VN_data_out( 3125 downto 3120 );
    VN520_sign_out <= VN_sign_out( 3125 downto 3120 );
    VN521_data_out <= VN_data_out( 3131 downto 3126 );
    VN521_sign_out <= VN_sign_out( 3131 downto 3126 );
    VN522_data_out <= VN_data_out( 3137 downto 3132 );
    VN522_sign_out <= VN_sign_out( 3137 downto 3132 );
    VN523_data_out <= VN_data_out( 3143 downto 3138 );
    VN523_sign_out <= VN_sign_out( 3143 downto 3138 );
    VN524_data_out <= VN_data_out( 3149 downto 3144 );
    VN524_sign_out <= VN_sign_out( 3149 downto 3144 );
    VN525_data_out <= VN_data_out( 3155 downto 3150 );
    VN525_sign_out <= VN_sign_out( 3155 downto 3150 );
    VN526_data_out <= VN_data_out( 3161 downto 3156 );
    VN526_sign_out <= VN_sign_out( 3161 downto 3156 );
    VN527_data_out <= VN_data_out( 3167 downto 3162 );
    VN527_sign_out <= VN_sign_out( 3167 downto 3162 );
    VN528_data_out <= VN_data_out( 3173 downto 3168 );
    VN528_sign_out <= VN_sign_out( 3173 downto 3168 );
    VN529_data_out <= VN_data_out( 3179 downto 3174 );
    VN529_sign_out <= VN_sign_out( 3179 downto 3174 );
    VN530_data_out <= VN_data_out( 3185 downto 3180 );
    VN530_sign_out <= VN_sign_out( 3185 downto 3180 );
    VN531_data_out <= VN_data_out( 3191 downto 3186 );
    VN531_sign_out <= VN_sign_out( 3191 downto 3186 );
    VN532_data_out <= VN_data_out( 3197 downto 3192 );
    VN532_sign_out <= VN_sign_out( 3197 downto 3192 );
    VN533_data_out <= VN_data_out( 3203 downto 3198 );
    VN533_sign_out <= VN_sign_out( 3203 downto 3198 );
    VN534_data_out <= VN_data_out( 3209 downto 3204 );
    VN534_sign_out <= VN_sign_out( 3209 downto 3204 );
    VN535_data_out <= VN_data_out( 3215 downto 3210 );
    VN535_sign_out <= VN_sign_out( 3215 downto 3210 );
    VN536_data_out <= VN_data_out( 3221 downto 3216 );
    VN536_sign_out <= VN_sign_out( 3221 downto 3216 );
    VN537_data_out <= VN_data_out( 3227 downto 3222 );
    VN537_sign_out <= VN_sign_out( 3227 downto 3222 );
    VN538_data_out <= VN_data_out( 3233 downto 3228 );
    VN538_sign_out <= VN_sign_out( 3233 downto 3228 );
    VN539_data_out <= VN_data_out( 3239 downto 3234 );
    VN539_sign_out <= VN_sign_out( 3239 downto 3234 );
    VN540_data_out <= VN_data_out( 3245 downto 3240 );
    VN540_sign_out <= VN_sign_out( 3245 downto 3240 );
    VN541_data_out <= VN_data_out( 3251 downto 3246 );
    VN541_sign_out <= VN_sign_out( 3251 downto 3246 );
    VN542_data_out <= VN_data_out( 3257 downto 3252 );
    VN542_sign_out <= VN_sign_out( 3257 downto 3252 );
    VN543_data_out <= VN_data_out( 3263 downto 3258 );
    VN543_sign_out <= VN_sign_out( 3263 downto 3258 );
    VN544_data_out <= VN_data_out( 3269 downto 3264 );
    VN544_sign_out <= VN_sign_out( 3269 downto 3264 );
    VN545_data_out <= VN_data_out( 3275 downto 3270 );
    VN545_sign_out <= VN_sign_out( 3275 downto 3270 );
    VN546_data_out <= VN_data_out( 3281 downto 3276 );
    VN546_sign_out <= VN_sign_out( 3281 downto 3276 );
    VN547_data_out <= VN_data_out( 3287 downto 3282 );
    VN547_sign_out <= VN_sign_out( 3287 downto 3282 );
    VN548_data_out <= VN_data_out( 3293 downto 3288 );
    VN548_sign_out <= VN_sign_out( 3293 downto 3288 );
    VN549_data_out <= VN_data_out( 3299 downto 3294 );
    VN549_sign_out <= VN_sign_out( 3299 downto 3294 );
    VN550_data_out <= VN_data_out( 3305 downto 3300 );
    VN550_sign_out <= VN_sign_out( 3305 downto 3300 );
    VN551_data_out <= VN_data_out( 3311 downto 3306 );
    VN551_sign_out <= VN_sign_out( 3311 downto 3306 );
    VN552_data_out <= VN_data_out( 3317 downto 3312 );
    VN552_sign_out <= VN_sign_out( 3317 downto 3312 );
    VN553_data_out <= VN_data_out( 3323 downto 3318 );
    VN553_sign_out <= VN_sign_out( 3323 downto 3318 );
    VN554_data_out <= VN_data_out( 3329 downto 3324 );
    VN554_sign_out <= VN_sign_out( 3329 downto 3324 );
    VN555_data_out <= VN_data_out( 3335 downto 3330 );
    VN555_sign_out <= VN_sign_out( 3335 downto 3330 );
    VN556_data_out <= VN_data_out( 3341 downto 3336 );
    VN556_sign_out <= VN_sign_out( 3341 downto 3336 );
    VN557_data_out <= VN_data_out( 3347 downto 3342 );
    VN557_sign_out <= VN_sign_out( 3347 downto 3342 );
    VN558_data_out <= VN_data_out( 3353 downto 3348 );
    VN558_sign_out <= VN_sign_out( 3353 downto 3348 );
    VN559_data_out <= VN_data_out( 3359 downto 3354 );
    VN559_sign_out <= VN_sign_out( 3359 downto 3354 );
    VN560_data_out <= VN_data_out( 3365 downto 3360 );
    VN560_sign_out <= VN_sign_out( 3365 downto 3360 );
    VN561_data_out <= VN_data_out( 3371 downto 3366 );
    VN561_sign_out <= VN_sign_out( 3371 downto 3366 );
    VN562_data_out <= VN_data_out( 3377 downto 3372 );
    VN562_sign_out <= VN_sign_out( 3377 downto 3372 );
    VN563_data_out <= VN_data_out( 3383 downto 3378 );
    VN563_sign_out <= VN_sign_out( 3383 downto 3378 );
    VN564_data_out <= VN_data_out( 3389 downto 3384 );
    VN564_sign_out <= VN_sign_out( 3389 downto 3384 );
    VN565_data_out <= VN_data_out( 3395 downto 3390 );
    VN565_sign_out <= VN_sign_out( 3395 downto 3390 );
    VN566_data_out <= VN_data_out( 3401 downto 3396 );
    VN566_sign_out <= VN_sign_out( 3401 downto 3396 );
    VN567_data_out <= VN_data_out( 3407 downto 3402 );
    VN567_sign_out <= VN_sign_out( 3407 downto 3402 );
    VN568_data_out <= VN_data_out( 3413 downto 3408 );
    VN568_sign_out <= VN_sign_out( 3413 downto 3408 );
    VN569_data_out <= VN_data_out( 3419 downto 3414 );
    VN569_sign_out <= VN_sign_out( 3419 downto 3414 );
    VN570_data_out <= VN_data_out( 3425 downto 3420 );
    VN570_sign_out <= VN_sign_out( 3425 downto 3420 );
    VN571_data_out <= VN_data_out( 3431 downto 3426 );
    VN571_sign_out <= VN_sign_out( 3431 downto 3426 );
    VN572_data_out <= VN_data_out( 3437 downto 3432 );
    VN572_sign_out <= VN_sign_out( 3437 downto 3432 );
    VN573_data_out <= VN_data_out( 3443 downto 3438 );
    VN573_sign_out <= VN_sign_out( 3443 downto 3438 );
    VN574_data_out <= VN_data_out( 3449 downto 3444 );
    VN574_sign_out <= VN_sign_out( 3449 downto 3444 );
    VN575_data_out <= VN_data_out( 3455 downto 3450 );
    VN575_sign_out <= VN_sign_out( 3455 downto 3450 );
    VN576_data_out <= VN_data_out( 3461 downto 3456 );
    VN576_sign_out <= VN_sign_out( 3461 downto 3456 );
    VN577_data_out <= VN_data_out( 3467 downto 3462 );
    VN577_sign_out <= VN_sign_out( 3467 downto 3462 );
    VN578_data_out <= VN_data_out( 3473 downto 3468 );
    VN578_sign_out <= VN_sign_out( 3473 downto 3468 );
    VN579_data_out <= VN_data_out( 3479 downto 3474 );
    VN579_sign_out <= VN_sign_out( 3479 downto 3474 );
    VN580_data_out <= VN_data_out( 3485 downto 3480 );
    VN580_sign_out <= VN_sign_out( 3485 downto 3480 );
    VN581_data_out <= VN_data_out( 3491 downto 3486 );
    VN581_sign_out <= VN_sign_out( 3491 downto 3486 );
    VN582_data_out <= VN_data_out( 3497 downto 3492 );
    VN582_sign_out <= VN_sign_out( 3497 downto 3492 );
    VN583_data_out <= VN_data_out( 3503 downto 3498 );
    VN583_sign_out <= VN_sign_out( 3503 downto 3498 );
    VN584_data_out <= VN_data_out( 3509 downto 3504 );
    VN584_sign_out <= VN_sign_out( 3509 downto 3504 );
    VN585_data_out <= VN_data_out( 3515 downto 3510 );
    VN585_sign_out <= VN_sign_out( 3515 downto 3510 );
    VN586_data_out <= VN_data_out( 3521 downto 3516 );
    VN586_sign_out <= VN_sign_out( 3521 downto 3516 );
    VN587_data_out <= VN_data_out( 3527 downto 3522 );
    VN587_sign_out <= VN_sign_out( 3527 downto 3522 );
    VN588_data_out <= VN_data_out( 3533 downto 3528 );
    VN588_sign_out <= VN_sign_out( 3533 downto 3528 );
    VN589_data_out <= VN_data_out( 3539 downto 3534 );
    VN589_sign_out <= VN_sign_out( 3539 downto 3534 );
    VN590_data_out <= VN_data_out( 3545 downto 3540 );
    VN590_sign_out <= VN_sign_out( 3545 downto 3540 );
    VN591_data_out <= VN_data_out( 3551 downto 3546 );
    VN591_sign_out <= VN_sign_out( 3551 downto 3546 );
    VN592_data_out <= VN_data_out( 3557 downto 3552 );
    VN592_sign_out <= VN_sign_out( 3557 downto 3552 );
    VN593_data_out <= VN_data_out( 3563 downto 3558 );
    VN593_sign_out <= VN_sign_out( 3563 downto 3558 );
    VN594_data_out <= VN_data_out( 3569 downto 3564 );
    VN594_sign_out <= VN_sign_out( 3569 downto 3564 );
    VN595_data_out <= VN_data_out( 3575 downto 3570 );
    VN595_sign_out <= VN_sign_out( 3575 downto 3570 );
    VN596_data_out <= VN_data_out( 3581 downto 3576 );
    VN596_sign_out <= VN_sign_out( 3581 downto 3576 );
    VN597_data_out <= VN_data_out( 3587 downto 3582 );
    VN597_sign_out <= VN_sign_out( 3587 downto 3582 );
    VN598_data_out <= VN_data_out( 3593 downto 3588 );
    VN598_sign_out <= VN_sign_out( 3593 downto 3588 );
    VN599_data_out <= VN_data_out( 3599 downto 3594 );
    VN599_sign_out <= VN_sign_out( 3599 downto 3594 );
    VN600_data_out <= VN_data_out( 3605 downto 3600 );
    VN600_sign_out <= VN_sign_out( 3605 downto 3600 );
    VN601_data_out <= VN_data_out( 3611 downto 3606 );
    VN601_sign_out <= VN_sign_out( 3611 downto 3606 );
    VN602_data_out <= VN_data_out( 3617 downto 3612 );
    VN602_sign_out <= VN_sign_out( 3617 downto 3612 );
    VN603_data_out <= VN_data_out( 3623 downto 3618 );
    VN603_sign_out <= VN_sign_out( 3623 downto 3618 );
    VN604_data_out <= VN_data_out( 3629 downto 3624 );
    VN604_sign_out <= VN_sign_out( 3629 downto 3624 );
    VN605_data_out <= VN_data_out( 3635 downto 3630 );
    VN605_sign_out <= VN_sign_out( 3635 downto 3630 );
    VN606_data_out <= VN_data_out( 3641 downto 3636 );
    VN606_sign_out <= VN_sign_out( 3641 downto 3636 );
    VN607_data_out <= VN_data_out( 3647 downto 3642 );
    VN607_sign_out <= VN_sign_out( 3647 downto 3642 );
    VN608_data_out <= VN_data_out( 3653 downto 3648 );
    VN608_sign_out <= VN_sign_out( 3653 downto 3648 );
    VN609_data_out <= VN_data_out( 3659 downto 3654 );
    VN609_sign_out <= VN_sign_out( 3659 downto 3654 );
    VN610_data_out <= VN_data_out( 3665 downto 3660 );
    VN610_sign_out <= VN_sign_out( 3665 downto 3660 );
    VN611_data_out <= VN_data_out( 3671 downto 3666 );
    VN611_sign_out <= VN_sign_out( 3671 downto 3666 );
    VN612_data_out <= VN_data_out( 3677 downto 3672 );
    VN612_sign_out <= VN_sign_out( 3677 downto 3672 );
    VN613_data_out <= VN_data_out( 3683 downto 3678 );
    VN613_sign_out <= VN_sign_out( 3683 downto 3678 );
    VN614_data_out <= VN_data_out( 3689 downto 3684 );
    VN614_sign_out <= VN_sign_out( 3689 downto 3684 );
    VN615_data_out <= VN_data_out( 3695 downto 3690 );
    VN615_sign_out <= VN_sign_out( 3695 downto 3690 );
    VN616_data_out <= VN_data_out( 3701 downto 3696 );
    VN616_sign_out <= VN_sign_out( 3701 downto 3696 );
    VN617_data_out <= VN_data_out( 3707 downto 3702 );
    VN617_sign_out <= VN_sign_out( 3707 downto 3702 );
    VN618_data_out <= VN_data_out( 3713 downto 3708 );
    VN618_sign_out <= VN_sign_out( 3713 downto 3708 );
    VN619_data_out <= VN_data_out( 3719 downto 3714 );
    VN619_sign_out <= VN_sign_out( 3719 downto 3714 );
    VN620_data_out <= VN_data_out( 3725 downto 3720 );
    VN620_sign_out <= VN_sign_out( 3725 downto 3720 );
    VN621_data_out <= VN_data_out( 3731 downto 3726 );
    VN621_sign_out <= VN_sign_out( 3731 downto 3726 );
    VN622_data_out <= VN_data_out( 3737 downto 3732 );
    VN622_sign_out <= VN_sign_out( 3737 downto 3732 );
    VN623_data_out <= VN_data_out( 3743 downto 3738 );
    VN623_sign_out <= VN_sign_out( 3743 downto 3738 );
    VN624_data_out <= VN_data_out( 3749 downto 3744 );
    VN624_sign_out <= VN_sign_out( 3749 downto 3744 );
    VN625_data_out <= VN_data_out( 3755 downto 3750 );
    VN625_sign_out <= VN_sign_out( 3755 downto 3750 );
    VN626_data_out <= VN_data_out( 3761 downto 3756 );
    VN626_sign_out <= VN_sign_out( 3761 downto 3756 );
    VN627_data_out <= VN_data_out( 3767 downto 3762 );
    VN627_sign_out <= VN_sign_out( 3767 downto 3762 );
    VN628_data_out <= VN_data_out( 3773 downto 3768 );
    VN628_sign_out <= VN_sign_out( 3773 downto 3768 );
    VN629_data_out <= VN_data_out( 3779 downto 3774 );
    VN629_sign_out <= VN_sign_out( 3779 downto 3774 );
    VN630_data_out <= VN_data_out( 3785 downto 3780 );
    VN630_sign_out <= VN_sign_out( 3785 downto 3780 );
    VN631_data_out <= VN_data_out( 3791 downto 3786 );
    VN631_sign_out <= VN_sign_out( 3791 downto 3786 );
    VN632_data_out <= VN_data_out( 3797 downto 3792 );
    VN632_sign_out <= VN_sign_out( 3797 downto 3792 );
    VN633_data_out <= VN_data_out( 3803 downto 3798 );
    VN633_sign_out <= VN_sign_out( 3803 downto 3798 );
    VN634_data_out <= VN_data_out( 3809 downto 3804 );
    VN634_sign_out <= VN_sign_out( 3809 downto 3804 );
    VN635_data_out <= VN_data_out( 3815 downto 3810 );
    VN635_sign_out <= VN_sign_out( 3815 downto 3810 );
    VN636_data_out <= VN_data_out( 3821 downto 3816 );
    VN636_sign_out <= VN_sign_out( 3821 downto 3816 );
    VN637_data_out <= VN_data_out( 3827 downto 3822 );
    VN637_sign_out <= VN_sign_out( 3827 downto 3822 );
    VN638_data_out <= VN_data_out( 3833 downto 3828 );
    VN638_sign_out <= VN_sign_out( 3833 downto 3828 );
    VN639_data_out <= VN_data_out( 3839 downto 3834 );
    VN639_sign_out <= VN_sign_out( 3839 downto 3834 );
    VN640_data_out <= VN_data_out( 3845 downto 3840 );
    VN640_sign_out <= VN_sign_out( 3845 downto 3840 );
    VN641_data_out <= VN_data_out( 3851 downto 3846 );
    VN641_sign_out <= VN_sign_out( 3851 downto 3846 );
    VN642_data_out <= VN_data_out( 3857 downto 3852 );
    VN642_sign_out <= VN_sign_out( 3857 downto 3852 );
    VN643_data_out <= VN_data_out( 3863 downto 3858 );
    VN643_sign_out <= VN_sign_out( 3863 downto 3858 );
    VN644_data_out <= VN_data_out( 3869 downto 3864 );
    VN644_sign_out <= VN_sign_out( 3869 downto 3864 );
    VN645_data_out <= VN_data_out( 3875 downto 3870 );
    VN645_sign_out <= VN_sign_out( 3875 downto 3870 );
    VN646_data_out <= VN_data_out( 3881 downto 3876 );
    VN646_sign_out <= VN_sign_out( 3881 downto 3876 );
    VN647_data_out <= VN_data_out( 3887 downto 3882 );
    VN647_sign_out <= VN_sign_out( 3887 downto 3882 );
    VN648_data_out <= VN_data_out( 3893 downto 3888 );
    VN648_sign_out <= VN_sign_out( 3893 downto 3888 );
    VN649_data_out <= VN_data_out( 3899 downto 3894 );
    VN649_sign_out <= VN_sign_out( 3899 downto 3894 );
    VN650_data_out <= VN_data_out( 3905 downto 3900 );
    VN650_sign_out <= VN_sign_out( 3905 downto 3900 );
    VN651_data_out <= VN_data_out( 3911 downto 3906 );
    VN651_sign_out <= VN_sign_out( 3911 downto 3906 );
    VN652_data_out <= VN_data_out( 3917 downto 3912 );
    VN652_sign_out <= VN_sign_out( 3917 downto 3912 );
    VN653_data_out <= VN_data_out( 3923 downto 3918 );
    VN653_sign_out <= VN_sign_out( 3923 downto 3918 );
    VN654_data_out <= VN_data_out( 3929 downto 3924 );
    VN654_sign_out <= VN_sign_out( 3929 downto 3924 );
    VN655_data_out <= VN_data_out( 3935 downto 3930 );
    VN655_sign_out <= VN_sign_out( 3935 downto 3930 );
    VN656_data_out <= VN_data_out( 3941 downto 3936 );
    VN656_sign_out <= VN_sign_out( 3941 downto 3936 );
    VN657_data_out <= VN_data_out( 3947 downto 3942 );
    VN657_sign_out <= VN_sign_out( 3947 downto 3942 );
    VN658_data_out <= VN_data_out( 3953 downto 3948 );
    VN658_sign_out <= VN_sign_out( 3953 downto 3948 );
    VN659_data_out <= VN_data_out( 3959 downto 3954 );
    VN659_sign_out <= VN_sign_out( 3959 downto 3954 );
    VN660_data_out <= VN_data_out( 3965 downto 3960 );
    VN660_sign_out <= VN_sign_out( 3965 downto 3960 );
    VN661_data_out <= VN_data_out( 3971 downto 3966 );
    VN661_sign_out <= VN_sign_out( 3971 downto 3966 );
    VN662_data_out <= VN_data_out( 3977 downto 3972 );
    VN662_sign_out <= VN_sign_out( 3977 downto 3972 );
    VN663_data_out <= VN_data_out( 3983 downto 3978 );
    VN663_sign_out <= VN_sign_out( 3983 downto 3978 );
    VN664_data_out <= VN_data_out( 3989 downto 3984 );
    VN664_sign_out <= VN_sign_out( 3989 downto 3984 );
    VN665_data_out <= VN_data_out( 3995 downto 3990 );
    VN665_sign_out <= VN_sign_out( 3995 downto 3990 );
    VN666_data_out <= VN_data_out( 4001 downto 3996 );
    VN666_sign_out <= VN_sign_out( 4001 downto 3996 );
    VN667_data_out <= VN_data_out( 4007 downto 4002 );
    VN667_sign_out <= VN_sign_out( 4007 downto 4002 );
    VN668_data_out <= VN_data_out( 4013 downto 4008 );
    VN668_sign_out <= VN_sign_out( 4013 downto 4008 );
    VN669_data_out <= VN_data_out( 4019 downto 4014 );
    VN669_sign_out <= VN_sign_out( 4019 downto 4014 );
    VN670_data_out <= VN_data_out( 4025 downto 4020 );
    VN670_sign_out <= VN_sign_out( 4025 downto 4020 );
    VN671_data_out <= VN_data_out( 4031 downto 4026 );
    VN671_sign_out <= VN_sign_out( 4031 downto 4026 );
    VN672_data_out <= VN_data_out( 4037 downto 4032 );
    VN672_sign_out <= VN_sign_out( 4037 downto 4032 );
    VN673_data_out <= VN_data_out( 4043 downto 4038 );
    VN673_sign_out <= VN_sign_out( 4043 downto 4038 );
    VN674_data_out <= VN_data_out( 4049 downto 4044 );
    VN674_sign_out <= VN_sign_out( 4049 downto 4044 );
    VN675_data_out <= VN_data_out( 4055 downto 4050 );
    VN675_sign_out <= VN_sign_out( 4055 downto 4050 );
    VN676_data_out <= VN_data_out( 4061 downto 4056 );
    VN676_sign_out <= VN_sign_out( 4061 downto 4056 );
    VN677_data_out <= VN_data_out( 4067 downto 4062 );
    VN677_sign_out <= VN_sign_out( 4067 downto 4062 );
    VN678_data_out <= VN_data_out( 4073 downto 4068 );
    VN678_sign_out <= VN_sign_out( 4073 downto 4068 );
    VN679_data_out <= VN_data_out( 4079 downto 4074 );
    VN679_sign_out <= VN_sign_out( 4079 downto 4074 );
    VN680_data_out <= VN_data_out( 4085 downto 4080 );
    VN680_sign_out <= VN_sign_out( 4085 downto 4080 );
    VN681_data_out <= VN_data_out( 4091 downto 4086 );
    VN681_sign_out <= VN_sign_out( 4091 downto 4086 );
    VN682_data_out <= VN_data_out( 4097 downto 4092 );
    VN682_sign_out <= VN_sign_out( 4097 downto 4092 );
    VN683_data_out <= VN_data_out( 4103 downto 4098 );
    VN683_sign_out <= VN_sign_out( 4103 downto 4098 );
    VN684_data_out <= VN_data_out( 4109 downto 4104 );
    VN684_sign_out <= VN_sign_out( 4109 downto 4104 );
    VN685_data_out <= VN_data_out( 4115 downto 4110 );
    VN685_sign_out <= VN_sign_out( 4115 downto 4110 );
    VN686_data_out <= VN_data_out( 4121 downto 4116 );
    VN686_sign_out <= VN_sign_out( 4121 downto 4116 );
    VN687_data_out <= VN_data_out( 4127 downto 4122 );
    VN687_sign_out <= VN_sign_out( 4127 downto 4122 );
    VN688_data_out <= VN_data_out( 4133 downto 4128 );
    VN688_sign_out <= VN_sign_out( 4133 downto 4128 );
    VN689_data_out <= VN_data_out( 4139 downto 4134 );
    VN689_sign_out <= VN_sign_out( 4139 downto 4134 );
    VN690_data_out <= VN_data_out( 4145 downto 4140 );
    VN690_sign_out <= VN_sign_out( 4145 downto 4140 );
    VN691_data_out <= VN_data_out( 4151 downto 4146 );
    VN691_sign_out <= VN_sign_out( 4151 downto 4146 );
    VN692_data_out <= VN_data_out( 4157 downto 4152 );
    VN692_sign_out <= VN_sign_out( 4157 downto 4152 );
    VN693_data_out <= VN_data_out( 4163 downto 4158 );
    VN693_sign_out <= VN_sign_out( 4163 downto 4158 );
    VN694_data_out <= VN_data_out( 4169 downto 4164 );
    VN694_sign_out <= VN_sign_out( 4169 downto 4164 );
    VN695_data_out <= VN_data_out( 4175 downto 4170 );
    VN695_sign_out <= VN_sign_out( 4175 downto 4170 );
    VN696_data_out <= VN_data_out( 4181 downto 4176 );
    VN696_sign_out <= VN_sign_out( 4181 downto 4176 );
    VN697_data_out <= VN_data_out( 4187 downto 4182 );
    VN697_sign_out <= VN_sign_out( 4187 downto 4182 );
    VN698_data_out <= VN_data_out( 4193 downto 4188 );
    VN698_sign_out <= VN_sign_out( 4193 downto 4188 );
    VN699_data_out <= VN_data_out( 4199 downto 4194 );
    VN699_sign_out <= VN_sign_out( 4199 downto 4194 );
    VN700_data_out <= VN_data_out( 4205 downto 4200 );
    VN700_sign_out <= VN_sign_out( 4205 downto 4200 );
    VN701_data_out <= VN_data_out( 4211 downto 4206 );
    VN701_sign_out <= VN_sign_out( 4211 downto 4206 );
    VN702_data_out <= VN_data_out( 4217 downto 4212 );
    VN702_sign_out <= VN_sign_out( 4217 downto 4212 );
    VN703_data_out <= VN_data_out( 4223 downto 4218 );
    VN703_sign_out <= VN_sign_out( 4223 downto 4218 );
    VN704_data_out <= VN_data_out( 4229 downto 4224 );
    VN704_sign_out <= VN_sign_out( 4229 downto 4224 );
    VN705_data_out <= VN_data_out( 4235 downto 4230 );
    VN705_sign_out <= VN_sign_out( 4235 downto 4230 );
    VN706_data_out <= VN_data_out( 4241 downto 4236 );
    VN706_sign_out <= VN_sign_out( 4241 downto 4236 );
    VN707_data_out <= VN_data_out( 4247 downto 4242 );
    VN707_sign_out <= VN_sign_out( 4247 downto 4242 );
    VN708_data_out <= VN_data_out( 4253 downto 4248 );
    VN708_sign_out <= VN_sign_out( 4253 downto 4248 );
    VN709_data_out <= VN_data_out( 4259 downto 4254 );
    VN709_sign_out <= VN_sign_out( 4259 downto 4254 );
    VN710_data_out <= VN_data_out( 4265 downto 4260 );
    VN710_sign_out <= VN_sign_out( 4265 downto 4260 );
    VN711_data_out <= VN_data_out( 4271 downto 4266 );
    VN711_sign_out <= VN_sign_out( 4271 downto 4266 );
    VN712_data_out <= VN_data_out( 4277 downto 4272 );
    VN712_sign_out <= VN_sign_out( 4277 downto 4272 );
    VN713_data_out <= VN_data_out( 4283 downto 4278 );
    VN713_sign_out <= VN_sign_out( 4283 downto 4278 );
    VN714_data_out <= VN_data_out( 4289 downto 4284 );
    VN714_sign_out <= VN_sign_out( 4289 downto 4284 );
    VN715_data_out <= VN_data_out( 4295 downto 4290 );
    VN715_sign_out <= VN_sign_out( 4295 downto 4290 );
    VN716_data_out <= VN_data_out( 4301 downto 4296 );
    VN716_sign_out <= VN_sign_out( 4301 downto 4296 );
    VN717_data_out <= VN_data_out( 4307 downto 4302 );
    VN717_sign_out <= VN_sign_out( 4307 downto 4302 );
    VN718_data_out <= VN_data_out( 4313 downto 4308 );
    VN718_sign_out <= VN_sign_out( 4313 downto 4308 );
    VN719_data_out <= VN_data_out( 4319 downto 4314 );
    VN719_sign_out <= VN_sign_out( 4319 downto 4314 );
    VN720_data_out <= VN_data_out( 4325 downto 4320 );
    VN720_sign_out <= VN_sign_out( 4325 downto 4320 );
    VN721_data_out <= VN_data_out( 4331 downto 4326 );
    VN721_sign_out <= VN_sign_out( 4331 downto 4326 );
    VN722_data_out <= VN_data_out( 4337 downto 4332 );
    VN722_sign_out <= VN_sign_out( 4337 downto 4332 );
    VN723_data_out <= VN_data_out( 4343 downto 4338 );
    VN723_sign_out <= VN_sign_out( 4343 downto 4338 );
    VN724_data_out <= VN_data_out( 4349 downto 4344 );
    VN724_sign_out <= VN_sign_out( 4349 downto 4344 );
    VN725_data_out <= VN_data_out( 4355 downto 4350 );
    VN725_sign_out <= VN_sign_out( 4355 downto 4350 );
    VN726_data_out <= VN_data_out( 4361 downto 4356 );
    VN726_sign_out <= VN_sign_out( 4361 downto 4356 );
    VN727_data_out <= VN_data_out( 4367 downto 4362 );
    VN727_sign_out <= VN_sign_out( 4367 downto 4362 );
    VN728_data_out <= VN_data_out( 4373 downto 4368 );
    VN728_sign_out <= VN_sign_out( 4373 downto 4368 );
    VN729_data_out <= VN_data_out( 4379 downto 4374 );
    VN729_sign_out <= VN_sign_out( 4379 downto 4374 );
    VN730_data_out <= VN_data_out( 4385 downto 4380 );
    VN730_sign_out <= VN_sign_out( 4385 downto 4380 );
    VN731_data_out <= VN_data_out( 4391 downto 4386 );
    VN731_sign_out <= VN_sign_out( 4391 downto 4386 );
    VN732_data_out <= VN_data_out( 4397 downto 4392 );
    VN732_sign_out <= VN_sign_out( 4397 downto 4392 );
    VN733_data_out <= VN_data_out( 4403 downto 4398 );
    VN733_sign_out <= VN_sign_out( 4403 downto 4398 );
    VN734_data_out <= VN_data_out( 4409 downto 4404 );
    VN734_sign_out <= VN_sign_out( 4409 downto 4404 );
    VN735_data_out <= VN_data_out( 4415 downto 4410 );
    VN735_sign_out <= VN_sign_out( 4415 downto 4410 );
    VN736_data_out <= VN_data_out( 4421 downto 4416 );
    VN736_sign_out <= VN_sign_out( 4421 downto 4416 );
    VN737_data_out <= VN_data_out( 4427 downto 4422 );
    VN737_sign_out <= VN_sign_out( 4427 downto 4422 );
    VN738_data_out <= VN_data_out( 4433 downto 4428 );
    VN738_sign_out <= VN_sign_out( 4433 downto 4428 );
    VN739_data_out <= VN_data_out( 4439 downto 4434 );
    VN739_sign_out <= VN_sign_out( 4439 downto 4434 );
    VN740_data_out <= VN_data_out( 4445 downto 4440 );
    VN740_sign_out <= VN_sign_out( 4445 downto 4440 );
    VN741_data_out <= VN_data_out( 4451 downto 4446 );
    VN741_sign_out <= VN_sign_out( 4451 downto 4446 );
    VN742_data_out <= VN_data_out( 4457 downto 4452 );
    VN742_sign_out <= VN_sign_out( 4457 downto 4452 );
    VN743_data_out <= VN_data_out( 4463 downto 4458 );
    VN743_sign_out <= VN_sign_out( 4463 downto 4458 );
    VN744_data_out <= VN_data_out( 4469 downto 4464 );
    VN744_sign_out <= VN_sign_out( 4469 downto 4464 );
    VN745_data_out <= VN_data_out( 4475 downto 4470 );
    VN745_sign_out <= VN_sign_out( 4475 downto 4470 );
    VN746_data_out <= VN_data_out( 4481 downto 4476 );
    VN746_sign_out <= VN_sign_out( 4481 downto 4476 );
    VN747_data_out <= VN_data_out( 4487 downto 4482 );
    VN747_sign_out <= VN_sign_out( 4487 downto 4482 );
    VN748_data_out <= VN_data_out( 4493 downto 4488 );
    VN748_sign_out <= VN_sign_out( 4493 downto 4488 );
    VN749_data_out <= VN_data_out( 4499 downto 4494 );
    VN749_sign_out <= VN_sign_out( 4499 downto 4494 );
    VN750_data_out <= VN_data_out( 4505 downto 4500 );
    VN750_sign_out <= VN_sign_out( 4505 downto 4500 );
    VN751_data_out <= VN_data_out( 4511 downto 4506 );
    VN751_sign_out <= VN_sign_out( 4511 downto 4506 );
    VN752_data_out <= VN_data_out( 4517 downto 4512 );
    VN752_sign_out <= VN_sign_out( 4517 downto 4512 );
    VN753_data_out <= VN_data_out( 4523 downto 4518 );
    VN753_sign_out <= VN_sign_out( 4523 downto 4518 );
    VN754_data_out <= VN_data_out( 4529 downto 4524 );
    VN754_sign_out <= VN_sign_out( 4529 downto 4524 );
    VN755_data_out <= VN_data_out( 4535 downto 4530 );
    VN755_sign_out <= VN_sign_out( 4535 downto 4530 );
    VN756_data_out <= VN_data_out( 4541 downto 4536 );
    VN756_sign_out <= VN_sign_out( 4541 downto 4536 );
    VN757_data_out <= VN_data_out( 4547 downto 4542 );
    VN757_sign_out <= VN_sign_out( 4547 downto 4542 );
    VN758_data_out <= VN_data_out( 4553 downto 4548 );
    VN758_sign_out <= VN_sign_out( 4553 downto 4548 );
    VN759_data_out <= VN_data_out( 4559 downto 4554 );
    VN759_sign_out <= VN_sign_out( 4559 downto 4554 );
    VN760_data_out <= VN_data_out( 4565 downto 4560 );
    VN760_sign_out <= VN_sign_out( 4565 downto 4560 );
    VN761_data_out <= VN_data_out( 4571 downto 4566 );
    VN761_sign_out <= VN_sign_out( 4571 downto 4566 );
    VN762_data_out <= VN_data_out( 4577 downto 4572 );
    VN762_sign_out <= VN_sign_out( 4577 downto 4572 );
    VN763_data_out <= VN_data_out( 4583 downto 4578 );
    VN763_sign_out <= VN_sign_out( 4583 downto 4578 );
    VN764_data_out <= VN_data_out( 4589 downto 4584 );
    VN764_sign_out <= VN_sign_out( 4589 downto 4584 );
    VN765_data_out <= VN_data_out( 4595 downto 4590 );
    VN765_sign_out <= VN_sign_out( 4595 downto 4590 );
    VN766_data_out <= VN_data_out( 4601 downto 4596 );
    VN766_sign_out <= VN_sign_out( 4601 downto 4596 );
    VN767_data_out <= VN_data_out( 4607 downto 4602 );
    VN767_sign_out <= VN_sign_out( 4607 downto 4602 );
    VN768_data_out <= VN_data_out( 4613 downto 4608 );
    VN768_sign_out <= VN_sign_out( 4613 downto 4608 );
    VN769_data_out <= VN_data_out( 4619 downto 4614 );
    VN769_sign_out <= VN_sign_out( 4619 downto 4614 );
    VN770_data_out <= VN_data_out( 4625 downto 4620 );
    VN770_sign_out <= VN_sign_out( 4625 downto 4620 );
    VN771_data_out <= VN_data_out( 4631 downto 4626 );
    VN771_sign_out <= VN_sign_out( 4631 downto 4626 );
    VN772_data_out <= VN_data_out( 4637 downto 4632 );
    VN772_sign_out <= VN_sign_out( 4637 downto 4632 );
    VN773_data_out <= VN_data_out( 4643 downto 4638 );
    VN773_sign_out <= VN_sign_out( 4643 downto 4638 );
    VN774_data_out <= VN_data_out( 4649 downto 4644 );
    VN774_sign_out <= VN_sign_out( 4649 downto 4644 );
    VN775_data_out <= VN_data_out( 4655 downto 4650 );
    VN775_sign_out <= VN_sign_out( 4655 downto 4650 );
    VN776_data_out <= VN_data_out( 4661 downto 4656 );
    VN776_sign_out <= VN_sign_out( 4661 downto 4656 );
    VN777_data_out <= VN_data_out( 4667 downto 4662 );
    VN777_sign_out <= VN_sign_out( 4667 downto 4662 );
    VN778_data_out <= VN_data_out( 4673 downto 4668 );
    VN778_sign_out <= VN_sign_out( 4673 downto 4668 );
    VN779_data_out <= VN_data_out( 4679 downto 4674 );
    VN779_sign_out <= VN_sign_out( 4679 downto 4674 );
    VN780_data_out <= VN_data_out( 4685 downto 4680 );
    VN780_sign_out <= VN_sign_out( 4685 downto 4680 );
    VN781_data_out <= VN_data_out( 4691 downto 4686 );
    VN781_sign_out <= VN_sign_out( 4691 downto 4686 );
    VN782_data_out <= VN_data_out( 4697 downto 4692 );
    VN782_sign_out <= VN_sign_out( 4697 downto 4692 );
    VN783_data_out <= VN_data_out( 4703 downto 4698 );
    VN783_sign_out <= VN_sign_out( 4703 downto 4698 );
    VN784_data_out <= VN_data_out( 4709 downto 4704 );
    VN784_sign_out <= VN_sign_out( 4709 downto 4704 );
    VN785_data_out <= VN_data_out( 4715 downto 4710 );
    VN785_sign_out <= VN_sign_out( 4715 downto 4710 );
    VN786_data_out <= VN_data_out( 4721 downto 4716 );
    VN786_sign_out <= VN_sign_out( 4721 downto 4716 );
    VN787_data_out <= VN_data_out( 4727 downto 4722 );
    VN787_sign_out <= VN_sign_out( 4727 downto 4722 );
    VN788_data_out <= VN_data_out( 4733 downto 4728 );
    VN788_sign_out <= VN_sign_out( 4733 downto 4728 );
    VN789_data_out <= VN_data_out( 4739 downto 4734 );
    VN789_sign_out <= VN_sign_out( 4739 downto 4734 );
    VN790_data_out <= VN_data_out( 4745 downto 4740 );
    VN790_sign_out <= VN_sign_out( 4745 downto 4740 );
    VN791_data_out <= VN_data_out( 4751 downto 4746 );
    VN791_sign_out <= VN_sign_out( 4751 downto 4746 );
    VN792_data_out <= VN_data_out( 4757 downto 4752 );
    VN792_sign_out <= VN_sign_out( 4757 downto 4752 );
    VN793_data_out <= VN_data_out( 4763 downto 4758 );
    VN793_sign_out <= VN_sign_out( 4763 downto 4758 );
    VN794_data_out <= VN_data_out( 4769 downto 4764 );
    VN794_sign_out <= VN_sign_out( 4769 downto 4764 );
    VN795_data_out <= VN_data_out( 4775 downto 4770 );
    VN795_sign_out <= VN_sign_out( 4775 downto 4770 );
    VN796_data_out <= VN_data_out( 4781 downto 4776 );
    VN796_sign_out <= VN_sign_out( 4781 downto 4776 );
    VN797_data_out <= VN_data_out( 4787 downto 4782 );
    VN797_sign_out <= VN_sign_out( 4787 downto 4782 );
    VN798_data_out <= VN_data_out( 4793 downto 4788 );
    VN798_sign_out <= VN_sign_out( 4793 downto 4788 );
    VN799_data_out <= VN_data_out( 4799 downto 4794 );
    VN799_sign_out <= VN_sign_out( 4799 downto 4794 );
    VN800_data_out <= VN_data_out( 4805 downto 4800 );
    VN800_sign_out <= VN_sign_out( 4805 downto 4800 );
    VN801_data_out <= VN_data_out( 4811 downto 4806 );
    VN801_sign_out <= VN_sign_out( 4811 downto 4806 );
    VN802_data_out <= VN_data_out( 4817 downto 4812 );
    VN802_sign_out <= VN_sign_out( 4817 downto 4812 );
    VN803_data_out <= VN_data_out( 4823 downto 4818 );
    VN803_sign_out <= VN_sign_out( 4823 downto 4818 );
    VN804_data_out <= VN_data_out( 4829 downto 4824 );
    VN804_sign_out <= VN_sign_out( 4829 downto 4824 );
    VN805_data_out <= VN_data_out( 4835 downto 4830 );
    VN805_sign_out <= VN_sign_out( 4835 downto 4830 );
    VN806_data_out <= VN_data_out( 4841 downto 4836 );
    VN806_sign_out <= VN_sign_out( 4841 downto 4836 );
    VN807_data_out <= VN_data_out( 4847 downto 4842 );
    VN807_sign_out <= VN_sign_out( 4847 downto 4842 );
    VN808_data_out <= VN_data_out( 4853 downto 4848 );
    VN808_sign_out <= VN_sign_out( 4853 downto 4848 );
    VN809_data_out <= VN_data_out( 4859 downto 4854 );
    VN809_sign_out <= VN_sign_out( 4859 downto 4854 );
    VN810_data_out <= VN_data_out( 4865 downto 4860 );
    VN810_sign_out <= VN_sign_out( 4865 downto 4860 );
    VN811_data_out <= VN_data_out( 4871 downto 4866 );
    VN811_sign_out <= VN_sign_out( 4871 downto 4866 );
    VN812_data_out <= VN_data_out( 4877 downto 4872 );
    VN812_sign_out <= VN_sign_out( 4877 downto 4872 );
    VN813_data_out <= VN_data_out( 4883 downto 4878 );
    VN813_sign_out <= VN_sign_out( 4883 downto 4878 );
    VN814_data_out <= VN_data_out( 4889 downto 4884 );
    VN814_sign_out <= VN_sign_out( 4889 downto 4884 );
    VN815_data_out <= VN_data_out( 4895 downto 4890 );
    VN815_sign_out <= VN_sign_out( 4895 downto 4890 );
    VN816_data_out <= VN_data_out( 4901 downto 4896 );
    VN816_sign_out <= VN_sign_out( 4901 downto 4896 );
    VN817_data_out <= VN_data_out( 4907 downto 4902 );
    VN817_sign_out <= VN_sign_out( 4907 downto 4902 );
    VN818_data_out <= VN_data_out( 4913 downto 4908 );
    VN818_sign_out <= VN_sign_out( 4913 downto 4908 );
    VN819_data_out <= VN_data_out( 4919 downto 4914 );
    VN819_sign_out <= VN_sign_out( 4919 downto 4914 );
    VN820_data_out <= VN_data_out( 4925 downto 4920 );
    VN820_sign_out <= VN_sign_out( 4925 downto 4920 );
    VN821_data_out <= VN_data_out( 4931 downto 4926 );
    VN821_sign_out <= VN_sign_out( 4931 downto 4926 );
    VN822_data_out <= VN_data_out( 4937 downto 4932 );
    VN822_sign_out <= VN_sign_out( 4937 downto 4932 );
    VN823_data_out <= VN_data_out( 4943 downto 4938 );
    VN823_sign_out <= VN_sign_out( 4943 downto 4938 );
    VN824_data_out <= VN_data_out( 4949 downto 4944 );
    VN824_sign_out <= VN_sign_out( 4949 downto 4944 );
    VN825_data_out <= VN_data_out( 4955 downto 4950 );
    VN825_sign_out <= VN_sign_out( 4955 downto 4950 );
    VN826_data_out <= VN_data_out( 4961 downto 4956 );
    VN826_sign_out <= VN_sign_out( 4961 downto 4956 );
    VN827_data_out <= VN_data_out( 4967 downto 4962 );
    VN827_sign_out <= VN_sign_out( 4967 downto 4962 );
    VN828_data_out <= VN_data_out( 4973 downto 4968 );
    VN828_sign_out <= VN_sign_out( 4973 downto 4968 );
    VN829_data_out <= VN_data_out( 4979 downto 4974 );
    VN829_sign_out <= VN_sign_out( 4979 downto 4974 );
    VN830_data_out <= VN_data_out( 4985 downto 4980 );
    VN830_sign_out <= VN_sign_out( 4985 downto 4980 );
    VN831_data_out <= VN_data_out( 4991 downto 4986 );
    VN831_sign_out <= VN_sign_out( 4991 downto 4986 );
    VN832_data_out <= VN_data_out( 4997 downto 4992 );
    VN832_sign_out <= VN_sign_out( 4997 downto 4992 );
    VN833_data_out <= VN_data_out( 5003 downto 4998 );
    VN833_sign_out <= VN_sign_out( 5003 downto 4998 );
    VN834_data_out <= VN_data_out( 5009 downto 5004 );
    VN834_sign_out <= VN_sign_out( 5009 downto 5004 );
    VN835_data_out <= VN_data_out( 5015 downto 5010 );
    VN835_sign_out <= VN_sign_out( 5015 downto 5010 );
    VN836_data_out <= VN_data_out( 5021 downto 5016 );
    VN836_sign_out <= VN_sign_out( 5021 downto 5016 );
    VN837_data_out <= VN_data_out( 5027 downto 5022 );
    VN837_sign_out <= VN_sign_out( 5027 downto 5022 );
    VN838_data_out <= VN_data_out( 5033 downto 5028 );
    VN838_sign_out <= VN_sign_out( 5033 downto 5028 );
    VN839_data_out <= VN_data_out( 5039 downto 5034 );
    VN839_sign_out <= VN_sign_out( 5039 downto 5034 );
    VN840_data_out <= VN_data_out( 5045 downto 5040 );
    VN840_sign_out <= VN_sign_out( 5045 downto 5040 );
    VN841_data_out <= VN_data_out( 5051 downto 5046 );
    VN841_sign_out <= VN_sign_out( 5051 downto 5046 );
    VN842_data_out <= VN_data_out( 5057 downto 5052 );
    VN842_sign_out <= VN_sign_out( 5057 downto 5052 );
    VN843_data_out <= VN_data_out( 5063 downto 5058 );
    VN843_sign_out <= VN_sign_out( 5063 downto 5058 );
    VN844_data_out <= VN_data_out( 5069 downto 5064 );
    VN844_sign_out <= VN_sign_out( 5069 downto 5064 );
    VN845_data_out <= VN_data_out( 5075 downto 5070 );
    VN845_sign_out <= VN_sign_out( 5075 downto 5070 );
    VN846_data_out <= VN_data_out( 5081 downto 5076 );
    VN846_sign_out <= VN_sign_out( 5081 downto 5076 );
    VN847_data_out <= VN_data_out( 5087 downto 5082 );
    VN847_sign_out <= VN_sign_out( 5087 downto 5082 );
    VN848_data_out <= VN_data_out( 5093 downto 5088 );
    VN848_sign_out <= VN_sign_out( 5093 downto 5088 );
    VN849_data_out <= VN_data_out( 5099 downto 5094 );
    VN849_sign_out <= VN_sign_out( 5099 downto 5094 );
    VN850_data_out <= VN_data_out( 5105 downto 5100 );
    VN850_sign_out <= VN_sign_out( 5105 downto 5100 );
    VN851_data_out <= VN_data_out( 5111 downto 5106 );
    VN851_sign_out <= VN_sign_out( 5111 downto 5106 );
    VN852_data_out <= VN_data_out( 5117 downto 5112 );
    VN852_sign_out <= VN_sign_out( 5117 downto 5112 );
    VN853_data_out <= VN_data_out( 5123 downto 5118 );
    VN853_sign_out <= VN_sign_out( 5123 downto 5118 );
    VN854_data_out <= VN_data_out( 5129 downto 5124 );
    VN854_sign_out <= VN_sign_out( 5129 downto 5124 );
    VN855_data_out <= VN_data_out( 5135 downto 5130 );
    VN855_sign_out <= VN_sign_out( 5135 downto 5130 );
    VN856_data_out <= VN_data_out( 5141 downto 5136 );
    VN856_sign_out <= VN_sign_out( 5141 downto 5136 );
    VN857_data_out <= VN_data_out( 5147 downto 5142 );
    VN857_sign_out <= VN_sign_out( 5147 downto 5142 );
    VN858_data_out <= VN_data_out( 5153 downto 5148 );
    VN858_sign_out <= VN_sign_out( 5153 downto 5148 );
    VN859_data_out <= VN_data_out( 5159 downto 5154 );
    VN859_sign_out <= VN_sign_out( 5159 downto 5154 );
    VN860_data_out <= VN_data_out( 5165 downto 5160 );
    VN860_sign_out <= VN_sign_out( 5165 downto 5160 );
    VN861_data_out <= VN_data_out( 5171 downto 5166 );
    VN861_sign_out <= VN_sign_out( 5171 downto 5166 );
    VN862_data_out <= VN_data_out( 5177 downto 5172 );
    VN862_sign_out <= VN_sign_out( 5177 downto 5172 );
    VN863_data_out <= VN_data_out( 5183 downto 5178 );
    VN863_sign_out <= VN_sign_out( 5183 downto 5178 );
    VN864_data_out <= VN_data_out( 5189 downto 5184 );
    VN864_sign_out <= VN_sign_out( 5189 downto 5184 );
    VN865_data_out <= VN_data_out( 5195 downto 5190 );
    VN865_sign_out <= VN_sign_out( 5195 downto 5190 );
    VN866_data_out <= VN_data_out( 5201 downto 5196 );
    VN866_sign_out <= VN_sign_out( 5201 downto 5196 );
    VN867_data_out <= VN_data_out( 5207 downto 5202 );
    VN867_sign_out <= VN_sign_out( 5207 downto 5202 );
    VN868_data_out <= VN_data_out( 5213 downto 5208 );
    VN868_sign_out <= VN_sign_out( 5213 downto 5208 );
    VN869_data_out <= VN_data_out( 5219 downto 5214 );
    VN869_sign_out <= VN_sign_out( 5219 downto 5214 );
    VN870_data_out <= VN_data_out( 5225 downto 5220 );
    VN870_sign_out <= VN_sign_out( 5225 downto 5220 );
    VN871_data_out <= VN_data_out( 5231 downto 5226 );
    VN871_sign_out <= VN_sign_out( 5231 downto 5226 );
    VN872_data_out <= VN_data_out( 5237 downto 5232 );
    VN872_sign_out <= VN_sign_out( 5237 downto 5232 );
    VN873_data_out <= VN_data_out( 5243 downto 5238 );
    VN873_sign_out <= VN_sign_out( 5243 downto 5238 );
    VN874_data_out <= VN_data_out( 5249 downto 5244 );
    VN874_sign_out <= VN_sign_out( 5249 downto 5244 );
    VN875_data_out <= VN_data_out( 5255 downto 5250 );
    VN875_sign_out <= VN_sign_out( 5255 downto 5250 );
    VN876_data_out <= VN_data_out( 5261 downto 5256 );
    VN876_sign_out <= VN_sign_out( 5261 downto 5256 );
    VN877_data_out <= VN_data_out( 5267 downto 5262 );
    VN877_sign_out <= VN_sign_out( 5267 downto 5262 );
    VN878_data_out <= VN_data_out( 5273 downto 5268 );
    VN878_sign_out <= VN_sign_out( 5273 downto 5268 );
    VN879_data_out <= VN_data_out( 5279 downto 5274 );
    VN879_sign_out <= VN_sign_out( 5279 downto 5274 );
    VN880_data_out <= VN_data_out( 5285 downto 5280 );
    VN880_sign_out <= VN_sign_out( 5285 downto 5280 );
    VN881_data_out <= VN_data_out( 5291 downto 5286 );
    VN881_sign_out <= VN_sign_out( 5291 downto 5286 );
    VN882_data_out <= VN_data_out( 5297 downto 5292 );
    VN882_sign_out <= VN_sign_out( 5297 downto 5292 );
    VN883_data_out <= VN_data_out( 5303 downto 5298 );
    VN883_sign_out <= VN_sign_out( 5303 downto 5298 );
    VN884_data_out <= VN_data_out( 5309 downto 5304 );
    VN884_sign_out <= VN_sign_out( 5309 downto 5304 );
    VN885_data_out <= VN_data_out( 5315 downto 5310 );
    VN885_sign_out <= VN_sign_out( 5315 downto 5310 );
    VN886_data_out <= VN_data_out( 5321 downto 5316 );
    VN886_sign_out <= VN_sign_out( 5321 downto 5316 );
    VN887_data_out <= VN_data_out( 5327 downto 5322 );
    VN887_sign_out <= VN_sign_out( 5327 downto 5322 );
    VN888_data_out <= VN_data_out( 5333 downto 5328 );
    VN888_sign_out <= VN_sign_out( 5333 downto 5328 );
    VN889_data_out <= VN_data_out( 5339 downto 5334 );
    VN889_sign_out <= VN_sign_out( 5339 downto 5334 );
    VN890_data_out <= VN_data_out( 5345 downto 5340 );
    VN890_sign_out <= VN_sign_out( 5345 downto 5340 );
    VN891_data_out <= VN_data_out( 5351 downto 5346 );
    VN891_sign_out <= VN_sign_out( 5351 downto 5346 );
    VN892_data_out <= VN_data_out( 5357 downto 5352 );
    VN892_sign_out <= VN_sign_out( 5357 downto 5352 );
    VN893_data_out <= VN_data_out( 5363 downto 5358 );
    VN893_sign_out <= VN_sign_out( 5363 downto 5358 );
    VN894_data_out <= VN_data_out( 5369 downto 5364 );
    VN894_sign_out <= VN_sign_out( 5369 downto 5364 );
    VN895_data_out <= VN_data_out( 5375 downto 5370 );
    VN895_sign_out <= VN_sign_out( 5375 downto 5370 );
    VN896_data_out <= VN_data_out( 5381 downto 5376 );
    VN896_sign_out <= VN_sign_out( 5381 downto 5376 );
    VN897_data_out <= VN_data_out( 5387 downto 5382 );
    VN897_sign_out <= VN_sign_out( 5387 downto 5382 );
    VN898_data_out <= VN_data_out( 5393 downto 5388 );
    VN898_sign_out <= VN_sign_out( 5393 downto 5388 );
    VN899_data_out <= VN_data_out( 5399 downto 5394 );
    VN899_sign_out <= VN_sign_out( 5399 downto 5394 );
    VN900_data_out <= VN_data_out( 5405 downto 5400 );
    VN900_sign_out <= VN_sign_out( 5405 downto 5400 );
    VN901_data_out <= VN_data_out( 5411 downto 5406 );
    VN901_sign_out <= VN_sign_out( 5411 downto 5406 );
    VN902_data_out <= VN_data_out( 5417 downto 5412 );
    VN902_sign_out <= VN_sign_out( 5417 downto 5412 );
    VN903_data_out <= VN_data_out( 5423 downto 5418 );
    VN903_sign_out <= VN_sign_out( 5423 downto 5418 );
    VN904_data_out <= VN_data_out( 5429 downto 5424 );
    VN904_sign_out <= VN_sign_out( 5429 downto 5424 );
    VN905_data_out <= VN_data_out( 5435 downto 5430 );
    VN905_sign_out <= VN_sign_out( 5435 downto 5430 );
    VN906_data_out <= VN_data_out( 5441 downto 5436 );
    VN906_sign_out <= VN_sign_out( 5441 downto 5436 );
    VN907_data_out <= VN_data_out( 5447 downto 5442 );
    VN907_sign_out <= VN_sign_out( 5447 downto 5442 );
    VN908_data_out <= VN_data_out( 5453 downto 5448 );
    VN908_sign_out <= VN_sign_out( 5453 downto 5448 );
    VN909_data_out <= VN_data_out( 5459 downto 5454 );
    VN909_sign_out <= VN_sign_out( 5459 downto 5454 );
    VN910_data_out <= VN_data_out( 5465 downto 5460 );
    VN910_sign_out <= VN_sign_out( 5465 downto 5460 );
    VN911_data_out <= VN_data_out( 5471 downto 5466 );
    VN911_sign_out <= VN_sign_out( 5471 downto 5466 );
    VN912_data_out <= VN_data_out( 5477 downto 5472 );
    VN912_sign_out <= VN_sign_out( 5477 downto 5472 );
    VN913_data_out <= VN_data_out( 5483 downto 5478 );
    VN913_sign_out <= VN_sign_out( 5483 downto 5478 );
    VN914_data_out <= VN_data_out( 5489 downto 5484 );
    VN914_sign_out <= VN_sign_out( 5489 downto 5484 );
    VN915_data_out <= VN_data_out( 5495 downto 5490 );
    VN915_sign_out <= VN_sign_out( 5495 downto 5490 );
    VN916_data_out <= VN_data_out( 5501 downto 5496 );
    VN916_sign_out <= VN_sign_out( 5501 downto 5496 );
    VN917_data_out <= VN_data_out( 5507 downto 5502 );
    VN917_sign_out <= VN_sign_out( 5507 downto 5502 );
    VN918_data_out <= VN_data_out( 5513 downto 5508 );
    VN918_sign_out <= VN_sign_out( 5513 downto 5508 );
    VN919_data_out <= VN_data_out( 5519 downto 5514 );
    VN919_sign_out <= VN_sign_out( 5519 downto 5514 );
    VN920_data_out <= VN_data_out( 5525 downto 5520 );
    VN920_sign_out <= VN_sign_out( 5525 downto 5520 );
    VN921_data_out <= VN_data_out( 5531 downto 5526 );
    VN921_sign_out <= VN_sign_out( 5531 downto 5526 );
    VN922_data_out <= VN_data_out( 5537 downto 5532 );
    VN922_sign_out <= VN_sign_out( 5537 downto 5532 );
    VN923_data_out <= VN_data_out( 5543 downto 5538 );
    VN923_sign_out <= VN_sign_out( 5543 downto 5538 );
    VN924_data_out <= VN_data_out( 5549 downto 5544 );
    VN924_sign_out <= VN_sign_out( 5549 downto 5544 );
    VN925_data_out <= VN_data_out( 5555 downto 5550 );
    VN925_sign_out <= VN_sign_out( 5555 downto 5550 );
    VN926_data_out <= VN_data_out( 5561 downto 5556 );
    VN926_sign_out <= VN_sign_out( 5561 downto 5556 );
    VN927_data_out <= VN_data_out( 5567 downto 5562 );
    VN927_sign_out <= VN_sign_out( 5567 downto 5562 );
    VN928_data_out <= VN_data_out( 5573 downto 5568 );
    VN928_sign_out <= VN_sign_out( 5573 downto 5568 );
    VN929_data_out <= VN_data_out( 5579 downto 5574 );
    VN929_sign_out <= VN_sign_out( 5579 downto 5574 );
    VN930_data_out <= VN_data_out( 5585 downto 5580 );
    VN930_sign_out <= VN_sign_out( 5585 downto 5580 );
    VN931_data_out <= VN_data_out( 5591 downto 5586 );
    VN931_sign_out <= VN_sign_out( 5591 downto 5586 );
    VN932_data_out <= VN_data_out( 5597 downto 5592 );
    VN932_sign_out <= VN_sign_out( 5597 downto 5592 );
    VN933_data_out <= VN_data_out( 5603 downto 5598 );
    VN933_sign_out <= VN_sign_out( 5603 downto 5598 );
    VN934_data_out <= VN_data_out( 5609 downto 5604 );
    VN934_sign_out <= VN_sign_out( 5609 downto 5604 );
    VN935_data_out <= VN_data_out( 5615 downto 5610 );
    VN935_sign_out <= VN_sign_out( 5615 downto 5610 );
    VN936_data_out <= VN_data_out( 5621 downto 5616 );
    VN936_sign_out <= VN_sign_out( 5621 downto 5616 );
    VN937_data_out <= VN_data_out( 5627 downto 5622 );
    VN937_sign_out <= VN_sign_out( 5627 downto 5622 );
    VN938_data_out <= VN_data_out( 5633 downto 5628 );
    VN938_sign_out <= VN_sign_out( 5633 downto 5628 );
    VN939_data_out <= VN_data_out( 5639 downto 5634 );
    VN939_sign_out <= VN_sign_out( 5639 downto 5634 );
    VN940_data_out <= VN_data_out( 5645 downto 5640 );
    VN940_sign_out <= VN_sign_out( 5645 downto 5640 );
    VN941_data_out <= VN_data_out( 5651 downto 5646 );
    VN941_sign_out <= VN_sign_out( 5651 downto 5646 );
    VN942_data_out <= VN_data_out( 5657 downto 5652 );
    VN942_sign_out <= VN_sign_out( 5657 downto 5652 );
    VN943_data_out <= VN_data_out( 5663 downto 5658 );
    VN943_sign_out <= VN_sign_out( 5663 downto 5658 );
    VN944_data_out <= VN_data_out( 5669 downto 5664 );
    VN944_sign_out <= VN_sign_out( 5669 downto 5664 );
    VN945_data_out <= VN_data_out( 5675 downto 5670 );
    VN945_sign_out <= VN_sign_out( 5675 downto 5670 );
    VN946_data_out <= VN_data_out( 5681 downto 5676 );
    VN946_sign_out <= VN_sign_out( 5681 downto 5676 );
    VN947_data_out <= VN_data_out( 5687 downto 5682 );
    VN947_sign_out <= VN_sign_out( 5687 downto 5682 );
    VN948_data_out <= VN_data_out( 5693 downto 5688 );
    VN948_sign_out <= VN_sign_out( 5693 downto 5688 );
    VN949_data_out <= VN_data_out( 5699 downto 5694 );
    VN949_sign_out <= VN_sign_out( 5699 downto 5694 );
    VN950_data_out <= VN_data_out( 5705 downto 5700 );
    VN950_sign_out <= VN_sign_out( 5705 downto 5700 );
    VN951_data_out <= VN_data_out( 5711 downto 5706 );
    VN951_sign_out <= VN_sign_out( 5711 downto 5706 );
    VN952_data_out <= VN_data_out( 5717 downto 5712 );
    VN952_sign_out <= VN_sign_out( 5717 downto 5712 );
    VN953_data_out <= VN_data_out( 5723 downto 5718 );
    VN953_sign_out <= VN_sign_out( 5723 downto 5718 );
    VN954_data_out <= VN_data_out( 5729 downto 5724 );
    VN954_sign_out <= VN_sign_out( 5729 downto 5724 );
    VN955_data_out <= VN_data_out( 5735 downto 5730 );
    VN955_sign_out <= VN_sign_out( 5735 downto 5730 );
    VN956_data_out <= VN_data_out( 5741 downto 5736 );
    VN956_sign_out <= VN_sign_out( 5741 downto 5736 );
    VN957_data_out <= VN_data_out( 5747 downto 5742 );
    VN957_sign_out <= VN_sign_out( 5747 downto 5742 );
    VN958_data_out <= VN_data_out( 5753 downto 5748 );
    VN958_sign_out <= VN_sign_out( 5753 downto 5748 );
    VN959_data_out <= VN_data_out( 5759 downto 5754 );
    VN959_sign_out <= VN_sign_out( 5759 downto 5754 );
    VN960_data_out <= VN_data_out( 5765 downto 5760 );
    VN960_sign_out <= VN_sign_out( 5765 downto 5760 );
    VN961_data_out <= VN_data_out( 5771 downto 5766 );
    VN961_sign_out <= VN_sign_out( 5771 downto 5766 );
    VN962_data_out <= VN_data_out( 5777 downto 5772 );
    VN962_sign_out <= VN_sign_out( 5777 downto 5772 );
    VN963_data_out <= VN_data_out( 5783 downto 5778 );
    VN963_sign_out <= VN_sign_out( 5783 downto 5778 );
    VN964_data_out <= VN_data_out( 5789 downto 5784 );
    VN964_sign_out <= VN_sign_out( 5789 downto 5784 );
    VN965_data_out <= VN_data_out( 5795 downto 5790 );
    VN965_sign_out <= VN_sign_out( 5795 downto 5790 );
    VN966_data_out <= VN_data_out( 5801 downto 5796 );
    VN966_sign_out <= VN_sign_out( 5801 downto 5796 );
    VN967_data_out <= VN_data_out( 5807 downto 5802 );
    VN967_sign_out <= VN_sign_out( 5807 downto 5802 );
    VN968_data_out <= VN_data_out( 5813 downto 5808 );
    VN968_sign_out <= VN_sign_out( 5813 downto 5808 );
    VN969_data_out <= VN_data_out( 5819 downto 5814 );
    VN969_sign_out <= VN_sign_out( 5819 downto 5814 );
    VN970_data_out <= VN_data_out( 5825 downto 5820 );
    VN970_sign_out <= VN_sign_out( 5825 downto 5820 );
    VN971_data_out <= VN_data_out( 5831 downto 5826 );
    VN971_sign_out <= VN_sign_out( 5831 downto 5826 );
    VN972_data_out <= VN_data_out( 5837 downto 5832 );
    VN972_sign_out <= VN_sign_out( 5837 downto 5832 );
    VN973_data_out <= VN_data_out( 5843 downto 5838 );
    VN973_sign_out <= VN_sign_out( 5843 downto 5838 );
    VN974_data_out <= VN_data_out( 5849 downto 5844 );
    VN974_sign_out <= VN_sign_out( 5849 downto 5844 );
    VN975_data_out <= VN_data_out( 5855 downto 5850 );
    VN975_sign_out <= VN_sign_out( 5855 downto 5850 );
    VN976_data_out <= VN_data_out( 5861 downto 5856 );
    VN976_sign_out <= VN_sign_out( 5861 downto 5856 );
    VN977_data_out <= VN_data_out( 5867 downto 5862 );
    VN977_sign_out <= VN_sign_out( 5867 downto 5862 );
    VN978_data_out <= VN_data_out( 5873 downto 5868 );
    VN978_sign_out <= VN_sign_out( 5873 downto 5868 );
    VN979_data_out <= VN_data_out( 5879 downto 5874 );
    VN979_sign_out <= VN_sign_out( 5879 downto 5874 );
    VN980_data_out <= VN_data_out( 5885 downto 5880 );
    VN980_sign_out <= VN_sign_out( 5885 downto 5880 );
    VN981_data_out <= VN_data_out( 5891 downto 5886 );
    VN981_sign_out <= VN_sign_out( 5891 downto 5886 );
    VN982_data_out <= VN_data_out( 5897 downto 5892 );
    VN982_sign_out <= VN_sign_out( 5897 downto 5892 );
    VN983_data_out <= VN_data_out( 5903 downto 5898 );
    VN983_sign_out <= VN_sign_out( 5903 downto 5898 );
    VN984_data_out <= VN_data_out( 5909 downto 5904 );
    VN984_sign_out <= VN_sign_out( 5909 downto 5904 );
    VN985_data_out <= VN_data_out( 5915 downto 5910 );
    VN985_sign_out <= VN_sign_out( 5915 downto 5910 );
    VN986_data_out <= VN_data_out( 5921 downto 5916 );
    VN986_sign_out <= VN_sign_out( 5921 downto 5916 );
    VN987_data_out <= VN_data_out( 5927 downto 5922 );
    VN987_sign_out <= VN_sign_out( 5927 downto 5922 );
    VN988_data_out <= VN_data_out( 5933 downto 5928 );
    VN988_sign_out <= VN_sign_out( 5933 downto 5928 );
    VN989_data_out <= VN_data_out( 5939 downto 5934 );
    VN989_sign_out <= VN_sign_out( 5939 downto 5934 );
    VN990_data_out <= VN_data_out( 5945 downto 5940 );
    VN990_sign_out <= VN_sign_out( 5945 downto 5940 );
    VN991_data_out <= VN_data_out( 5951 downto 5946 );
    VN991_sign_out <= VN_sign_out( 5951 downto 5946 );
    VN992_data_out <= VN_data_out( 5957 downto 5952 );
    VN992_sign_out <= VN_sign_out( 5957 downto 5952 );
    VN993_data_out <= VN_data_out( 5963 downto 5958 );
    VN993_sign_out <= VN_sign_out( 5963 downto 5958 );
    VN994_data_out <= VN_data_out( 5969 downto 5964 );
    VN994_sign_out <= VN_sign_out( 5969 downto 5964 );
    VN995_data_out <= VN_data_out( 5975 downto 5970 );
    VN995_sign_out <= VN_sign_out( 5975 downto 5970 );
    VN996_data_out <= VN_data_out( 5981 downto 5976 );
    VN996_sign_out <= VN_sign_out( 5981 downto 5976 );
    VN997_data_out <= VN_data_out( 5987 downto 5982 );
    VN997_sign_out <= VN_sign_out( 5987 downto 5982 );
    VN998_data_out <= VN_data_out( 5993 downto 5988 );
    VN998_sign_out <= VN_sign_out( 5993 downto 5988 );
    VN999_data_out <= VN_data_out( 5999 downto 5994 );
    VN999_sign_out <= VN_sign_out( 5999 downto 5994 );
    VN1000_data_out <= VN_data_out( 6005 downto 6000 );
    VN1000_sign_out <= VN_sign_out( 6005 downto 6000 );
    VN1001_data_out <= VN_data_out( 6011 downto 6006 );
    VN1001_sign_out <= VN_sign_out( 6011 downto 6006 );
    VN1002_data_out <= VN_data_out( 6017 downto 6012 );
    VN1002_sign_out <= VN_sign_out( 6017 downto 6012 );
    VN1003_data_out <= VN_data_out( 6023 downto 6018 );
    VN1003_sign_out <= VN_sign_out( 6023 downto 6018 );
    VN1004_data_out <= VN_data_out( 6029 downto 6024 );
    VN1004_sign_out <= VN_sign_out( 6029 downto 6024 );
    VN1005_data_out <= VN_data_out( 6035 downto 6030 );
    VN1005_sign_out <= VN_sign_out( 6035 downto 6030 );
    VN1006_data_out <= VN_data_out( 6041 downto 6036 );
    VN1006_sign_out <= VN_sign_out( 6041 downto 6036 );
    VN1007_data_out <= VN_data_out( 6047 downto 6042 );
    VN1007_sign_out <= VN_sign_out( 6047 downto 6042 );
    VN1008_data_out <= VN_data_out( 6053 downto 6048 );
    VN1008_sign_out <= VN_sign_out( 6053 downto 6048 );
    VN1009_data_out <= VN_data_out( 6059 downto 6054 );
    VN1009_sign_out <= VN_sign_out( 6059 downto 6054 );
    VN1010_data_out <= VN_data_out( 6065 downto 6060 );
    VN1010_sign_out <= VN_sign_out( 6065 downto 6060 );
    VN1011_data_out <= VN_data_out( 6071 downto 6066 );
    VN1011_sign_out <= VN_sign_out( 6071 downto 6066 );
    VN1012_data_out <= VN_data_out( 6077 downto 6072 );
    VN1012_sign_out <= VN_sign_out( 6077 downto 6072 );
    VN1013_data_out <= VN_data_out( 6083 downto 6078 );
    VN1013_sign_out <= VN_sign_out( 6083 downto 6078 );
    VN1014_data_out <= VN_data_out( 6089 downto 6084 );
    VN1014_sign_out <= VN_sign_out( 6089 downto 6084 );
    VN1015_data_out <= VN_data_out( 6095 downto 6090 );
    VN1015_sign_out <= VN_sign_out( 6095 downto 6090 );
    VN1016_data_out <= VN_data_out( 6101 downto 6096 );
    VN1016_sign_out <= VN_sign_out( 6101 downto 6096 );
    VN1017_data_out <= VN_data_out( 6107 downto 6102 );
    VN1017_sign_out <= VN_sign_out( 6107 downto 6102 );
    VN1018_data_out <= VN_data_out( 6113 downto 6108 );
    VN1018_sign_out <= VN_sign_out( 6113 downto 6108 );
    VN1019_data_out <= VN_data_out( 6119 downto 6114 );
    VN1019_sign_out <= VN_sign_out( 6119 downto 6114 );
    VN1020_data_out <= VN_data_out( 6125 downto 6120 );
    VN1020_sign_out <= VN_sign_out( 6125 downto 6120 );
    VN1021_data_out <= VN_data_out( 6131 downto 6126 );
    VN1021_sign_out <= VN_sign_out( 6131 downto 6126 );
    VN1022_data_out <= VN_data_out( 6137 downto 6132 );
    VN1022_sign_out <= VN_sign_out( 6137 downto 6132 );
    VN1023_data_out <= VN_data_out( 6143 downto 6138 );
    VN1023_sign_out <= VN_sign_out( 6143 downto 6138 );
    VN1024_data_out <= VN_data_out( 6149 downto 6144 );
    VN1024_sign_out <= VN_sign_out( 6149 downto 6144 );
    VN1025_data_out <= VN_data_out( 6155 downto 6150 );
    VN1025_sign_out <= VN_sign_out( 6155 downto 6150 );
    VN1026_data_out <= VN_data_out( 6161 downto 6156 );
    VN1026_sign_out <= VN_sign_out( 6161 downto 6156 );
    VN1027_data_out <= VN_data_out( 6167 downto 6162 );
    VN1027_sign_out <= VN_sign_out( 6167 downto 6162 );
    VN1028_data_out <= VN_data_out( 6173 downto 6168 );
    VN1028_sign_out <= VN_sign_out( 6173 downto 6168 );
    VN1029_data_out <= VN_data_out( 6179 downto 6174 );
    VN1029_sign_out <= VN_sign_out( 6179 downto 6174 );
    VN1030_data_out <= VN_data_out( 6185 downto 6180 );
    VN1030_sign_out <= VN_sign_out( 6185 downto 6180 );
    VN1031_data_out <= VN_data_out( 6191 downto 6186 );
    VN1031_sign_out <= VN_sign_out( 6191 downto 6186 );
    VN1032_data_out <= VN_data_out( 6197 downto 6192 );
    VN1032_sign_out <= VN_sign_out( 6197 downto 6192 );
    VN1033_data_out <= VN_data_out( 6203 downto 6198 );
    VN1033_sign_out <= VN_sign_out( 6203 downto 6198 );
    VN1034_data_out <= VN_data_out( 6209 downto 6204 );
    VN1034_sign_out <= VN_sign_out( 6209 downto 6204 );
    VN1035_data_out <= VN_data_out( 6215 downto 6210 );
    VN1035_sign_out <= VN_sign_out( 6215 downto 6210 );
    VN1036_data_out <= VN_data_out( 6221 downto 6216 );
    VN1036_sign_out <= VN_sign_out( 6221 downto 6216 );
    VN1037_data_out <= VN_data_out( 6227 downto 6222 );
    VN1037_sign_out <= VN_sign_out( 6227 downto 6222 );
    VN1038_data_out <= VN_data_out( 6233 downto 6228 );
    VN1038_sign_out <= VN_sign_out( 6233 downto 6228 );
    VN1039_data_out <= VN_data_out( 6239 downto 6234 );
    VN1039_sign_out <= VN_sign_out( 6239 downto 6234 );
    VN1040_data_out <= VN_data_out( 6245 downto 6240 );
    VN1040_sign_out <= VN_sign_out( 6245 downto 6240 );
    VN1041_data_out <= VN_data_out( 6251 downto 6246 );
    VN1041_sign_out <= VN_sign_out( 6251 downto 6246 );
    VN1042_data_out <= VN_data_out( 6257 downto 6252 );
    VN1042_sign_out <= VN_sign_out( 6257 downto 6252 );
    VN1043_data_out <= VN_data_out( 6263 downto 6258 );
    VN1043_sign_out <= VN_sign_out( 6263 downto 6258 );
    VN1044_data_out <= VN_data_out( 6269 downto 6264 );
    VN1044_sign_out <= VN_sign_out( 6269 downto 6264 );
    VN1045_data_out <= VN_data_out( 6275 downto 6270 );
    VN1045_sign_out <= VN_sign_out( 6275 downto 6270 );
    VN1046_data_out <= VN_data_out( 6281 downto 6276 );
    VN1046_sign_out <= VN_sign_out( 6281 downto 6276 );
    VN1047_data_out <= VN_data_out( 6287 downto 6282 );
    VN1047_sign_out <= VN_sign_out( 6287 downto 6282 );
    VN1048_data_out <= VN_data_out( 6293 downto 6288 );
    VN1048_sign_out <= VN_sign_out( 6293 downto 6288 );
    VN1049_data_out <= VN_data_out( 6299 downto 6294 );
    VN1049_sign_out <= VN_sign_out( 6299 downto 6294 );
    VN1050_data_out <= VN_data_out( 6305 downto 6300 );
    VN1050_sign_out <= VN_sign_out( 6305 downto 6300 );
    VN1051_data_out <= VN_data_out( 6311 downto 6306 );
    VN1051_sign_out <= VN_sign_out( 6311 downto 6306 );
    VN1052_data_out <= VN_data_out( 6317 downto 6312 );
    VN1052_sign_out <= VN_sign_out( 6317 downto 6312 );
    VN1053_data_out <= VN_data_out( 6323 downto 6318 );
    VN1053_sign_out <= VN_sign_out( 6323 downto 6318 );
    VN1054_data_out <= VN_data_out( 6329 downto 6324 );
    VN1054_sign_out <= VN_sign_out( 6329 downto 6324 );
    VN1055_data_out <= VN_data_out( 6335 downto 6330 );
    VN1055_sign_out <= VN_sign_out( 6335 downto 6330 );
    VN1056_data_out <= VN_data_out( 6341 downto 6336 );
    VN1056_sign_out <= VN_sign_out( 6341 downto 6336 );
    VN1057_data_out <= VN_data_out( 6347 downto 6342 );
    VN1057_sign_out <= VN_sign_out( 6347 downto 6342 );
    VN1058_data_out <= VN_data_out( 6353 downto 6348 );
    VN1058_sign_out <= VN_sign_out( 6353 downto 6348 );
    VN1059_data_out <= VN_data_out( 6359 downto 6354 );
    VN1059_sign_out <= VN_sign_out( 6359 downto 6354 );
    VN1060_data_out <= VN_data_out( 6365 downto 6360 );
    VN1060_sign_out <= VN_sign_out( 6365 downto 6360 );
    VN1061_data_out <= VN_data_out( 6371 downto 6366 );
    VN1061_sign_out <= VN_sign_out( 6371 downto 6366 );
    VN1062_data_out <= VN_data_out( 6377 downto 6372 );
    VN1062_sign_out <= VN_sign_out( 6377 downto 6372 );
    VN1063_data_out <= VN_data_out( 6383 downto 6378 );
    VN1063_sign_out <= VN_sign_out( 6383 downto 6378 );
    VN1064_data_out <= VN_data_out( 6389 downto 6384 );
    VN1064_sign_out <= VN_sign_out( 6389 downto 6384 );
    VN1065_data_out <= VN_data_out( 6395 downto 6390 );
    VN1065_sign_out <= VN_sign_out( 6395 downto 6390 );
    VN1066_data_out <= VN_data_out( 6401 downto 6396 );
    VN1066_sign_out <= VN_sign_out( 6401 downto 6396 );
    VN1067_data_out <= VN_data_out( 6407 downto 6402 );
    VN1067_sign_out <= VN_sign_out( 6407 downto 6402 );
    VN1068_data_out <= VN_data_out( 6413 downto 6408 );
    VN1068_sign_out <= VN_sign_out( 6413 downto 6408 );
    VN1069_data_out <= VN_data_out( 6419 downto 6414 );
    VN1069_sign_out <= VN_sign_out( 6419 downto 6414 );
    VN1070_data_out <= VN_data_out( 6425 downto 6420 );
    VN1070_sign_out <= VN_sign_out( 6425 downto 6420 );
    VN1071_data_out <= VN_data_out( 6431 downto 6426 );
    VN1071_sign_out <= VN_sign_out( 6431 downto 6426 );
    VN1072_data_out <= VN_data_out( 6437 downto 6432 );
    VN1072_sign_out <= VN_sign_out( 6437 downto 6432 );
    VN1073_data_out <= VN_data_out( 6443 downto 6438 );
    VN1073_sign_out <= VN_sign_out( 6443 downto 6438 );
    VN1074_data_out <= VN_data_out( 6449 downto 6444 );
    VN1074_sign_out <= VN_sign_out( 6449 downto 6444 );
    VN1075_data_out <= VN_data_out( 6455 downto 6450 );
    VN1075_sign_out <= VN_sign_out( 6455 downto 6450 );
    VN1076_data_out <= VN_data_out( 6461 downto 6456 );
    VN1076_sign_out <= VN_sign_out( 6461 downto 6456 );
    VN1077_data_out <= VN_data_out( 6467 downto 6462 );
    VN1077_sign_out <= VN_sign_out( 6467 downto 6462 );
    VN1078_data_out <= VN_data_out( 6473 downto 6468 );
    VN1078_sign_out <= VN_sign_out( 6473 downto 6468 );
    VN1079_data_out <= VN_data_out( 6479 downto 6474 );
    VN1079_sign_out <= VN_sign_out( 6479 downto 6474 );
    VN1080_data_out <= VN_data_out( 6485 downto 6480 );
    VN1080_sign_out <= VN_sign_out( 6485 downto 6480 );
    VN1081_data_out <= VN_data_out( 6491 downto 6486 );
    VN1081_sign_out <= VN_sign_out( 6491 downto 6486 );
    VN1082_data_out <= VN_data_out( 6497 downto 6492 );
    VN1082_sign_out <= VN_sign_out( 6497 downto 6492 );
    VN1083_data_out <= VN_data_out( 6503 downto 6498 );
    VN1083_sign_out <= VN_sign_out( 6503 downto 6498 );
    VN1084_data_out <= VN_data_out( 6509 downto 6504 );
    VN1084_sign_out <= VN_sign_out( 6509 downto 6504 );
    VN1085_data_out <= VN_data_out( 6515 downto 6510 );
    VN1085_sign_out <= VN_sign_out( 6515 downto 6510 );
    VN1086_data_out <= VN_data_out( 6521 downto 6516 );
    VN1086_sign_out <= VN_sign_out( 6521 downto 6516 );
    VN1087_data_out <= VN_data_out( 6527 downto 6522 );
    VN1087_sign_out <= VN_sign_out( 6527 downto 6522 );
    VN1088_data_out <= VN_data_out( 6533 downto 6528 );
    VN1088_sign_out <= VN_sign_out( 6533 downto 6528 );
    VN1089_data_out <= VN_data_out( 6539 downto 6534 );
    VN1089_sign_out <= VN_sign_out( 6539 downto 6534 );
    VN1090_data_out <= VN_data_out( 6545 downto 6540 );
    VN1090_sign_out <= VN_sign_out( 6545 downto 6540 );
    VN1091_data_out <= VN_data_out( 6551 downto 6546 );
    VN1091_sign_out <= VN_sign_out( 6551 downto 6546 );
    VN1092_data_out <= VN_data_out( 6557 downto 6552 );
    VN1092_sign_out <= VN_sign_out( 6557 downto 6552 );
    VN1093_data_out <= VN_data_out( 6563 downto 6558 );
    VN1093_sign_out <= VN_sign_out( 6563 downto 6558 );
    VN1094_data_out <= VN_data_out( 6569 downto 6564 );
    VN1094_sign_out <= VN_sign_out( 6569 downto 6564 );
    VN1095_data_out <= VN_data_out( 6575 downto 6570 );
    VN1095_sign_out <= VN_sign_out( 6575 downto 6570 );
    VN1096_data_out <= VN_data_out( 6581 downto 6576 );
    VN1096_sign_out <= VN_sign_out( 6581 downto 6576 );
    VN1097_data_out <= VN_data_out( 6587 downto 6582 );
    VN1097_sign_out <= VN_sign_out( 6587 downto 6582 );
    VN1098_data_out <= VN_data_out( 6593 downto 6588 );
    VN1098_sign_out <= VN_sign_out( 6593 downto 6588 );
    VN1099_data_out <= VN_data_out( 6599 downto 6594 );
    VN1099_sign_out <= VN_sign_out( 6599 downto 6594 );
    VN1100_data_out <= VN_data_out( 6605 downto 6600 );
    VN1100_sign_out <= VN_sign_out( 6605 downto 6600 );
    VN1101_data_out <= VN_data_out( 6611 downto 6606 );
    VN1101_sign_out <= VN_sign_out( 6611 downto 6606 );
    VN1102_data_out <= VN_data_out( 6617 downto 6612 );
    VN1102_sign_out <= VN_sign_out( 6617 downto 6612 );
    VN1103_data_out <= VN_data_out( 6623 downto 6618 );
    VN1103_sign_out <= VN_sign_out( 6623 downto 6618 );
    VN1104_data_out <= VN_data_out( 6629 downto 6624 );
    VN1104_sign_out <= VN_sign_out( 6629 downto 6624 );
    VN1105_data_out <= VN_data_out( 6635 downto 6630 );
    VN1105_sign_out <= VN_sign_out( 6635 downto 6630 );
    VN1106_data_out <= VN_data_out( 6641 downto 6636 );
    VN1106_sign_out <= VN_sign_out( 6641 downto 6636 );
    VN1107_data_out <= VN_data_out( 6647 downto 6642 );
    VN1107_sign_out <= VN_sign_out( 6647 downto 6642 );
    VN1108_data_out <= VN_data_out( 6653 downto 6648 );
    VN1108_sign_out <= VN_sign_out( 6653 downto 6648 );
    VN1109_data_out <= VN_data_out( 6659 downto 6654 );
    VN1109_sign_out <= VN_sign_out( 6659 downto 6654 );
    VN1110_data_out <= VN_data_out( 6665 downto 6660 );
    VN1110_sign_out <= VN_sign_out( 6665 downto 6660 );
    VN1111_data_out <= VN_data_out( 6671 downto 6666 );
    VN1111_sign_out <= VN_sign_out( 6671 downto 6666 );
    VN1112_data_out <= VN_data_out( 6677 downto 6672 );
    VN1112_sign_out <= VN_sign_out( 6677 downto 6672 );
    VN1113_data_out <= VN_data_out( 6683 downto 6678 );
    VN1113_sign_out <= VN_sign_out( 6683 downto 6678 );
    VN1114_data_out <= VN_data_out( 6689 downto 6684 );
    VN1114_sign_out <= VN_sign_out( 6689 downto 6684 );
    VN1115_data_out <= VN_data_out( 6695 downto 6690 );
    VN1115_sign_out <= VN_sign_out( 6695 downto 6690 );
    VN1116_data_out <= VN_data_out( 6701 downto 6696 );
    VN1116_sign_out <= VN_sign_out( 6701 downto 6696 );
    VN1117_data_out <= VN_data_out( 6707 downto 6702 );
    VN1117_sign_out <= VN_sign_out( 6707 downto 6702 );
    VN1118_data_out <= VN_data_out( 6713 downto 6708 );
    VN1118_sign_out <= VN_sign_out( 6713 downto 6708 );
    VN1119_data_out <= VN_data_out( 6719 downto 6714 );
    VN1119_sign_out <= VN_sign_out( 6719 downto 6714 );
    VN1120_data_out <= VN_data_out( 6725 downto 6720 );
    VN1120_sign_out <= VN_sign_out( 6725 downto 6720 );
    VN1121_data_out <= VN_data_out( 6731 downto 6726 );
    VN1121_sign_out <= VN_sign_out( 6731 downto 6726 );
    VN1122_data_out <= VN_data_out( 6737 downto 6732 );
    VN1122_sign_out <= VN_sign_out( 6737 downto 6732 );
    VN1123_data_out <= VN_data_out( 6743 downto 6738 );
    VN1123_sign_out <= VN_sign_out( 6743 downto 6738 );
    VN1124_data_out <= VN_data_out( 6749 downto 6744 );
    VN1124_sign_out <= VN_sign_out( 6749 downto 6744 );
    VN1125_data_out <= VN_data_out( 6755 downto 6750 );
    VN1125_sign_out <= VN_sign_out( 6755 downto 6750 );
    VN1126_data_out <= VN_data_out( 6761 downto 6756 );
    VN1126_sign_out <= VN_sign_out( 6761 downto 6756 );
    VN1127_data_out <= VN_data_out( 6767 downto 6762 );
    VN1127_sign_out <= VN_sign_out( 6767 downto 6762 );
    VN1128_data_out <= VN_data_out( 6773 downto 6768 );
    VN1128_sign_out <= VN_sign_out( 6773 downto 6768 );
    VN1129_data_out <= VN_data_out( 6779 downto 6774 );
    VN1129_sign_out <= VN_sign_out( 6779 downto 6774 );
    VN1130_data_out <= VN_data_out( 6785 downto 6780 );
    VN1130_sign_out <= VN_sign_out( 6785 downto 6780 );
    VN1131_data_out <= VN_data_out( 6791 downto 6786 );
    VN1131_sign_out <= VN_sign_out( 6791 downto 6786 );
    VN1132_data_out <= VN_data_out( 6797 downto 6792 );
    VN1132_sign_out <= VN_sign_out( 6797 downto 6792 );
    VN1133_data_out <= VN_data_out( 6803 downto 6798 );
    VN1133_sign_out <= VN_sign_out( 6803 downto 6798 );
    VN1134_data_out <= VN_data_out( 6809 downto 6804 );
    VN1134_sign_out <= VN_sign_out( 6809 downto 6804 );
    VN1135_data_out <= VN_data_out( 6815 downto 6810 );
    VN1135_sign_out <= VN_sign_out( 6815 downto 6810 );
    VN1136_data_out <= VN_data_out( 6821 downto 6816 );
    VN1136_sign_out <= VN_sign_out( 6821 downto 6816 );
    VN1137_data_out <= VN_data_out( 6827 downto 6822 );
    VN1137_sign_out <= VN_sign_out( 6827 downto 6822 );
    VN1138_data_out <= VN_data_out( 6833 downto 6828 );
    VN1138_sign_out <= VN_sign_out( 6833 downto 6828 );
    VN1139_data_out <= VN_data_out( 6839 downto 6834 );
    VN1139_sign_out <= VN_sign_out( 6839 downto 6834 );
    VN1140_data_out <= VN_data_out( 6845 downto 6840 );
    VN1140_sign_out <= VN_sign_out( 6845 downto 6840 );
    VN1141_data_out <= VN_data_out( 6851 downto 6846 );
    VN1141_sign_out <= VN_sign_out( 6851 downto 6846 );
    VN1142_data_out <= VN_data_out( 6857 downto 6852 );
    VN1142_sign_out <= VN_sign_out( 6857 downto 6852 );
    VN1143_data_out <= VN_data_out( 6863 downto 6858 );
    VN1143_sign_out <= VN_sign_out( 6863 downto 6858 );
    VN1144_data_out <= VN_data_out( 6869 downto 6864 );
    VN1144_sign_out <= VN_sign_out( 6869 downto 6864 );
    VN1145_data_out <= VN_data_out( 6875 downto 6870 );
    VN1145_sign_out <= VN_sign_out( 6875 downto 6870 );
    VN1146_data_out <= VN_data_out( 6881 downto 6876 );
    VN1146_sign_out <= VN_sign_out( 6881 downto 6876 );
    VN1147_data_out <= VN_data_out( 6887 downto 6882 );
    VN1147_sign_out <= VN_sign_out( 6887 downto 6882 );
    VN1148_data_out <= VN_data_out( 6893 downto 6888 );
    VN1148_sign_out <= VN_sign_out( 6893 downto 6888 );
    VN1149_data_out <= VN_data_out( 6899 downto 6894 );
    VN1149_sign_out <= VN_sign_out( 6899 downto 6894 );
    VN1150_data_out <= VN_data_out( 6905 downto 6900 );
    VN1150_sign_out <= VN_sign_out( 6905 downto 6900 );
    VN1151_data_out <= VN_data_out( 6911 downto 6906 );
    VN1151_sign_out <= VN_sign_out( 6911 downto 6906 );
    VN1152_data_out <= VN_data_out( 6917 downto 6912 );
    VN1152_sign_out <= VN_sign_out( 6917 downto 6912 );
    VN1153_data_out <= VN_data_out( 6923 downto 6918 );
    VN1153_sign_out <= VN_sign_out( 6923 downto 6918 );
    VN1154_data_out <= VN_data_out( 6929 downto 6924 );
    VN1154_sign_out <= VN_sign_out( 6929 downto 6924 );
    VN1155_data_out <= VN_data_out( 6935 downto 6930 );
    VN1155_sign_out <= VN_sign_out( 6935 downto 6930 );
    VN1156_data_out <= VN_data_out( 6941 downto 6936 );
    VN1156_sign_out <= VN_sign_out( 6941 downto 6936 );
    VN1157_data_out <= VN_data_out( 6947 downto 6942 );
    VN1157_sign_out <= VN_sign_out( 6947 downto 6942 );
    VN1158_data_out <= VN_data_out( 6953 downto 6948 );
    VN1158_sign_out <= VN_sign_out( 6953 downto 6948 );
    VN1159_data_out <= VN_data_out( 6959 downto 6954 );
    VN1159_sign_out <= VN_sign_out( 6959 downto 6954 );
    VN1160_data_out <= VN_data_out( 6965 downto 6960 );
    VN1160_sign_out <= VN_sign_out( 6965 downto 6960 );
    VN1161_data_out <= VN_data_out( 6971 downto 6966 );
    VN1161_sign_out <= VN_sign_out( 6971 downto 6966 );
    VN1162_data_out <= VN_data_out( 6977 downto 6972 );
    VN1162_sign_out <= VN_sign_out( 6977 downto 6972 );
    VN1163_data_out <= VN_data_out( 6983 downto 6978 );
    VN1163_sign_out <= VN_sign_out( 6983 downto 6978 );
    VN1164_data_out <= VN_data_out( 6989 downto 6984 );
    VN1164_sign_out <= VN_sign_out( 6989 downto 6984 );
    VN1165_data_out <= VN_data_out( 6995 downto 6990 );
    VN1165_sign_out <= VN_sign_out( 6995 downto 6990 );
    VN1166_data_out <= VN_data_out( 7001 downto 6996 );
    VN1166_sign_out <= VN_sign_out( 7001 downto 6996 );
    VN1167_data_out <= VN_data_out( 7007 downto 7002 );
    VN1167_sign_out <= VN_sign_out( 7007 downto 7002 );
    VN1168_data_out <= VN_data_out( 7013 downto 7008 );
    VN1168_sign_out <= VN_sign_out( 7013 downto 7008 );
    VN1169_data_out <= VN_data_out( 7019 downto 7014 );
    VN1169_sign_out <= VN_sign_out( 7019 downto 7014 );
    VN1170_data_out <= VN_data_out( 7025 downto 7020 );
    VN1170_sign_out <= VN_sign_out( 7025 downto 7020 );
    VN1171_data_out <= VN_data_out( 7031 downto 7026 );
    VN1171_sign_out <= VN_sign_out( 7031 downto 7026 );
    VN1172_data_out <= VN_data_out( 7037 downto 7032 );
    VN1172_sign_out <= VN_sign_out( 7037 downto 7032 );
    VN1173_data_out <= VN_data_out( 7043 downto 7038 );
    VN1173_sign_out <= VN_sign_out( 7043 downto 7038 );
    VN1174_data_out <= VN_data_out( 7049 downto 7044 );
    VN1174_sign_out <= VN_sign_out( 7049 downto 7044 );
    VN1175_data_out <= VN_data_out( 7055 downto 7050 );
    VN1175_sign_out <= VN_sign_out( 7055 downto 7050 );
    VN1176_data_out <= VN_data_out( 7061 downto 7056 );
    VN1176_sign_out <= VN_sign_out( 7061 downto 7056 );
    VN1177_data_out <= VN_data_out( 7067 downto 7062 );
    VN1177_sign_out <= VN_sign_out( 7067 downto 7062 );
    VN1178_data_out <= VN_data_out( 7073 downto 7068 );
    VN1178_sign_out <= VN_sign_out( 7073 downto 7068 );
    VN1179_data_out <= VN_data_out( 7079 downto 7074 );
    VN1179_sign_out <= VN_sign_out( 7079 downto 7074 );
    VN1180_data_out <= VN_data_out( 7085 downto 7080 );
    VN1180_sign_out <= VN_sign_out( 7085 downto 7080 );
    VN1181_data_out <= VN_data_out( 7091 downto 7086 );
    VN1181_sign_out <= VN_sign_out( 7091 downto 7086 );
    VN1182_data_out <= VN_data_out( 7097 downto 7092 );
    VN1182_sign_out <= VN_sign_out( 7097 downto 7092 );
    VN1183_data_out <= VN_data_out( 7103 downto 7098 );
    VN1183_sign_out <= VN_sign_out( 7103 downto 7098 );
    VN1184_data_out <= VN_data_out( 7109 downto 7104 );
    VN1184_sign_out <= VN_sign_out( 7109 downto 7104 );
    VN1185_data_out <= VN_data_out( 7115 downto 7110 );
    VN1185_sign_out <= VN_sign_out( 7115 downto 7110 );
    VN1186_data_out <= VN_data_out( 7121 downto 7116 );
    VN1186_sign_out <= VN_sign_out( 7121 downto 7116 );
    VN1187_data_out <= VN_data_out( 7127 downto 7122 );
    VN1187_sign_out <= VN_sign_out( 7127 downto 7122 );
    VN1188_data_out <= VN_data_out( 7133 downto 7128 );
    VN1188_sign_out <= VN_sign_out( 7133 downto 7128 );
    VN1189_data_out <= VN_data_out( 7139 downto 7134 );
    VN1189_sign_out <= VN_sign_out( 7139 downto 7134 );
    VN1190_data_out <= VN_data_out( 7145 downto 7140 );
    VN1190_sign_out <= VN_sign_out( 7145 downto 7140 );
    VN1191_data_out <= VN_data_out( 7151 downto 7146 );
    VN1191_sign_out <= VN_sign_out( 7151 downto 7146 );
    VN1192_data_out <= VN_data_out( 7157 downto 7152 );
    VN1192_sign_out <= VN_sign_out( 7157 downto 7152 );
    VN1193_data_out <= VN_data_out( 7163 downto 7158 );
    VN1193_sign_out <= VN_sign_out( 7163 downto 7158 );
    VN1194_data_out <= VN_data_out( 7169 downto 7164 );
    VN1194_sign_out <= VN_sign_out( 7169 downto 7164 );
    VN1195_data_out <= VN_data_out( 7175 downto 7170 );
    VN1195_sign_out <= VN_sign_out( 7175 downto 7170 );
    VN1196_data_out <= VN_data_out( 7181 downto 7176 );
    VN1196_sign_out <= VN_sign_out( 7181 downto 7176 );
    VN1197_data_out <= VN_data_out( 7187 downto 7182 );
    VN1197_sign_out <= VN_sign_out( 7187 downto 7182 );
    VN1198_data_out <= VN_data_out( 7193 downto 7188 );
    VN1198_sign_out <= VN_sign_out( 7193 downto 7188 );
    VN1199_data_out <= VN_data_out( 7199 downto 7194 );
    VN1199_sign_out <= VN_sign_out( 7199 downto 7194 );
    VN1200_data_out <= VN_data_out( 7205 downto 7200 );
    VN1200_sign_out <= VN_sign_out( 7205 downto 7200 );
    VN1201_data_out <= VN_data_out( 7211 downto 7206 );
    VN1201_sign_out <= VN_sign_out( 7211 downto 7206 );
    VN1202_data_out <= VN_data_out( 7217 downto 7212 );
    VN1202_sign_out <= VN_sign_out( 7217 downto 7212 );
    VN1203_data_out <= VN_data_out( 7223 downto 7218 );
    VN1203_sign_out <= VN_sign_out( 7223 downto 7218 );
    VN1204_data_out <= VN_data_out( 7229 downto 7224 );
    VN1204_sign_out <= VN_sign_out( 7229 downto 7224 );
    VN1205_data_out <= VN_data_out( 7235 downto 7230 );
    VN1205_sign_out <= VN_sign_out( 7235 downto 7230 );
    VN1206_data_out <= VN_data_out( 7241 downto 7236 );
    VN1206_sign_out <= VN_sign_out( 7241 downto 7236 );
    VN1207_data_out <= VN_data_out( 7247 downto 7242 );
    VN1207_sign_out <= VN_sign_out( 7247 downto 7242 );
    VN1208_data_out <= VN_data_out( 7253 downto 7248 );
    VN1208_sign_out <= VN_sign_out( 7253 downto 7248 );
    VN1209_data_out <= VN_data_out( 7259 downto 7254 );
    VN1209_sign_out <= VN_sign_out( 7259 downto 7254 );
    VN1210_data_out <= VN_data_out( 7265 downto 7260 );
    VN1210_sign_out <= VN_sign_out( 7265 downto 7260 );
    VN1211_data_out <= VN_data_out( 7271 downto 7266 );
    VN1211_sign_out <= VN_sign_out( 7271 downto 7266 );
    VN1212_data_out <= VN_data_out( 7277 downto 7272 );
    VN1212_sign_out <= VN_sign_out( 7277 downto 7272 );
    VN1213_data_out <= VN_data_out( 7283 downto 7278 );
    VN1213_sign_out <= VN_sign_out( 7283 downto 7278 );
    VN1214_data_out <= VN_data_out( 7289 downto 7284 );
    VN1214_sign_out <= VN_sign_out( 7289 downto 7284 );
    VN1215_data_out <= VN_data_out( 7295 downto 7290 );
    VN1215_sign_out <= VN_sign_out( 7295 downto 7290 );
    VN1216_data_out <= VN_data_out( 7301 downto 7296 );
    VN1216_sign_out <= VN_sign_out( 7301 downto 7296 );
    VN1217_data_out <= VN_data_out( 7307 downto 7302 );
    VN1217_sign_out <= VN_sign_out( 7307 downto 7302 );
    VN1218_data_out <= VN_data_out( 7313 downto 7308 );
    VN1218_sign_out <= VN_sign_out( 7313 downto 7308 );
    VN1219_data_out <= VN_data_out( 7319 downto 7314 );
    VN1219_sign_out <= VN_sign_out( 7319 downto 7314 );
    VN1220_data_out <= VN_data_out( 7325 downto 7320 );
    VN1220_sign_out <= VN_sign_out( 7325 downto 7320 );
    VN1221_data_out <= VN_data_out( 7331 downto 7326 );
    VN1221_sign_out <= VN_sign_out( 7331 downto 7326 );
    VN1222_data_out <= VN_data_out( 7337 downto 7332 );
    VN1222_sign_out <= VN_sign_out( 7337 downto 7332 );
    VN1223_data_out <= VN_data_out( 7343 downto 7338 );
    VN1223_sign_out <= VN_sign_out( 7343 downto 7338 );
    VN1224_data_out <= VN_data_out( 7349 downto 7344 );
    VN1224_sign_out <= VN_sign_out( 7349 downto 7344 );
    VN1225_data_out <= VN_data_out( 7355 downto 7350 );
    VN1225_sign_out <= VN_sign_out( 7355 downto 7350 );
    VN1226_data_out <= VN_data_out( 7361 downto 7356 );
    VN1226_sign_out <= VN_sign_out( 7361 downto 7356 );
    VN1227_data_out <= VN_data_out( 7367 downto 7362 );
    VN1227_sign_out <= VN_sign_out( 7367 downto 7362 );
    VN1228_data_out <= VN_data_out( 7373 downto 7368 );
    VN1228_sign_out <= VN_sign_out( 7373 downto 7368 );
    VN1229_data_out <= VN_data_out( 7379 downto 7374 );
    VN1229_sign_out <= VN_sign_out( 7379 downto 7374 );
    VN1230_data_out <= VN_data_out( 7385 downto 7380 );
    VN1230_sign_out <= VN_sign_out( 7385 downto 7380 );
    VN1231_data_out <= VN_data_out( 7391 downto 7386 );
    VN1231_sign_out <= VN_sign_out( 7391 downto 7386 );
    VN1232_data_out <= VN_data_out( 7397 downto 7392 );
    VN1232_sign_out <= VN_sign_out( 7397 downto 7392 );
    VN1233_data_out <= VN_data_out( 7403 downto 7398 );
    VN1233_sign_out <= VN_sign_out( 7403 downto 7398 );
    VN1234_data_out <= VN_data_out( 7409 downto 7404 );
    VN1234_sign_out <= VN_sign_out( 7409 downto 7404 );
    VN1235_data_out <= VN_data_out( 7415 downto 7410 );
    VN1235_sign_out <= VN_sign_out( 7415 downto 7410 );
    VN1236_data_out <= VN_data_out( 7421 downto 7416 );
    VN1236_sign_out <= VN_sign_out( 7421 downto 7416 );
    VN1237_data_out <= VN_data_out( 7427 downto 7422 );
    VN1237_sign_out <= VN_sign_out( 7427 downto 7422 );
    VN1238_data_out <= VN_data_out( 7433 downto 7428 );
    VN1238_sign_out <= VN_sign_out( 7433 downto 7428 );
    VN1239_data_out <= VN_data_out( 7439 downto 7434 );
    VN1239_sign_out <= VN_sign_out( 7439 downto 7434 );
    VN1240_data_out <= VN_data_out( 7445 downto 7440 );
    VN1240_sign_out <= VN_sign_out( 7445 downto 7440 );
    VN1241_data_out <= VN_data_out( 7451 downto 7446 );
    VN1241_sign_out <= VN_sign_out( 7451 downto 7446 );
    VN1242_data_out <= VN_data_out( 7457 downto 7452 );
    VN1242_sign_out <= VN_sign_out( 7457 downto 7452 );
    VN1243_data_out <= VN_data_out( 7463 downto 7458 );
    VN1243_sign_out <= VN_sign_out( 7463 downto 7458 );
    VN1244_data_out <= VN_data_out( 7469 downto 7464 );
    VN1244_sign_out <= VN_sign_out( 7469 downto 7464 );
    VN1245_data_out <= VN_data_out( 7475 downto 7470 );
    VN1245_sign_out <= VN_sign_out( 7475 downto 7470 );
    VN1246_data_out <= VN_data_out( 7481 downto 7476 );
    VN1246_sign_out <= VN_sign_out( 7481 downto 7476 );
    VN1247_data_out <= VN_data_out( 7487 downto 7482 );
    VN1247_sign_out <= VN_sign_out( 7487 downto 7482 );
    VN1248_data_out <= VN_data_out( 7493 downto 7488 );
    VN1248_sign_out <= VN_sign_out( 7493 downto 7488 );
    VN1249_data_out <= VN_data_out( 7499 downto 7494 );
    VN1249_sign_out <= VN_sign_out( 7499 downto 7494 );
    VN1250_data_out <= VN_data_out( 7505 downto 7500 );
    VN1250_sign_out <= VN_sign_out( 7505 downto 7500 );
    VN1251_data_out <= VN_data_out( 7511 downto 7506 );
    VN1251_sign_out <= VN_sign_out( 7511 downto 7506 );
    VN1252_data_out <= VN_data_out( 7517 downto 7512 );
    VN1252_sign_out <= VN_sign_out( 7517 downto 7512 );
    VN1253_data_out <= VN_data_out( 7523 downto 7518 );
    VN1253_sign_out <= VN_sign_out( 7523 downto 7518 );
    VN1254_data_out <= VN_data_out( 7529 downto 7524 );
    VN1254_sign_out <= VN_sign_out( 7529 downto 7524 );
    VN1255_data_out <= VN_data_out( 7535 downto 7530 );
    VN1255_sign_out <= VN_sign_out( 7535 downto 7530 );
    VN1256_data_out <= VN_data_out( 7541 downto 7536 );
    VN1256_sign_out <= VN_sign_out( 7541 downto 7536 );
    VN1257_data_out <= VN_data_out( 7547 downto 7542 );
    VN1257_sign_out <= VN_sign_out( 7547 downto 7542 );
    VN1258_data_out <= VN_data_out( 7553 downto 7548 );
    VN1258_sign_out <= VN_sign_out( 7553 downto 7548 );
    VN1259_data_out <= VN_data_out( 7559 downto 7554 );
    VN1259_sign_out <= VN_sign_out( 7559 downto 7554 );
    VN1260_data_out <= VN_data_out( 7565 downto 7560 );
    VN1260_sign_out <= VN_sign_out( 7565 downto 7560 );
    VN1261_data_out <= VN_data_out( 7571 downto 7566 );
    VN1261_sign_out <= VN_sign_out( 7571 downto 7566 );
    VN1262_data_out <= VN_data_out( 7577 downto 7572 );
    VN1262_sign_out <= VN_sign_out( 7577 downto 7572 );
    VN1263_data_out <= VN_data_out( 7583 downto 7578 );
    VN1263_sign_out <= VN_sign_out( 7583 downto 7578 );
    VN1264_data_out <= VN_data_out( 7589 downto 7584 );
    VN1264_sign_out <= VN_sign_out( 7589 downto 7584 );
    VN1265_data_out <= VN_data_out( 7595 downto 7590 );
    VN1265_sign_out <= VN_sign_out( 7595 downto 7590 );
    VN1266_data_out <= VN_data_out( 7601 downto 7596 );
    VN1266_sign_out <= VN_sign_out( 7601 downto 7596 );
    VN1267_data_out <= VN_data_out( 7607 downto 7602 );
    VN1267_sign_out <= VN_sign_out( 7607 downto 7602 );
    VN1268_data_out <= VN_data_out( 7613 downto 7608 );
    VN1268_sign_out <= VN_sign_out( 7613 downto 7608 );
    VN1269_data_out <= VN_data_out( 7619 downto 7614 );
    VN1269_sign_out <= VN_sign_out( 7619 downto 7614 );
    VN1270_data_out <= VN_data_out( 7625 downto 7620 );
    VN1270_sign_out <= VN_sign_out( 7625 downto 7620 );
    VN1271_data_out <= VN_data_out( 7631 downto 7626 );
    VN1271_sign_out <= VN_sign_out( 7631 downto 7626 );
    VN1272_data_out <= VN_data_out( 7637 downto 7632 );
    VN1272_sign_out <= VN_sign_out( 7637 downto 7632 );
    VN1273_data_out <= VN_data_out( 7643 downto 7638 );
    VN1273_sign_out <= VN_sign_out( 7643 downto 7638 );
    VN1274_data_out <= VN_data_out( 7649 downto 7644 );
    VN1274_sign_out <= VN_sign_out( 7649 downto 7644 );
    VN1275_data_out <= VN_data_out( 7655 downto 7650 );
    VN1275_sign_out <= VN_sign_out( 7655 downto 7650 );
    VN1276_data_out <= VN_data_out( 7661 downto 7656 );
    VN1276_sign_out <= VN_sign_out( 7661 downto 7656 );
    VN1277_data_out <= VN_data_out( 7667 downto 7662 );
    VN1277_sign_out <= VN_sign_out( 7667 downto 7662 );
    VN1278_data_out <= VN_data_out( 7673 downto 7668 );
    VN1278_sign_out <= VN_sign_out( 7673 downto 7668 );
    VN1279_data_out <= VN_data_out( 7679 downto 7674 );
    VN1279_sign_out <= VN_sign_out( 7679 downto 7674 );
    VN1280_data_out <= VN_data_out( 7685 downto 7680 );
    VN1280_sign_out <= VN_sign_out( 7685 downto 7680 );
    VN1281_data_out <= VN_data_out( 7691 downto 7686 );
    VN1281_sign_out <= VN_sign_out( 7691 downto 7686 );
    VN1282_data_out <= VN_data_out( 7697 downto 7692 );
    VN1282_sign_out <= VN_sign_out( 7697 downto 7692 );
    VN1283_data_out <= VN_data_out( 7703 downto 7698 );
    VN1283_sign_out <= VN_sign_out( 7703 downto 7698 );
    VN1284_data_out <= VN_data_out( 7709 downto 7704 );
    VN1284_sign_out <= VN_sign_out( 7709 downto 7704 );
    VN1285_data_out <= VN_data_out( 7715 downto 7710 );
    VN1285_sign_out <= VN_sign_out( 7715 downto 7710 );
    VN1286_data_out <= VN_data_out( 7721 downto 7716 );
    VN1286_sign_out <= VN_sign_out( 7721 downto 7716 );
    VN1287_data_out <= VN_data_out( 7727 downto 7722 );
    VN1287_sign_out <= VN_sign_out( 7727 downto 7722 );
    VN1288_data_out <= VN_data_out( 7733 downto 7728 );
    VN1288_sign_out <= VN_sign_out( 7733 downto 7728 );
    VN1289_data_out <= VN_data_out( 7739 downto 7734 );
    VN1289_sign_out <= VN_sign_out( 7739 downto 7734 );
    VN1290_data_out <= VN_data_out( 7745 downto 7740 );
    VN1290_sign_out <= VN_sign_out( 7745 downto 7740 );
    VN1291_data_out <= VN_data_out( 7751 downto 7746 );
    VN1291_sign_out <= VN_sign_out( 7751 downto 7746 );
    VN1292_data_out <= VN_data_out( 7757 downto 7752 );
    VN1292_sign_out <= VN_sign_out( 7757 downto 7752 );
    VN1293_data_out <= VN_data_out( 7763 downto 7758 );
    VN1293_sign_out <= VN_sign_out( 7763 downto 7758 );
    VN1294_data_out <= VN_data_out( 7769 downto 7764 );
    VN1294_sign_out <= VN_sign_out( 7769 downto 7764 );
    VN1295_data_out <= VN_data_out( 7775 downto 7770 );
    VN1295_sign_out <= VN_sign_out( 7775 downto 7770 );
    VN1296_data_out <= VN_data_out( 7781 downto 7776 );
    VN1296_sign_out <= VN_sign_out( 7781 downto 7776 );
    VN1297_data_out <= VN_data_out( 7787 downto 7782 );
    VN1297_sign_out <= VN_sign_out( 7787 downto 7782 );
    VN1298_data_out <= VN_data_out( 7793 downto 7788 );
    VN1298_sign_out <= VN_sign_out( 7793 downto 7788 );
    VN1299_data_out <= VN_data_out( 7799 downto 7794 );
    VN1299_sign_out <= VN_sign_out( 7799 downto 7794 );
    VN1300_data_out <= VN_data_out( 7805 downto 7800 );
    VN1300_sign_out <= VN_sign_out( 7805 downto 7800 );
    VN1301_data_out <= VN_data_out( 7811 downto 7806 );
    VN1301_sign_out <= VN_sign_out( 7811 downto 7806 );
    VN1302_data_out <= VN_data_out( 7817 downto 7812 );
    VN1302_sign_out <= VN_sign_out( 7817 downto 7812 );
    VN1303_data_out <= VN_data_out( 7823 downto 7818 );
    VN1303_sign_out <= VN_sign_out( 7823 downto 7818 );
    VN1304_data_out <= VN_data_out( 7829 downto 7824 );
    VN1304_sign_out <= VN_sign_out( 7829 downto 7824 );
    VN1305_data_out <= VN_data_out( 7835 downto 7830 );
    VN1305_sign_out <= VN_sign_out( 7835 downto 7830 );
    VN1306_data_out <= VN_data_out( 7841 downto 7836 );
    VN1306_sign_out <= VN_sign_out( 7841 downto 7836 );
    VN1307_data_out <= VN_data_out( 7847 downto 7842 );
    VN1307_sign_out <= VN_sign_out( 7847 downto 7842 );
    VN1308_data_out <= VN_data_out( 7853 downto 7848 );
    VN1308_sign_out <= VN_sign_out( 7853 downto 7848 );
    VN1309_data_out <= VN_data_out( 7859 downto 7854 );
    VN1309_sign_out <= VN_sign_out( 7859 downto 7854 );
    VN1310_data_out <= VN_data_out( 7865 downto 7860 );
    VN1310_sign_out <= VN_sign_out( 7865 downto 7860 );
    VN1311_data_out <= VN_data_out( 7871 downto 7866 );
    VN1311_sign_out <= VN_sign_out( 7871 downto 7866 );
    VN1312_data_out <= VN_data_out( 7877 downto 7872 );
    VN1312_sign_out <= VN_sign_out( 7877 downto 7872 );
    VN1313_data_out <= VN_data_out( 7883 downto 7878 );
    VN1313_sign_out <= VN_sign_out( 7883 downto 7878 );
    VN1314_data_out <= VN_data_out( 7889 downto 7884 );
    VN1314_sign_out <= VN_sign_out( 7889 downto 7884 );
    VN1315_data_out <= VN_data_out( 7895 downto 7890 );
    VN1315_sign_out <= VN_sign_out( 7895 downto 7890 );
    VN1316_data_out <= VN_data_out( 7901 downto 7896 );
    VN1316_sign_out <= VN_sign_out( 7901 downto 7896 );
    VN1317_data_out <= VN_data_out( 7907 downto 7902 );
    VN1317_sign_out <= VN_sign_out( 7907 downto 7902 );
    VN1318_data_out <= VN_data_out( 7913 downto 7908 );
    VN1318_sign_out <= VN_sign_out( 7913 downto 7908 );
    VN1319_data_out <= VN_data_out( 7919 downto 7914 );
    VN1319_sign_out <= VN_sign_out( 7919 downto 7914 );
    VN1320_data_out <= VN_data_out( 7925 downto 7920 );
    VN1320_sign_out <= VN_sign_out( 7925 downto 7920 );
    VN1321_data_out <= VN_data_out( 7931 downto 7926 );
    VN1321_sign_out <= VN_sign_out( 7931 downto 7926 );
    VN1322_data_out <= VN_data_out( 7937 downto 7932 );
    VN1322_sign_out <= VN_sign_out( 7937 downto 7932 );
    VN1323_data_out <= VN_data_out( 7943 downto 7938 );
    VN1323_sign_out <= VN_sign_out( 7943 downto 7938 );
    VN1324_data_out <= VN_data_out( 7949 downto 7944 );
    VN1324_sign_out <= VN_sign_out( 7949 downto 7944 );
    VN1325_data_out <= VN_data_out( 7955 downto 7950 );
    VN1325_sign_out <= VN_sign_out( 7955 downto 7950 );
    VN1326_data_out <= VN_data_out( 7961 downto 7956 );
    VN1326_sign_out <= VN_sign_out( 7961 downto 7956 );
    VN1327_data_out <= VN_data_out( 7967 downto 7962 );
    VN1327_sign_out <= VN_sign_out( 7967 downto 7962 );
    VN1328_data_out <= VN_data_out( 7973 downto 7968 );
    VN1328_sign_out <= VN_sign_out( 7973 downto 7968 );
    VN1329_data_out <= VN_data_out( 7979 downto 7974 );
    VN1329_sign_out <= VN_sign_out( 7979 downto 7974 );
    VN1330_data_out <= VN_data_out( 7985 downto 7980 );
    VN1330_sign_out <= VN_sign_out( 7985 downto 7980 );
    VN1331_data_out <= VN_data_out( 7991 downto 7986 );
    VN1331_sign_out <= VN_sign_out( 7991 downto 7986 );
    VN1332_data_out <= VN_data_out( 7997 downto 7992 );
    VN1332_sign_out <= VN_sign_out( 7997 downto 7992 );
    VN1333_data_out <= VN_data_out( 8003 downto 7998 );
    VN1333_sign_out <= VN_sign_out( 8003 downto 7998 );
    VN1334_data_out <= VN_data_out( 8009 downto 8004 );
    VN1334_sign_out <= VN_sign_out( 8009 downto 8004 );
    VN1335_data_out <= VN_data_out( 8015 downto 8010 );
    VN1335_sign_out <= VN_sign_out( 8015 downto 8010 );
    VN1336_data_out <= VN_data_out( 8021 downto 8016 );
    VN1336_sign_out <= VN_sign_out( 8021 downto 8016 );
    VN1337_data_out <= VN_data_out( 8027 downto 8022 );
    VN1337_sign_out <= VN_sign_out( 8027 downto 8022 );
    VN1338_data_out <= VN_data_out( 8033 downto 8028 );
    VN1338_sign_out <= VN_sign_out( 8033 downto 8028 );
    VN1339_data_out <= VN_data_out( 8039 downto 8034 );
    VN1339_sign_out <= VN_sign_out( 8039 downto 8034 );
    VN1340_data_out <= VN_data_out( 8045 downto 8040 );
    VN1340_sign_out <= VN_sign_out( 8045 downto 8040 );
    VN1341_data_out <= VN_data_out( 8051 downto 8046 );
    VN1341_sign_out <= VN_sign_out( 8051 downto 8046 );
    VN1342_data_out <= VN_data_out( 8057 downto 8052 );
    VN1342_sign_out <= VN_sign_out( 8057 downto 8052 );
    VN1343_data_out <= VN_data_out( 8063 downto 8058 );
    VN1343_sign_out <= VN_sign_out( 8063 downto 8058 );
    VN1344_data_out <= VN_data_out( 8069 downto 8064 );
    VN1344_sign_out <= VN_sign_out( 8069 downto 8064 );
    VN1345_data_out <= VN_data_out( 8075 downto 8070 );
    VN1345_sign_out <= VN_sign_out( 8075 downto 8070 );
    VN1346_data_out <= VN_data_out( 8081 downto 8076 );
    VN1346_sign_out <= VN_sign_out( 8081 downto 8076 );
    VN1347_data_out <= VN_data_out( 8087 downto 8082 );
    VN1347_sign_out <= VN_sign_out( 8087 downto 8082 );
    VN1348_data_out <= VN_data_out( 8093 downto 8088 );
    VN1348_sign_out <= VN_sign_out( 8093 downto 8088 );
    VN1349_data_out <= VN_data_out( 8099 downto 8094 );
    VN1349_sign_out <= VN_sign_out( 8099 downto 8094 );
    VN1350_data_out <= VN_data_out( 8105 downto 8100 );
    VN1350_sign_out <= VN_sign_out( 8105 downto 8100 );
    VN1351_data_out <= VN_data_out( 8111 downto 8106 );
    VN1351_sign_out <= VN_sign_out( 8111 downto 8106 );
    VN1352_data_out <= VN_data_out( 8117 downto 8112 );
    VN1352_sign_out <= VN_sign_out( 8117 downto 8112 );
    VN1353_data_out <= VN_data_out( 8123 downto 8118 );
    VN1353_sign_out <= VN_sign_out( 8123 downto 8118 );
    VN1354_data_out <= VN_data_out( 8129 downto 8124 );
    VN1354_sign_out <= VN_sign_out( 8129 downto 8124 );
    VN1355_data_out <= VN_data_out( 8135 downto 8130 );
    VN1355_sign_out <= VN_sign_out( 8135 downto 8130 );
    VN1356_data_out <= VN_data_out( 8141 downto 8136 );
    VN1356_sign_out <= VN_sign_out( 8141 downto 8136 );
    VN1357_data_out <= VN_data_out( 8147 downto 8142 );
    VN1357_sign_out <= VN_sign_out( 8147 downto 8142 );
    VN1358_data_out <= VN_data_out( 8153 downto 8148 );
    VN1358_sign_out <= VN_sign_out( 8153 downto 8148 );
    VN1359_data_out <= VN_data_out( 8159 downto 8154 );
    VN1359_sign_out <= VN_sign_out( 8159 downto 8154 );
    VN1360_data_out <= VN_data_out( 8165 downto 8160 );
    VN1360_sign_out <= VN_sign_out( 8165 downto 8160 );
    VN1361_data_out <= VN_data_out( 8171 downto 8166 );
    VN1361_sign_out <= VN_sign_out( 8171 downto 8166 );
    VN1362_data_out <= VN_data_out( 8177 downto 8172 );
    VN1362_sign_out <= VN_sign_out( 8177 downto 8172 );
    VN1363_data_out <= VN_data_out( 8183 downto 8178 );
    VN1363_sign_out <= VN_sign_out( 8183 downto 8178 );
    VN1364_data_out <= VN_data_out( 8189 downto 8184 );
    VN1364_sign_out <= VN_sign_out( 8189 downto 8184 );
    VN1365_data_out <= VN_data_out( 8195 downto 8190 );
    VN1365_sign_out <= VN_sign_out( 8195 downto 8190 );
    VN1366_data_out <= VN_data_out( 8201 downto 8196 );
    VN1366_sign_out <= VN_sign_out( 8201 downto 8196 );
    VN1367_data_out <= VN_data_out( 8207 downto 8202 );
    VN1367_sign_out <= VN_sign_out( 8207 downto 8202 );
    VN1368_data_out <= VN_data_out( 8213 downto 8208 );
    VN1368_sign_out <= VN_sign_out( 8213 downto 8208 );
    VN1369_data_out <= VN_data_out( 8219 downto 8214 );
    VN1369_sign_out <= VN_sign_out( 8219 downto 8214 );
    VN1370_data_out <= VN_data_out( 8225 downto 8220 );
    VN1370_sign_out <= VN_sign_out( 8225 downto 8220 );
    VN1371_data_out <= VN_data_out( 8231 downto 8226 );
    VN1371_sign_out <= VN_sign_out( 8231 downto 8226 );
    VN1372_data_out <= VN_data_out( 8237 downto 8232 );
    VN1372_sign_out <= VN_sign_out( 8237 downto 8232 );
    VN1373_data_out <= VN_data_out( 8243 downto 8238 );
    VN1373_sign_out <= VN_sign_out( 8243 downto 8238 );
    VN1374_data_out <= VN_data_out( 8249 downto 8244 );
    VN1374_sign_out <= VN_sign_out( 8249 downto 8244 );
    VN1375_data_out <= VN_data_out( 8255 downto 8250 );
    VN1375_sign_out <= VN_sign_out( 8255 downto 8250 );
    VN1376_data_out <= VN_data_out( 8261 downto 8256 );
    VN1376_sign_out <= VN_sign_out( 8261 downto 8256 );
    VN1377_data_out <= VN_data_out( 8267 downto 8262 );
    VN1377_sign_out <= VN_sign_out( 8267 downto 8262 );
    VN1378_data_out <= VN_data_out( 8273 downto 8268 );
    VN1378_sign_out <= VN_sign_out( 8273 downto 8268 );
    VN1379_data_out <= VN_data_out( 8279 downto 8274 );
    VN1379_sign_out <= VN_sign_out( 8279 downto 8274 );
    VN1380_data_out <= VN_data_out( 8285 downto 8280 );
    VN1380_sign_out <= VN_sign_out( 8285 downto 8280 );
    VN1381_data_out <= VN_data_out( 8291 downto 8286 );
    VN1381_sign_out <= VN_sign_out( 8291 downto 8286 );
    VN1382_data_out <= VN_data_out( 8297 downto 8292 );
    VN1382_sign_out <= VN_sign_out( 8297 downto 8292 );
    VN1383_data_out <= VN_data_out( 8303 downto 8298 );
    VN1383_sign_out <= VN_sign_out( 8303 downto 8298 );
    VN1384_data_out <= VN_data_out( 8309 downto 8304 );
    VN1384_sign_out <= VN_sign_out( 8309 downto 8304 );
    VN1385_data_out <= VN_data_out( 8315 downto 8310 );
    VN1385_sign_out <= VN_sign_out( 8315 downto 8310 );
    VN1386_data_out <= VN_data_out( 8321 downto 8316 );
    VN1386_sign_out <= VN_sign_out( 8321 downto 8316 );
    VN1387_data_out <= VN_data_out( 8327 downto 8322 );
    VN1387_sign_out <= VN_sign_out( 8327 downto 8322 );
    VN1388_data_out <= VN_data_out( 8333 downto 8328 );
    VN1388_sign_out <= VN_sign_out( 8333 downto 8328 );
    VN1389_data_out <= VN_data_out( 8339 downto 8334 );
    VN1389_sign_out <= VN_sign_out( 8339 downto 8334 );
    VN1390_data_out <= VN_data_out( 8345 downto 8340 );
    VN1390_sign_out <= VN_sign_out( 8345 downto 8340 );
    VN1391_data_out <= VN_data_out( 8351 downto 8346 );
    VN1391_sign_out <= VN_sign_out( 8351 downto 8346 );
    VN1392_data_out <= VN_data_out( 8357 downto 8352 );
    VN1392_sign_out <= VN_sign_out( 8357 downto 8352 );
    VN1393_data_out <= VN_data_out( 8363 downto 8358 );
    VN1393_sign_out <= VN_sign_out( 8363 downto 8358 );
    VN1394_data_out <= VN_data_out( 8369 downto 8364 );
    VN1394_sign_out <= VN_sign_out( 8369 downto 8364 );
    VN1395_data_out <= VN_data_out( 8375 downto 8370 );
    VN1395_sign_out <= VN_sign_out( 8375 downto 8370 );
    VN1396_data_out <= VN_data_out( 8381 downto 8376 );
    VN1396_sign_out <= VN_sign_out( 8381 downto 8376 );
    VN1397_data_out <= VN_data_out( 8387 downto 8382 );
    VN1397_sign_out <= VN_sign_out( 8387 downto 8382 );
    VN1398_data_out <= VN_data_out( 8393 downto 8388 );
    VN1398_sign_out <= VN_sign_out( 8393 downto 8388 );
    VN1399_data_out <= VN_data_out( 8399 downto 8394 );
    VN1399_sign_out <= VN_sign_out( 8399 downto 8394 );
    VN1400_data_out <= VN_data_out( 8405 downto 8400 );
    VN1400_sign_out <= VN_sign_out( 8405 downto 8400 );
    VN1401_data_out <= VN_data_out( 8411 downto 8406 );
    VN1401_sign_out <= VN_sign_out( 8411 downto 8406 );
    VN1402_data_out <= VN_data_out( 8417 downto 8412 );
    VN1402_sign_out <= VN_sign_out( 8417 downto 8412 );
    VN1403_data_out <= VN_data_out( 8423 downto 8418 );
    VN1403_sign_out <= VN_sign_out( 8423 downto 8418 );
    VN1404_data_out <= VN_data_out( 8429 downto 8424 );
    VN1404_sign_out <= VN_sign_out( 8429 downto 8424 );
    VN1405_data_out <= VN_data_out( 8435 downto 8430 );
    VN1405_sign_out <= VN_sign_out( 8435 downto 8430 );
    VN1406_data_out <= VN_data_out( 8441 downto 8436 );
    VN1406_sign_out <= VN_sign_out( 8441 downto 8436 );
    VN1407_data_out <= VN_data_out( 8447 downto 8442 );
    VN1407_sign_out <= VN_sign_out( 8447 downto 8442 );
    VN1408_data_out <= VN_data_out( 8453 downto 8448 );
    VN1408_sign_out <= VN_sign_out( 8453 downto 8448 );
    VN1409_data_out <= VN_data_out( 8459 downto 8454 );
    VN1409_sign_out <= VN_sign_out( 8459 downto 8454 );
    VN1410_data_out <= VN_data_out( 8465 downto 8460 );
    VN1410_sign_out <= VN_sign_out( 8465 downto 8460 );
    VN1411_data_out <= VN_data_out( 8471 downto 8466 );
    VN1411_sign_out <= VN_sign_out( 8471 downto 8466 );
    VN1412_data_out <= VN_data_out( 8477 downto 8472 );
    VN1412_sign_out <= VN_sign_out( 8477 downto 8472 );
    VN1413_data_out <= VN_data_out( 8483 downto 8478 );
    VN1413_sign_out <= VN_sign_out( 8483 downto 8478 );
    VN1414_data_out <= VN_data_out( 8489 downto 8484 );
    VN1414_sign_out <= VN_sign_out( 8489 downto 8484 );
    VN1415_data_out <= VN_data_out( 8495 downto 8490 );
    VN1415_sign_out <= VN_sign_out( 8495 downto 8490 );
    VN1416_data_out <= VN_data_out( 8501 downto 8496 );
    VN1416_sign_out <= VN_sign_out( 8501 downto 8496 );
    VN1417_data_out <= VN_data_out( 8507 downto 8502 );
    VN1417_sign_out <= VN_sign_out( 8507 downto 8502 );
    VN1418_data_out <= VN_data_out( 8513 downto 8508 );
    VN1418_sign_out <= VN_sign_out( 8513 downto 8508 );
    VN1419_data_out <= VN_data_out( 8519 downto 8514 );
    VN1419_sign_out <= VN_sign_out( 8519 downto 8514 );
    VN1420_data_out <= VN_data_out( 8525 downto 8520 );
    VN1420_sign_out <= VN_sign_out( 8525 downto 8520 );
    VN1421_data_out <= VN_data_out( 8531 downto 8526 );
    VN1421_sign_out <= VN_sign_out( 8531 downto 8526 );
    VN1422_data_out <= VN_data_out( 8537 downto 8532 );
    VN1422_sign_out <= VN_sign_out( 8537 downto 8532 );
    VN1423_data_out <= VN_data_out( 8543 downto 8538 );
    VN1423_sign_out <= VN_sign_out( 8543 downto 8538 );
    VN1424_data_out <= VN_data_out( 8549 downto 8544 );
    VN1424_sign_out <= VN_sign_out( 8549 downto 8544 );
    VN1425_data_out <= VN_data_out( 8555 downto 8550 );
    VN1425_sign_out <= VN_sign_out( 8555 downto 8550 );
    VN1426_data_out <= VN_data_out( 8561 downto 8556 );
    VN1426_sign_out <= VN_sign_out( 8561 downto 8556 );
    VN1427_data_out <= VN_data_out( 8567 downto 8562 );
    VN1427_sign_out <= VN_sign_out( 8567 downto 8562 );
    VN1428_data_out <= VN_data_out( 8573 downto 8568 );
    VN1428_sign_out <= VN_sign_out( 8573 downto 8568 );
    VN1429_data_out <= VN_data_out( 8579 downto 8574 );
    VN1429_sign_out <= VN_sign_out( 8579 downto 8574 );
    VN1430_data_out <= VN_data_out( 8585 downto 8580 );
    VN1430_sign_out <= VN_sign_out( 8585 downto 8580 );
    VN1431_data_out <= VN_data_out( 8591 downto 8586 );
    VN1431_sign_out <= VN_sign_out( 8591 downto 8586 );
    VN1432_data_out <= VN_data_out( 8597 downto 8592 );
    VN1432_sign_out <= VN_sign_out( 8597 downto 8592 );
    VN1433_data_out <= VN_data_out( 8603 downto 8598 );
    VN1433_sign_out <= VN_sign_out( 8603 downto 8598 );
    VN1434_data_out <= VN_data_out( 8609 downto 8604 );
    VN1434_sign_out <= VN_sign_out( 8609 downto 8604 );
    VN1435_data_out <= VN_data_out( 8615 downto 8610 );
    VN1435_sign_out <= VN_sign_out( 8615 downto 8610 );
    VN1436_data_out <= VN_data_out( 8621 downto 8616 );
    VN1436_sign_out <= VN_sign_out( 8621 downto 8616 );
    VN1437_data_out <= VN_data_out( 8627 downto 8622 );
    VN1437_sign_out <= VN_sign_out( 8627 downto 8622 );
    VN1438_data_out <= VN_data_out( 8633 downto 8628 );
    VN1438_sign_out <= VN_sign_out( 8633 downto 8628 );
    VN1439_data_out <= VN_data_out( 8639 downto 8634 );
    VN1439_sign_out <= VN_sign_out( 8639 downto 8634 );
    VN1440_data_out <= VN_data_out( 8645 downto 8640 );
    VN1440_sign_out <= VN_sign_out( 8645 downto 8640 );
    VN1441_data_out <= VN_data_out( 8651 downto 8646 );
    VN1441_sign_out <= VN_sign_out( 8651 downto 8646 );
    VN1442_data_out <= VN_data_out( 8657 downto 8652 );
    VN1442_sign_out <= VN_sign_out( 8657 downto 8652 );
    VN1443_data_out <= VN_data_out( 8663 downto 8658 );
    VN1443_sign_out <= VN_sign_out( 8663 downto 8658 );
    VN1444_data_out <= VN_data_out( 8669 downto 8664 );
    VN1444_sign_out <= VN_sign_out( 8669 downto 8664 );
    VN1445_data_out <= VN_data_out( 8675 downto 8670 );
    VN1445_sign_out <= VN_sign_out( 8675 downto 8670 );
    VN1446_data_out <= VN_data_out( 8681 downto 8676 );
    VN1446_sign_out <= VN_sign_out( 8681 downto 8676 );
    VN1447_data_out <= VN_data_out( 8687 downto 8682 );
    VN1447_sign_out <= VN_sign_out( 8687 downto 8682 );
    VN1448_data_out <= VN_data_out( 8693 downto 8688 );
    VN1448_sign_out <= VN_sign_out( 8693 downto 8688 );
    VN1449_data_out <= VN_data_out( 8699 downto 8694 );
    VN1449_sign_out <= VN_sign_out( 8699 downto 8694 );
    VN1450_data_out <= VN_data_out( 8705 downto 8700 );
    VN1450_sign_out <= VN_sign_out( 8705 downto 8700 );
    VN1451_data_out <= VN_data_out( 8711 downto 8706 );
    VN1451_sign_out <= VN_sign_out( 8711 downto 8706 );
    VN1452_data_out <= VN_data_out( 8717 downto 8712 );
    VN1452_sign_out <= VN_sign_out( 8717 downto 8712 );
    VN1453_data_out <= VN_data_out( 8723 downto 8718 );
    VN1453_sign_out <= VN_sign_out( 8723 downto 8718 );
    VN1454_data_out <= VN_data_out( 8729 downto 8724 );
    VN1454_sign_out <= VN_sign_out( 8729 downto 8724 );
    VN1455_data_out <= VN_data_out( 8735 downto 8730 );
    VN1455_sign_out <= VN_sign_out( 8735 downto 8730 );
    VN1456_data_out <= VN_data_out( 8741 downto 8736 );
    VN1456_sign_out <= VN_sign_out( 8741 downto 8736 );
    VN1457_data_out <= VN_data_out( 8747 downto 8742 );
    VN1457_sign_out <= VN_sign_out( 8747 downto 8742 );
    VN1458_data_out <= VN_data_out( 8753 downto 8748 );
    VN1458_sign_out <= VN_sign_out( 8753 downto 8748 );
    VN1459_data_out <= VN_data_out( 8759 downto 8754 );
    VN1459_sign_out <= VN_sign_out( 8759 downto 8754 );
    VN1460_data_out <= VN_data_out( 8765 downto 8760 );
    VN1460_sign_out <= VN_sign_out( 8765 downto 8760 );
    VN1461_data_out <= VN_data_out( 8771 downto 8766 );
    VN1461_sign_out <= VN_sign_out( 8771 downto 8766 );
    VN1462_data_out <= VN_data_out( 8777 downto 8772 );
    VN1462_sign_out <= VN_sign_out( 8777 downto 8772 );
    VN1463_data_out <= VN_data_out( 8783 downto 8778 );
    VN1463_sign_out <= VN_sign_out( 8783 downto 8778 );
    VN1464_data_out <= VN_data_out( 8789 downto 8784 );
    VN1464_sign_out <= VN_sign_out( 8789 downto 8784 );
    VN1465_data_out <= VN_data_out( 8795 downto 8790 );
    VN1465_sign_out <= VN_sign_out( 8795 downto 8790 );
    VN1466_data_out <= VN_data_out( 8801 downto 8796 );
    VN1466_sign_out <= VN_sign_out( 8801 downto 8796 );
    VN1467_data_out <= VN_data_out( 8807 downto 8802 );
    VN1467_sign_out <= VN_sign_out( 8807 downto 8802 );
    VN1468_data_out <= VN_data_out( 8813 downto 8808 );
    VN1468_sign_out <= VN_sign_out( 8813 downto 8808 );
    VN1469_data_out <= VN_data_out( 8819 downto 8814 );
    VN1469_sign_out <= VN_sign_out( 8819 downto 8814 );
    VN1470_data_out <= VN_data_out( 8825 downto 8820 );
    VN1470_sign_out <= VN_sign_out( 8825 downto 8820 );
    VN1471_data_out <= VN_data_out( 8831 downto 8826 );
    VN1471_sign_out <= VN_sign_out( 8831 downto 8826 );
    VN1472_data_out <= VN_data_out( 8837 downto 8832 );
    VN1472_sign_out <= VN_sign_out( 8837 downto 8832 );
    VN1473_data_out <= VN_data_out( 8843 downto 8838 );
    VN1473_sign_out <= VN_sign_out( 8843 downto 8838 );
    VN1474_data_out <= VN_data_out( 8849 downto 8844 );
    VN1474_sign_out <= VN_sign_out( 8849 downto 8844 );
    VN1475_data_out <= VN_data_out( 8855 downto 8850 );
    VN1475_sign_out <= VN_sign_out( 8855 downto 8850 );
    VN1476_data_out <= VN_data_out( 8861 downto 8856 );
    VN1476_sign_out <= VN_sign_out( 8861 downto 8856 );
    VN1477_data_out <= VN_data_out( 8867 downto 8862 );
    VN1477_sign_out <= VN_sign_out( 8867 downto 8862 );
    VN1478_data_out <= VN_data_out( 8873 downto 8868 );
    VN1478_sign_out <= VN_sign_out( 8873 downto 8868 );
    VN1479_data_out <= VN_data_out( 8879 downto 8874 );
    VN1479_sign_out <= VN_sign_out( 8879 downto 8874 );
    VN1480_data_out <= VN_data_out( 8885 downto 8880 );
    VN1480_sign_out <= VN_sign_out( 8885 downto 8880 );
    VN1481_data_out <= VN_data_out( 8891 downto 8886 );
    VN1481_sign_out <= VN_sign_out( 8891 downto 8886 );
    VN1482_data_out <= VN_data_out( 8897 downto 8892 );
    VN1482_sign_out <= VN_sign_out( 8897 downto 8892 );
    VN1483_data_out <= VN_data_out( 8903 downto 8898 );
    VN1483_sign_out <= VN_sign_out( 8903 downto 8898 );
    VN1484_data_out <= VN_data_out( 8909 downto 8904 );
    VN1484_sign_out <= VN_sign_out( 8909 downto 8904 );
    VN1485_data_out <= VN_data_out( 8915 downto 8910 );
    VN1485_sign_out <= VN_sign_out( 8915 downto 8910 );
    VN1486_data_out <= VN_data_out( 8921 downto 8916 );
    VN1486_sign_out <= VN_sign_out( 8921 downto 8916 );
    VN1487_data_out <= VN_data_out( 8927 downto 8922 );
    VN1487_sign_out <= VN_sign_out( 8927 downto 8922 );
    VN1488_data_out <= VN_data_out( 8933 downto 8928 );
    VN1488_sign_out <= VN_sign_out( 8933 downto 8928 );
    VN1489_data_out <= VN_data_out( 8939 downto 8934 );
    VN1489_sign_out <= VN_sign_out( 8939 downto 8934 );
    VN1490_data_out <= VN_data_out( 8945 downto 8940 );
    VN1490_sign_out <= VN_sign_out( 8945 downto 8940 );
    VN1491_data_out <= VN_data_out( 8951 downto 8946 );
    VN1491_sign_out <= VN_sign_out( 8951 downto 8946 );
    VN1492_data_out <= VN_data_out( 8957 downto 8952 );
    VN1492_sign_out <= VN_sign_out( 8957 downto 8952 );
    VN1493_data_out <= VN_data_out( 8963 downto 8958 );
    VN1493_sign_out <= VN_sign_out( 8963 downto 8958 );
    VN1494_data_out <= VN_data_out( 8969 downto 8964 );
    VN1494_sign_out <= VN_sign_out( 8969 downto 8964 );
    VN1495_data_out <= VN_data_out( 8975 downto 8970 );
    VN1495_sign_out <= VN_sign_out( 8975 downto 8970 );
    VN1496_data_out <= VN_data_out( 8981 downto 8976 );
    VN1496_sign_out <= VN_sign_out( 8981 downto 8976 );
    VN1497_data_out <= VN_data_out( 8987 downto 8982 );
    VN1497_sign_out <= VN_sign_out( 8987 downto 8982 );
    VN1498_data_out <= VN_data_out( 8993 downto 8988 );
    VN1498_sign_out <= VN_sign_out( 8993 downto 8988 );
    VN1499_data_out <= VN_data_out( 8999 downto 8994 );
    VN1499_sign_out <= VN_sign_out( 8999 downto 8994 );
    VN1500_data_out <= VN_data_out( 9005 downto 9000 );
    VN1500_sign_out <= VN_sign_out( 9005 downto 9000 );
    VN1501_data_out <= VN_data_out( 9011 downto 9006 );
    VN1501_sign_out <= VN_sign_out( 9011 downto 9006 );
    VN1502_data_out <= VN_data_out( 9017 downto 9012 );
    VN1502_sign_out <= VN_sign_out( 9017 downto 9012 );
    VN1503_data_out <= VN_data_out( 9023 downto 9018 );
    VN1503_sign_out <= VN_sign_out( 9023 downto 9018 );
    VN1504_data_out <= VN_data_out( 9029 downto 9024 );
    VN1504_sign_out <= VN_sign_out( 9029 downto 9024 );
    VN1505_data_out <= VN_data_out( 9035 downto 9030 );
    VN1505_sign_out <= VN_sign_out( 9035 downto 9030 );
    VN1506_data_out <= VN_data_out( 9041 downto 9036 );
    VN1506_sign_out <= VN_sign_out( 9041 downto 9036 );
    VN1507_data_out <= VN_data_out( 9047 downto 9042 );
    VN1507_sign_out <= VN_sign_out( 9047 downto 9042 );
    VN1508_data_out <= VN_data_out( 9053 downto 9048 );
    VN1508_sign_out <= VN_sign_out( 9053 downto 9048 );
    VN1509_data_out <= VN_data_out( 9059 downto 9054 );
    VN1509_sign_out <= VN_sign_out( 9059 downto 9054 );
    VN1510_data_out <= VN_data_out( 9065 downto 9060 );
    VN1510_sign_out <= VN_sign_out( 9065 downto 9060 );
    VN1511_data_out <= VN_data_out( 9071 downto 9066 );
    VN1511_sign_out <= VN_sign_out( 9071 downto 9066 );
    VN1512_data_out <= VN_data_out( 9077 downto 9072 );
    VN1512_sign_out <= VN_sign_out( 9077 downto 9072 );
    VN1513_data_out <= VN_data_out( 9083 downto 9078 );
    VN1513_sign_out <= VN_sign_out( 9083 downto 9078 );
    VN1514_data_out <= VN_data_out( 9089 downto 9084 );
    VN1514_sign_out <= VN_sign_out( 9089 downto 9084 );
    VN1515_data_out <= VN_data_out( 9095 downto 9090 );
    VN1515_sign_out <= VN_sign_out( 9095 downto 9090 );
    VN1516_data_out <= VN_data_out( 9101 downto 9096 );
    VN1516_sign_out <= VN_sign_out( 9101 downto 9096 );
    VN1517_data_out <= VN_data_out( 9107 downto 9102 );
    VN1517_sign_out <= VN_sign_out( 9107 downto 9102 );
    VN1518_data_out <= VN_data_out( 9113 downto 9108 );
    VN1518_sign_out <= VN_sign_out( 9113 downto 9108 );
    VN1519_data_out <= VN_data_out( 9119 downto 9114 );
    VN1519_sign_out <= VN_sign_out( 9119 downto 9114 );
    VN1520_data_out <= VN_data_out( 9125 downto 9120 );
    VN1520_sign_out <= VN_sign_out( 9125 downto 9120 );
    VN1521_data_out <= VN_data_out( 9131 downto 9126 );
    VN1521_sign_out <= VN_sign_out( 9131 downto 9126 );
    VN1522_data_out <= VN_data_out( 9137 downto 9132 );
    VN1522_sign_out <= VN_sign_out( 9137 downto 9132 );
    VN1523_data_out <= VN_data_out( 9143 downto 9138 );
    VN1523_sign_out <= VN_sign_out( 9143 downto 9138 );
    VN1524_data_out <= VN_data_out( 9149 downto 9144 );
    VN1524_sign_out <= VN_sign_out( 9149 downto 9144 );
    VN1525_data_out <= VN_data_out( 9155 downto 9150 );
    VN1525_sign_out <= VN_sign_out( 9155 downto 9150 );
    VN1526_data_out <= VN_data_out( 9161 downto 9156 );
    VN1526_sign_out <= VN_sign_out( 9161 downto 9156 );
    VN1527_data_out <= VN_data_out( 9167 downto 9162 );
    VN1527_sign_out <= VN_sign_out( 9167 downto 9162 );
    VN1528_data_out <= VN_data_out( 9173 downto 9168 );
    VN1528_sign_out <= VN_sign_out( 9173 downto 9168 );
    VN1529_data_out <= VN_data_out( 9179 downto 9174 );
    VN1529_sign_out <= VN_sign_out( 9179 downto 9174 );
    VN1530_data_out <= VN_data_out( 9185 downto 9180 );
    VN1530_sign_out <= VN_sign_out( 9185 downto 9180 );
    VN1531_data_out <= VN_data_out( 9191 downto 9186 );
    VN1531_sign_out <= VN_sign_out( 9191 downto 9186 );
    VN1532_data_out <= VN_data_out( 9197 downto 9192 );
    VN1532_sign_out <= VN_sign_out( 9197 downto 9192 );
    VN1533_data_out <= VN_data_out( 9203 downto 9198 );
    VN1533_sign_out <= VN_sign_out( 9203 downto 9198 );
    VN1534_data_out <= VN_data_out( 9209 downto 9204 );
    VN1534_sign_out <= VN_sign_out( 9209 downto 9204 );
    VN1535_data_out <= VN_data_out( 9215 downto 9210 );
    VN1535_sign_out <= VN_sign_out( 9215 downto 9210 );
    VN1536_data_out <= VN_data_out( 9221 downto 9216 );
    VN1536_sign_out <= VN_sign_out( 9221 downto 9216 );
    VN1537_data_out <= VN_data_out( 9227 downto 9222 );
    VN1537_sign_out <= VN_sign_out( 9227 downto 9222 );
    VN1538_data_out <= VN_data_out( 9233 downto 9228 );
    VN1538_sign_out <= VN_sign_out( 9233 downto 9228 );
    VN1539_data_out <= VN_data_out( 9239 downto 9234 );
    VN1539_sign_out <= VN_sign_out( 9239 downto 9234 );
    VN1540_data_out <= VN_data_out( 9245 downto 9240 );
    VN1540_sign_out <= VN_sign_out( 9245 downto 9240 );
    VN1541_data_out <= VN_data_out( 9251 downto 9246 );
    VN1541_sign_out <= VN_sign_out( 9251 downto 9246 );
    VN1542_data_out <= VN_data_out( 9257 downto 9252 );
    VN1542_sign_out <= VN_sign_out( 9257 downto 9252 );
    VN1543_data_out <= VN_data_out( 9263 downto 9258 );
    VN1543_sign_out <= VN_sign_out( 9263 downto 9258 );
    VN1544_data_out <= VN_data_out( 9269 downto 9264 );
    VN1544_sign_out <= VN_sign_out( 9269 downto 9264 );
    VN1545_data_out <= VN_data_out( 9275 downto 9270 );
    VN1545_sign_out <= VN_sign_out( 9275 downto 9270 );
    VN1546_data_out <= VN_data_out( 9281 downto 9276 );
    VN1546_sign_out <= VN_sign_out( 9281 downto 9276 );
    VN1547_data_out <= VN_data_out( 9287 downto 9282 );
    VN1547_sign_out <= VN_sign_out( 9287 downto 9282 );
    VN1548_data_out <= VN_data_out( 9293 downto 9288 );
    VN1548_sign_out <= VN_sign_out( 9293 downto 9288 );
    VN1549_data_out <= VN_data_out( 9299 downto 9294 );
    VN1549_sign_out <= VN_sign_out( 9299 downto 9294 );
    VN1550_data_out <= VN_data_out( 9305 downto 9300 );
    VN1550_sign_out <= VN_sign_out( 9305 downto 9300 );
    VN1551_data_out <= VN_data_out( 9311 downto 9306 );
    VN1551_sign_out <= VN_sign_out( 9311 downto 9306 );
    VN1552_data_out <= VN_data_out( 9317 downto 9312 );
    VN1552_sign_out <= VN_sign_out( 9317 downto 9312 );
    VN1553_data_out <= VN_data_out( 9323 downto 9318 );
    VN1553_sign_out <= VN_sign_out( 9323 downto 9318 );
    VN1554_data_out <= VN_data_out( 9329 downto 9324 );
    VN1554_sign_out <= VN_sign_out( 9329 downto 9324 );
    VN1555_data_out <= VN_data_out( 9335 downto 9330 );
    VN1555_sign_out <= VN_sign_out( 9335 downto 9330 );
    VN1556_data_out <= VN_data_out( 9341 downto 9336 );
    VN1556_sign_out <= VN_sign_out( 9341 downto 9336 );
    VN1557_data_out <= VN_data_out( 9347 downto 9342 );
    VN1557_sign_out <= VN_sign_out( 9347 downto 9342 );
    VN1558_data_out <= VN_data_out( 9353 downto 9348 );
    VN1558_sign_out <= VN_sign_out( 9353 downto 9348 );
    VN1559_data_out <= VN_data_out( 9359 downto 9354 );
    VN1559_sign_out <= VN_sign_out( 9359 downto 9354 );
    VN1560_data_out <= VN_data_out( 9365 downto 9360 );
    VN1560_sign_out <= VN_sign_out( 9365 downto 9360 );
    VN1561_data_out <= VN_data_out( 9371 downto 9366 );
    VN1561_sign_out <= VN_sign_out( 9371 downto 9366 );
    VN1562_data_out <= VN_data_out( 9377 downto 9372 );
    VN1562_sign_out <= VN_sign_out( 9377 downto 9372 );
    VN1563_data_out <= VN_data_out( 9383 downto 9378 );
    VN1563_sign_out <= VN_sign_out( 9383 downto 9378 );
    VN1564_data_out <= VN_data_out( 9389 downto 9384 );
    VN1564_sign_out <= VN_sign_out( 9389 downto 9384 );
    VN1565_data_out <= VN_data_out( 9395 downto 9390 );
    VN1565_sign_out <= VN_sign_out( 9395 downto 9390 );
    VN1566_data_out <= VN_data_out( 9401 downto 9396 );
    VN1566_sign_out <= VN_sign_out( 9401 downto 9396 );
    VN1567_data_out <= VN_data_out( 9407 downto 9402 );
    VN1567_sign_out <= VN_sign_out( 9407 downto 9402 );
    VN1568_data_out <= VN_data_out( 9413 downto 9408 );
    VN1568_sign_out <= VN_sign_out( 9413 downto 9408 );
    VN1569_data_out <= VN_data_out( 9419 downto 9414 );
    VN1569_sign_out <= VN_sign_out( 9419 downto 9414 );
    VN1570_data_out <= VN_data_out( 9425 downto 9420 );
    VN1570_sign_out <= VN_sign_out( 9425 downto 9420 );
    VN1571_data_out <= VN_data_out( 9431 downto 9426 );
    VN1571_sign_out <= VN_sign_out( 9431 downto 9426 );
    VN1572_data_out <= VN_data_out( 9437 downto 9432 );
    VN1572_sign_out <= VN_sign_out( 9437 downto 9432 );
    VN1573_data_out <= VN_data_out( 9443 downto 9438 );
    VN1573_sign_out <= VN_sign_out( 9443 downto 9438 );
    VN1574_data_out <= VN_data_out( 9449 downto 9444 );
    VN1574_sign_out <= VN_sign_out( 9449 downto 9444 );
    VN1575_data_out <= VN_data_out( 9455 downto 9450 );
    VN1575_sign_out <= VN_sign_out( 9455 downto 9450 );
    VN1576_data_out <= VN_data_out( 9461 downto 9456 );
    VN1576_sign_out <= VN_sign_out( 9461 downto 9456 );
    VN1577_data_out <= VN_data_out( 9467 downto 9462 );
    VN1577_sign_out <= VN_sign_out( 9467 downto 9462 );
    VN1578_data_out <= VN_data_out( 9473 downto 9468 );
    VN1578_sign_out <= VN_sign_out( 9473 downto 9468 );
    VN1579_data_out <= VN_data_out( 9479 downto 9474 );
    VN1579_sign_out <= VN_sign_out( 9479 downto 9474 );
    VN1580_data_out <= VN_data_out( 9485 downto 9480 );
    VN1580_sign_out <= VN_sign_out( 9485 downto 9480 );
    VN1581_data_out <= VN_data_out( 9491 downto 9486 );
    VN1581_sign_out <= VN_sign_out( 9491 downto 9486 );
    VN1582_data_out <= VN_data_out( 9497 downto 9492 );
    VN1582_sign_out <= VN_sign_out( 9497 downto 9492 );
    VN1583_data_out <= VN_data_out( 9503 downto 9498 );
    VN1583_sign_out <= VN_sign_out( 9503 downto 9498 );
    VN1584_data_out <= VN_data_out( 9509 downto 9504 );
    VN1584_sign_out <= VN_sign_out( 9509 downto 9504 );
    VN1585_data_out <= VN_data_out( 9515 downto 9510 );
    VN1585_sign_out <= VN_sign_out( 9515 downto 9510 );
    VN1586_data_out <= VN_data_out( 9521 downto 9516 );
    VN1586_sign_out <= VN_sign_out( 9521 downto 9516 );
    VN1587_data_out <= VN_data_out( 9527 downto 9522 );
    VN1587_sign_out <= VN_sign_out( 9527 downto 9522 );
    VN1588_data_out <= VN_data_out( 9533 downto 9528 );
    VN1588_sign_out <= VN_sign_out( 9533 downto 9528 );
    VN1589_data_out <= VN_data_out( 9539 downto 9534 );
    VN1589_sign_out <= VN_sign_out( 9539 downto 9534 );
    VN1590_data_out <= VN_data_out( 9545 downto 9540 );
    VN1590_sign_out <= VN_sign_out( 9545 downto 9540 );
    VN1591_data_out <= VN_data_out( 9551 downto 9546 );
    VN1591_sign_out <= VN_sign_out( 9551 downto 9546 );
    VN1592_data_out <= VN_data_out( 9557 downto 9552 );
    VN1592_sign_out <= VN_sign_out( 9557 downto 9552 );
    VN1593_data_out <= VN_data_out( 9563 downto 9558 );
    VN1593_sign_out <= VN_sign_out( 9563 downto 9558 );
    VN1594_data_out <= VN_data_out( 9569 downto 9564 );
    VN1594_sign_out <= VN_sign_out( 9569 downto 9564 );
    VN1595_data_out <= VN_data_out( 9575 downto 9570 );
    VN1595_sign_out <= VN_sign_out( 9575 downto 9570 );
    VN1596_data_out <= VN_data_out( 9581 downto 9576 );
    VN1596_sign_out <= VN_sign_out( 9581 downto 9576 );
    VN1597_data_out <= VN_data_out( 9587 downto 9582 );
    VN1597_sign_out <= VN_sign_out( 9587 downto 9582 );
    VN1598_data_out <= VN_data_out( 9593 downto 9588 );
    VN1598_sign_out <= VN_sign_out( 9593 downto 9588 );
    VN1599_data_out <= VN_data_out( 9599 downto 9594 );
    VN1599_sign_out <= VN_sign_out( 9599 downto 9594 );
    VN1600_data_out <= VN_data_out( 9605 downto 9600 );
    VN1600_sign_out <= VN_sign_out( 9605 downto 9600 );
    VN1601_data_out <= VN_data_out( 9611 downto 9606 );
    VN1601_sign_out <= VN_sign_out( 9611 downto 9606 );
    VN1602_data_out <= VN_data_out( 9617 downto 9612 );
    VN1602_sign_out <= VN_sign_out( 9617 downto 9612 );
    VN1603_data_out <= VN_data_out( 9623 downto 9618 );
    VN1603_sign_out <= VN_sign_out( 9623 downto 9618 );
    VN1604_data_out <= VN_data_out( 9629 downto 9624 );
    VN1604_sign_out <= VN_sign_out( 9629 downto 9624 );
    VN1605_data_out <= VN_data_out( 9635 downto 9630 );
    VN1605_sign_out <= VN_sign_out( 9635 downto 9630 );
    VN1606_data_out <= VN_data_out( 9641 downto 9636 );
    VN1606_sign_out <= VN_sign_out( 9641 downto 9636 );
    VN1607_data_out <= VN_data_out( 9647 downto 9642 );
    VN1607_sign_out <= VN_sign_out( 9647 downto 9642 );
    VN1608_data_out <= VN_data_out( 9653 downto 9648 );
    VN1608_sign_out <= VN_sign_out( 9653 downto 9648 );
    VN1609_data_out <= VN_data_out( 9659 downto 9654 );
    VN1609_sign_out <= VN_sign_out( 9659 downto 9654 );
    VN1610_data_out <= VN_data_out( 9665 downto 9660 );
    VN1610_sign_out <= VN_sign_out( 9665 downto 9660 );
    VN1611_data_out <= VN_data_out( 9671 downto 9666 );
    VN1611_sign_out <= VN_sign_out( 9671 downto 9666 );
    VN1612_data_out <= VN_data_out( 9677 downto 9672 );
    VN1612_sign_out <= VN_sign_out( 9677 downto 9672 );
    VN1613_data_out <= VN_data_out( 9683 downto 9678 );
    VN1613_sign_out <= VN_sign_out( 9683 downto 9678 );
    VN1614_data_out <= VN_data_out( 9689 downto 9684 );
    VN1614_sign_out <= VN_sign_out( 9689 downto 9684 );
    VN1615_data_out <= VN_data_out( 9695 downto 9690 );
    VN1615_sign_out <= VN_sign_out( 9695 downto 9690 );
    VN1616_data_out <= VN_data_out( 9701 downto 9696 );
    VN1616_sign_out <= VN_sign_out( 9701 downto 9696 );
    VN1617_data_out <= VN_data_out( 9707 downto 9702 );
    VN1617_sign_out <= VN_sign_out( 9707 downto 9702 );
    VN1618_data_out <= VN_data_out( 9713 downto 9708 );
    VN1618_sign_out <= VN_sign_out( 9713 downto 9708 );
    VN1619_data_out <= VN_data_out( 9719 downto 9714 );
    VN1619_sign_out <= VN_sign_out( 9719 downto 9714 );
    VN1620_data_out <= VN_data_out( 9725 downto 9720 );
    VN1620_sign_out <= VN_sign_out( 9725 downto 9720 );
    VN1621_data_out <= VN_data_out( 9731 downto 9726 );
    VN1621_sign_out <= VN_sign_out( 9731 downto 9726 );
    VN1622_data_out <= VN_data_out( 9737 downto 9732 );
    VN1622_sign_out <= VN_sign_out( 9737 downto 9732 );
    VN1623_data_out <= VN_data_out( 9743 downto 9738 );
    VN1623_sign_out <= VN_sign_out( 9743 downto 9738 );
    VN1624_data_out <= VN_data_out( 9749 downto 9744 );
    VN1624_sign_out <= VN_sign_out( 9749 downto 9744 );
    VN1625_data_out <= VN_data_out( 9755 downto 9750 );
    VN1625_sign_out <= VN_sign_out( 9755 downto 9750 );
    VN1626_data_out <= VN_data_out( 9761 downto 9756 );
    VN1626_sign_out <= VN_sign_out( 9761 downto 9756 );
    VN1627_data_out <= VN_data_out( 9767 downto 9762 );
    VN1627_sign_out <= VN_sign_out( 9767 downto 9762 );
    VN1628_data_out <= VN_data_out( 9773 downto 9768 );
    VN1628_sign_out <= VN_sign_out( 9773 downto 9768 );
    VN1629_data_out <= VN_data_out( 9779 downto 9774 );
    VN1629_sign_out <= VN_sign_out( 9779 downto 9774 );
    VN1630_data_out <= VN_data_out( 9785 downto 9780 );
    VN1630_sign_out <= VN_sign_out( 9785 downto 9780 );
    VN1631_data_out <= VN_data_out( 9791 downto 9786 );
    VN1631_sign_out <= VN_sign_out( 9791 downto 9786 );
    VN1632_data_out <= VN_data_out( 9797 downto 9792 );
    VN1632_sign_out <= VN_sign_out( 9797 downto 9792 );
    VN1633_data_out <= VN_data_out( 9803 downto 9798 );
    VN1633_sign_out <= VN_sign_out( 9803 downto 9798 );
    VN1634_data_out <= VN_data_out( 9809 downto 9804 );
    VN1634_sign_out <= VN_sign_out( 9809 downto 9804 );
    VN1635_data_out <= VN_data_out( 9815 downto 9810 );
    VN1635_sign_out <= VN_sign_out( 9815 downto 9810 );
    VN1636_data_out <= VN_data_out( 9821 downto 9816 );
    VN1636_sign_out <= VN_sign_out( 9821 downto 9816 );
    VN1637_data_out <= VN_data_out( 9827 downto 9822 );
    VN1637_sign_out <= VN_sign_out( 9827 downto 9822 );
    VN1638_data_out <= VN_data_out( 9833 downto 9828 );
    VN1638_sign_out <= VN_sign_out( 9833 downto 9828 );
    VN1639_data_out <= VN_data_out( 9839 downto 9834 );
    VN1639_sign_out <= VN_sign_out( 9839 downto 9834 );
    VN1640_data_out <= VN_data_out( 9845 downto 9840 );
    VN1640_sign_out <= VN_sign_out( 9845 downto 9840 );
    VN1641_data_out <= VN_data_out( 9851 downto 9846 );
    VN1641_sign_out <= VN_sign_out( 9851 downto 9846 );
    VN1642_data_out <= VN_data_out( 9857 downto 9852 );
    VN1642_sign_out <= VN_sign_out( 9857 downto 9852 );
    VN1643_data_out <= VN_data_out( 9863 downto 9858 );
    VN1643_sign_out <= VN_sign_out( 9863 downto 9858 );
    VN1644_data_out <= VN_data_out( 9869 downto 9864 );
    VN1644_sign_out <= VN_sign_out( 9869 downto 9864 );
    VN1645_data_out <= VN_data_out( 9875 downto 9870 );
    VN1645_sign_out <= VN_sign_out( 9875 downto 9870 );
    VN1646_data_out <= VN_data_out( 9881 downto 9876 );
    VN1646_sign_out <= VN_sign_out( 9881 downto 9876 );
    VN1647_data_out <= VN_data_out( 9887 downto 9882 );
    VN1647_sign_out <= VN_sign_out( 9887 downto 9882 );
    VN1648_data_out <= VN_data_out( 9893 downto 9888 );
    VN1648_sign_out <= VN_sign_out( 9893 downto 9888 );
    VN1649_data_out <= VN_data_out( 9899 downto 9894 );
    VN1649_sign_out <= VN_sign_out( 9899 downto 9894 );
    VN1650_data_out <= VN_data_out( 9905 downto 9900 );
    VN1650_sign_out <= VN_sign_out( 9905 downto 9900 );
    VN1651_data_out <= VN_data_out( 9911 downto 9906 );
    VN1651_sign_out <= VN_sign_out( 9911 downto 9906 );
    VN1652_data_out <= VN_data_out( 9917 downto 9912 );
    VN1652_sign_out <= VN_sign_out( 9917 downto 9912 );
    VN1653_data_out <= VN_data_out( 9923 downto 9918 );
    VN1653_sign_out <= VN_sign_out( 9923 downto 9918 );
    VN1654_data_out <= VN_data_out( 9929 downto 9924 );
    VN1654_sign_out <= VN_sign_out( 9929 downto 9924 );
    VN1655_data_out <= VN_data_out( 9935 downto 9930 );
    VN1655_sign_out <= VN_sign_out( 9935 downto 9930 );
    VN1656_data_out <= VN_data_out( 9941 downto 9936 );
    VN1656_sign_out <= VN_sign_out( 9941 downto 9936 );
    VN1657_data_out <= VN_data_out( 9947 downto 9942 );
    VN1657_sign_out <= VN_sign_out( 9947 downto 9942 );
    VN1658_data_out <= VN_data_out( 9953 downto 9948 );
    VN1658_sign_out <= VN_sign_out( 9953 downto 9948 );
    VN1659_data_out <= VN_data_out( 9959 downto 9954 );
    VN1659_sign_out <= VN_sign_out( 9959 downto 9954 );
    VN1660_data_out <= VN_data_out( 9965 downto 9960 );
    VN1660_sign_out <= VN_sign_out( 9965 downto 9960 );
    VN1661_data_out <= VN_data_out( 9971 downto 9966 );
    VN1661_sign_out <= VN_sign_out( 9971 downto 9966 );
    VN1662_data_out <= VN_data_out( 9977 downto 9972 );
    VN1662_sign_out <= VN_sign_out( 9977 downto 9972 );
    VN1663_data_out <= VN_data_out( 9983 downto 9978 );
    VN1663_sign_out <= VN_sign_out( 9983 downto 9978 );
    VN1664_data_out <= VN_data_out( 9989 downto 9984 );
    VN1664_sign_out <= VN_sign_out( 9989 downto 9984 );
    VN1665_data_out <= VN_data_out( 9995 downto 9990 );
    VN1665_sign_out <= VN_sign_out( 9995 downto 9990 );
    VN1666_data_out <= VN_data_out( 10001 downto 9996 );
    VN1666_sign_out <= VN_sign_out( 10001 downto 9996 );
    VN1667_data_out <= VN_data_out( 10007 downto 10002 );
    VN1667_sign_out <= VN_sign_out( 10007 downto 10002 );
    VN1668_data_out <= VN_data_out( 10013 downto 10008 );
    VN1668_sign_out <= VN_sign_out( 10013 downto 10008 );
    VN1669_data_out <= VN_data_out( 10019 downto 10014 );
    VN1669_sign_out <= VN_sign_out( 10019 downto 10014 );
    VN1670_data_out <= VN_data_out( 10025 downto 10020 );
    VN1670_sign_out <= VN_sign_out( 10025 downto 10020 );
    VN1671_data_out <= VN_data_out( 10031 downto 10026 );
    VN1671_sign_out <= VN_sign_out( 10031 downto 10026 );
    VN1672_data_out <= VN_data_out( 10037 downto 10032 );
    VN1672_sign_out <= VN_sign_out( 10037 downto 10032 );
    VN1673_data_out <= VN_data_out( 10043 downto 10038 );
    VN1673_sign_out <= VN_sign_out( 10043 downto 10038 );
    VN1674_data_out <= VN_data_out( 10049 downto 10044 );
    VN1674_sign_out <= VN_sign_out( 10049 downto 10044 );
    VN1675_data_out <= VN_data_out( 10055 downto 10050 );
    VN1675_sign_out <= VN_sign_out( 10055 downto 10050 );
    VN1676_data_out <= VN_data_out( 10061 downto 10056 );
    VN1676_sign_out <= VN_sign_out( 10061 downto 10056 );
    VN1677_data_out <= VN_data_out( 10067 downto 10062 );
    VN1677_sign_out <= VN_sign_out( 10067 downto 10062 );
    VN1678_data_out <= VN_data_out( 10073 downto 10068 );
    VN1678_sign_out <= VN_sign_out( 10073 downto 10068 );
    VN1679_data_out <= VN_data_out( 10079 downto 10074 );
    VN1679_sign_out <= VN_sign_out( 10079 downto 10074 );
    VN1680_data_out <= VN_data_out( 10085 downto 10080 );
    VN1680_sign_out <= VN_sign_out( 10085 downto 10080 );
    VN1681_data_out <= VN_data_out( 10091 downto 10086 );
    VN1681_sign_out <= VN_sign_out( 10091 downto 10086 );
    VN1682_data_out <= VN_data_out( 10097 downto 10092 );
    VN1682_sign_out <= VN_sign_out( 10097 downto 10092 );
    VN1683_data_out <= VN_data_out( 10103 downto 10098 );
    VN1683_sign_out <= VN_sign_out( 10103 downto 10098 );
    VN1684_data_out <= VN_data_out( 10109 downto 10104 );
    VN1684_sign_out <= VN_sign_out( 10109 downto 10104 );
    VN1685_data_out <= VN_data_out( 10115 downto 10110 );
    VN1685_sign_out <= VN_sign_out( 10115 downto 10110 );
    VN1686_data_out <= VN_data_out( 10121 downto 10116 );
    VN1686_sign_out <= VN_sign_out( 10121 downto 10116 );
    VN1687_data_out <= VN_data_out( 10127 downto 10122 );
    VN1687_sign_out <= VN_sign_out( 10127 downto 10122 );
    VN1688_data_out <= VN_data_out( 10133 downto 10128 );
    VN1688_sign_out <= VN_sign_out( 10133 downto 10128 );
    VN1689_data_out <= VN_data_out( 10139 downto 10134 );
    VN1689_sign_out <= VN_sign_out( 10139 downto 10134 );
    VN1690_data_out <= VN_data_out( 10145 downto 10140 );
    VN1690_sign_out <= VN_sign_out( 10145 downto 10140 );
    VN1691_data_out <= VN_data_out( 10151 downto 10146 );
    VN1691_sign_out <= VN_sign_out( 10151 downto 10146 );
    VN1692_data_out <= VN_data_out( 10157 downto 10152 );
    VN1692_sign_out <= VN_sign_out( 10157 downto 10152 );
    VN1693_data_out <= VN_data_out( 10163 downto 10158 );
    VN1693_sign_out <= VN_sign_out( 10163 downto 10158 );
    VN1694_data_out <= VN_data_out( 10169 downto 10164 );
    VN1694_sign_out <= VN_sign_out( 10169 downto 10164 );
    VN1695_data_out <= VN_data_out( 10175 downto 10170 );
    VN1695_sign_out <= VN_sign_out( 10175 downto 10170 );
    VN1696_data_out <= VN_data_out( 10181 downto 10176 );
    VN1696_sign_out <= VN_sign_out( 10181 downto 10176 );
    VN1697_data_out <= VN_data_out( 10187 downto 10182 );
    VN1697_sign_out <= VN_sign_out( 10187 downto 10182 );
    VN1698_data_out <= VN_data_out( 10193 downto 10188 );
    VN1698_sign_out <= VN_sign_out( 10193 downto 10188 );
    VN1699_data_out <= VN_data_out( 10199 downto 10194 );
    VN1699_sign_out <= VN_sign_out( 10199 downto 10194 );
    VN1700_data_out <= VN_data_out( 10205 downto 10200 );
    VN1700_sign_out <= VN_sign_out( 10205 downto 10200 );
    VN1701_data_out <= VN_data_out( 10211 downto 10206 );
    VN1701_sign_out <= VN_sign_out( 10211 downto 10206 );
    VN1702_data_out <= VN_data_out( 10217 downto 10212 );
    VN1702_sign_out <= VN_sign_out( 10217 downto 10212 );
    VN1703_data_out <= VN_data_out( 10223 downto 10218 );
    VN1703_sign_out <= VN_sign_out( 10223 downto 10218 );
    VN1704_data_out <= VN_data_out( 10229 downto 10224 );
    VN1704_sign_out <= VN_sign_out( 10229 downto 10224 );
    VN1705_data_out <= VN_data_out( 10235 downto 10230 );
    VN1705_sign_out <= VN_sign_out( 10235 downto 10230 );
    VN1706_data_out <= VN_data_out( 10241 downto 10236 );
    VN1706_sign_out <= VN_sign_out( 10241 downto 10236 );
    VN1707_data_out <= VN_data_out( 10247 downto 10242 );
    VN1707_sign_out <= VN_sign_out( 10247 downto 10242 );
    VN1708_data_out <= VN_data_out( 10253 downto 10248 );
    VN1708_sign_out <= VN_sign_out( 10253 downto 10248 );
    VN1709_data_out <= VN_data_out( 10259 downto 10254 );
    VN1709_sign_out <= VN_sign_out( 10259 downto 10254 );
    VN1710_data_out <= VN_data_out( 10265 downto 10260 );
    VN1710_sign_out <= VN_sign_out( 10265 downto 10260 );
    VN1711_data_out <= VN_data_out( 10271 downto 10266 );
    VN1711_sign_out <= VN_sign_out( 10271 downto 10266 );
    VN1712_data_out <= VN_data_out( 10277 downto 10272 );
    VN1712_sign_out <= VN_sign_out( 10277 downto 10272 );
    VN1713_data_out <= VN_data_out( 10283 downto 10278 );
    VN1713_sign_out <= VN_sign_out( 10283 downto 10278 );
    VN1714_data_out <= VN_data_out( 10289 downto 10284 );
    VN1714_sign_out <= VN_sign_out( 10289 downto 10284 );
    VN1715_data_out <= VN_data_out( 10295 downto 10290 );
    VN1715_sign_out <= VN_sign_out( 10295 downto 10290 );
    VN1716_data_out <= VN_data_out( 10301 downto 10296 );
    VN1716_sign_out <= VN_sign_out( 10301 downto 10296 );
    VN1717_data_out <= VN_data_out( 10307 downto 10302 );
    VN1717_sign_out <= VN_sign_out( 10307 downto 10302 );
    VN1718_data_out <= VN_data_out( 10313 downto 10308 );
    VN1718_sign_out <= VN_sign_out( 10313 downto 10308 );
    VN1719_data_out <= VN_data_out( 10319 downto 10314 );
    VN1719_sign_out <= VN_sign_out( 10319 downto 10314 );
    VN1720_data_out <= VN_data_out( 10325 downto 10320 );
    VN1720_sign_out <= VN_sign_out( 10325 downto 10320 );
    VN1721_data_out <= VN_data_out( 10331 downto 10326 );
    VN1721_sign_out <= VN_sign_out( 10331 downto 10326 );
    VN1722_data_out <= VN_data_out( 10337 downto 10332 );
    VN1722_sign_out <= VN_sign_out( 10337 downto 10332 );
    VN1723_data_out <= VN_data_out( 10343 downto 10338 );
    VN1723_sign_out <= VN_sign_out( 10343 downto 10338 );
    VN1724_data_out <= VN_data_out( 10349 downto 10344 );
    VN1724_sign_out <= VN_sign_out( 10349 downto 10344 );
    VN1725_data_out <= VN_data_out( 10355 downto 10350 );
    VN1725_sign_out <= VN_sign_out( 10355 downto 10350 );
    VN1726_data_out <= VN_data_out( 10361 downto 10356 );
    VN1726_sign_out <= VN_sign_out( 10361 downto 10356 );
    VN1727_data_out <= VN_data_out( 10367 downto 10362 );
    VN1727_sign_out <= VN_sign_out( 10367 downto 10362 );
    VN1728_data_out <= VN_data_out( 10373 downto 10368 );
    VN1728_sign_out <= VN_sign_out( 10373 downto 10368 );
    VN1729_data_out <= VN_data_out( 10379 downto 10374 );
    VN1729_sign_out <= VN_sign_out( 10379 downto 10374 );
    VN1730_data_out <= VN_data_out( 10385 downto 10380 );
    VN1730_sign_out <= VN_sign_out( 10385 downto 10380 );
    VN1731_data_out <= VN_data_out( 10391 downto 10386 );
    VN1731_sign_out <= VN_sign_out( 10391 downto 10386 );
    VN1732_data_out <= VN_data_out( 10397 downto 10392 );
    VN1732_sign_out <= VN_sign_out( 10397 downto 10392 );
    VN1733_data_out <= VN_data_out( 10403 downto 10398 );
    VN1733_sign_out <= VN_sign_out( 10403 downto 10398 );
    VN1734_data_out <= VN_data_out( 10409 downto 10404 );
    VN1734_sign_out <= VN_sign_out( 10409 downto 10404 );
    VN1735_data_out <= VN_data_out( 10415 downto 10410 );
    VN1735_sign_out <= VN_sign_out( 10415 downto 10410 );
    VN1736_data_out <= VN_data_out( 10421 downto 10416 );
    VN1736_sign_out <= VN_sign_out( 10421 downto 10416 );
    VN1737_data_out <= VN_data_out( 10427 downto 10422 );
    VN1737_sign_out <= VN_sign_out( 10427 downto 10422 );
    VN1738_data_out <= VN_data_out( 10433 downto 10428 );
    VN1738_sign_out <= VN_sign_out( 10433 downto 10428 );
    VN1739_data_out <= VN_data_out( 10439 downto 10434 );
    VN1739_sign_out <= VN_sign_out( 10439 downto 10434 );
    VN1740_data_out <= VN_data_out( 10445 downto 10440 );
    VN1740_sign_out <= VN_sign_out( 10445 downto 10440 );
    VN1741_data_out <= VN_data_out( 10451 downto 10446 );
    VN1741_sign_out <= VN_sign_out( 10451 downto 10446 );
    VN1742_data_out <= VN_data_out( 10457 downto 10452 );
    VN1742_sign_out <= VN_sign_out( 10457 downto 10452 );
    VN1743_data_out <= VN_data_out( 10463 downto 10458 );
    VN1743_sign_out <= VN_sign_out( 10463 downto 10458 );
    VN1744_data_out <= VN_data_out( 10469 downto 10464 );
    VN1744_sign_out <= VN_sign_out( 10469 downto 10464 );
    VN1745_data_out <= VN_data_out( 10475 downto 10470 );
    VN1745_sign_out <= VN_sign_out( 10475 downto 10470 );
    VN1746_data_out <= VN_data_out( 10481 downto 10476 );
    VN1746_sign_out <= VN_sign_out( 10481 downto 10476 );
    VN1747_data_out <= VN_data_out( 10487 downto 10482 );
    VN1747_sign_out <= VN_sign_out( 10487 downto 10482 );
    VN1748_data_out <= VN_data_out( 10493 downto 10488 );
    VN1748_sign_out <= VN_sign_out( 10493 downto 10488 );
    VN1749_data_out <= VN_data_out( 10499 downto 10494 );
    VN1749_sign_out <= VN_sign_out( 10499 downto 10494 );
    VN1750_data_out <= VN_data_out( 10505 downto 10500 );
    VN1750_sign_out <= VN_sign_out( 10505 downto 10500 );
    VN1751_data_out <= VN_data_out( 10511 downto 10506 );
    VN1751_sign_out <= VN_sign_out( 10511 downto 10506 );
    VN1752_data_out <= VN_data_out( 10517 downto 10512 );
    VN1752_sign_out <= VN_sign_out( 10517 downto 10512 );
    VN1753_data_out <= VN_data_out( 10523 downto 10518 );
    VN1753_sign_out <= VN_sign_out( 10523 downto 10518 );
    VN1754_data_out <= VN_data_out( 10529 downto 10524 );
    VN1754_sign_out <= VN_sign_out( 10529 downto 10524 );
    VN1755_data_out <= VN_data_out( 10535 downto 10530 );
    VN1755_sign_out <= VN_sign_out( 10535 downto 10530 );
    VN1756_data_out <= VN_data_out( 10541 downto 10536 );
    VN1756_sign_out <= VN_sign_out( 10541 downto 10536 );
    VN1757_data_out <= VN_data_out( 10547 downto 10542 );
    VN1757_sign_out <= VN_sign_out( 10547 downto 10542 );
    VN1758_data_out <= VN_data_out( 10553 downto 10548 );
    VN1758_sign_out <= VN_sign_out( 10553 downto 10548 );
    VN1759_data_out <= VN_data_out( 10559 downto 10554 );
    VN1759_sign_out <= VN_sign_out( 10559 downto 10554 );
    VN1760_data_out <= VN_data_out( 10565 downto 10560 );
    VN1760_sign_out <= VN_sign_out( 10565 downto 10560 );
    VN1761_data_out <= VN_data_out( 10571 downto 10566 );
    VN1761_sign_out <= VN_sign_out( 10571 downto 10566 );
    VN1762_data_out <= VN_data_out( 10577 downto 10572 );
    VN1762_sign_out <= VN_sign_out( 10577 downto 10572 );
    VN1763_data_out <= VN_data_out( 10583 downto 10578 );
    VN1763_sign_out <= VN_sign_out( 10583 downto 10578 );
    VN1764_data_out <= VN_data_out( 10589 downto 10584 );
    VN1764_sign_out <= VN_sign_out( 10589 downto 10584 );
    VN1765_data_out <= VN_data_out( 10595 downto 10590 );
    VN1765_sign_out <= VN_sign_out( 10595 downto 10590 );
    VN1766_data_out <= VN_data_out( 10601 downto 10596 );
    VN1766_sign_out <= VN_sign_out( 10601 downto 10596 );
    VN1767_data_out <= VN_data_out( 10607 downto 10602 );
    VN1767_sign_out <= VN_sign_out( 10607 downto 10602 );
    VN1768_data_out <= VN_data_out( 10613 downto 10608 );
    VN1768_sign_out <= VN_sign_out( 10613 downto 10608 );
    VN1769_data_out <= VN_data_out( 10619 downto 10614 );
    VN1769_sign_out <= VN_sign_out( 10619 downto 10614 );
    VN1770_data_out <= VN_data_out( 10625 downto 10620 );
    VN1770_sign_out <= VN_sign_out( 10625 downto 10620 );
    VN1771_data_out <= VN_data_out( 10631 downto 10626 );
    VN1771_sign_out <= VN_sign_out( 10631 downto 10626 );
    VN1772_data_out <= VN_data_out( 10637 downto 10632 );
    VN1772_sign_out <= VN_sign_out( 10637 downto 10632 );
    VN1773_data_out <= VN_data_out( 10643 downto 10638 );
    VN1773_sign_out <= VN_sign_out( 10643 downto 10638 );
    VN1774_data_out <= VN_data_out( 10649 downto 10644 );
    VN1774_sign_out <= VN_sign_out( 10649 downto 10644 );
    VN1775_data_out <= VN_data_out( 10655 downto 10650 );
    VN1775_sign_out <= VN_sign_out( 10655 downto 10650 );
    VN1776_data_out <= VN_data_out( 10661 downto 10656 );
    VN1776_sign_out <= VN_sign_out( 10661 downto 10656 );
    VN1777_data_out <= VN_data_out( 10667 downto 10662 );
    VN1777_sign_out <= VN_sign_out( 10667 downto 10662 );
    VN1778_data_out <= VN_data_out( 10673 downto 10668 );
    VN1778_sign_out <= VN_sign_out( 10673 downto 10668 );
    VN1779_data_out <= VN_data_out( 10679 downto 10674 );
    VN1779_sign_out <= VN_sign_out( 10679 downto 10674 );
    VN1780_data_out <= VN_data_out( 10685 downto 10680 );
    VN1780_sign_out <= VN_sign_out( 10685 downto 10680 );
    VN1781_data_out <= VN_data_out( 10691 downto 10686 );
    VN1781_sign_out <= VN_sign_out( 10691 downto 10686 );
    VN1782_data_out <= VN_data_out( 10697 downto 10692 );
    VN1782_sign_out <= VN_sign_out( 10697 downto 10692 );
    VN1783_data_out <= VN_data_out( 10703 downto 10698 );
    VN1783_sign_out <= VN_sign_out( 10703 downto 10698 );
    VN1784_data_out <= VN_data_out( 10709 downto 10704 );
    VN1784_sign_out <= VN_sign_out( 10709 downto 10704 );
    VN1785_data_out <= VN_data_out( 10715 downto 10710 );
    VN1785_sign_out <= VN_sign_out( 10715 downto 10710 );
    VN1786_data_out <= VN_data_out( 10721 downto 10716 );
    VN1786_sign_out <= VN_sign_out( 10721 downto 10716 );
    VN1787_data_out <= VN_data_out( 10727 downto 10722 );
    VN1787_sign_out <= VN_sign_out( 10727 downto 10722 );
    VN1788_data_out <= VN_data_out( 10733 downto 10728 );
    VN1788_sign_out <= VN_sign_out( 10733 downto 10728 );
    VN1789_data_out <= VN_data_out( 10739 downto 10734 );
    VN1789_sign_out <= VN_sign_out( 10739 downto 10734 );
    VN1790_data_out <= VN_data_out( 10745 downto 10740 );
    VN1790_sign_out <= VN_sign_out( 10745 downto 10740 );
    VN1791_data_out <= VN_data_out( 10751 downto 10746 );
    VN1791_sign_out <= VN_sign_out( 10751 downto 10746 );
    VN1792_data_out <= VN_data_out( 10757 downto 10752 );
    VN1792_sign_out <= VN_sign_out( 10757 downto 10752 );
    VN1793_data_out <= VN_data_out( 10763 downto 10758 );
    VN1793_sign_out <= VN_sign_out( 10763 downto 10758 );
    VN1794_data_out <= VN_data_out( 10769 downto 10764 );
    VN1794_sign_out <= VN_sign_out( 10769 downto 10764 );
    VN1795_data_out <= VN_data_out( 10775 downto 10770 );
    VN1795_sign_out <= VN_sign_out( 10775 downto 10770 );
    VN1796_data_out <= VN_data_out( 10781 downto 10776 );
    VN1796_sign_out <= VN_sign_out( 10781 downto 10776 );
    VN1797_data_out <= VN_data_out( 10787 downto 10782 );
    VN1797_sign_out <= VN_sign_out( 10787 downto 10782 );
    VN1798_data_out <= VN_data_out( 10793 downto 10788 );
    VN1798_sign_out <= VN_sign_out( 10793 downto 10788 );
    VN1799_data_out <= VN_data_out( 10799 downto 10794 );
    VN1799_sign_out <= VN_sign_out( 10799 downto 10794 );
    VN1800_data_out <= VN_data_out( 10805 downto 10800 );
    VN1800_sign_out <= VN_sign_out( 10805 downto 10800 );
    VN1801_data_out <= VN_data_out( 10811 downto 10806 );
    VN1801_sign_out <= VN_sign_out( 10811 downto 10806 );
    VN1802_data_out <= VN_data_out( 10817 downto 10812 );
    VN1802_sign_out <= VN_sign_out( 10817 downto 10812 );
    VN1803_data_out <= VN_data_out( 10823 downto 10818 );
    VN1803_sign_out <= VN_sign_out( 10823 downto 10818 );
    VN1804_data_out <= VN_data_out( 10829 downto 10824 );
    VN1804_sign_out <= VN_sign_out( 10829 downto 10824 );
    VN1805_data_out <= VN_data_out( 10835 downto 10830 );
    VN1805_sign_out <= VN_sign_out( 10835 downto 10830 );
    VN1806_data_out <= VN_data_out( 10841 downto 10836 );
    VN1806_sign_out <= VN_sign_out( 10841 downto 10836 );
    VN1807_data_out <= VN_data_out( 10847 downto 10842 );
    VN1807_sign_out <= VN_sign_out( 10847 downto 10842 );
    VN1808_data_out <= VN_data_out( 10853 downto 10848 );
    VN1808_sign_out <= VN_sign_out( 10853 downto 10848 );
    VN1809_data_out <= VN_data_out( 10859 downto 10854 );
    VN1809_sign_out <= VN_sign_out( 10859 downto 10854 );
    VN1810_data_out <= VN_data_out( 10865 downto 10860 );
    VN1810_sign_out <= VN_sign_out( 10865 downto 10860 );
    VN1811_data_out <= VN_data_out( 10871 downto 10866 );
    VN1811_sign_out <= VN_sign_out( 10871 downto 10866 );
    VN1812_data_out <= VN_data_out( 10877 downto 10872 );
    VN1812_sign_out <= VN_sign_out( 10877 downto 10872 );
    VN1813_data_out <= VN_data_out( 10883 downto 10878 );
    VN1813_sign_out <= VN_sign_out( 10883 downto 10878 );
    VN1814_data_out <= VN_data_out( 10889 downto 10884 );
    VN1814_sign_out <= VN_sign_out( 10889 downto 10884 );
    VN1815_data_out <= VN_data_out( 10895 downto 10890 );
    VN1815_sign_out <= VN_sign_out( 10895 downto 10890 );
    VN1816_data_out <= VN_data_out( 10901 downto 10896 );
    VN1816_sign_out <= VN_sign_out( 10901 downto 10896 );
    VN1817_data_out <= VN_data_out( 10907 downto 10902 );
    VN1817_sign_out <= VN_sign_out( 10907 downto 10902 );
    VN1818_data_out <= VN_data_out( 10913 downto 10908 );
    VN1818_sign_out <= VN_sign_out( 10913 downto 10908 );
    VN1819_data_out <= VN_data_out( 10919 downto 10914 );
    VN1819_sign_out <= VN_sign_out( 10919 downto 10914 );
    VN1820_data_out <= VN_data_out( 10925 downto 10920 );
    VN1820_sign_out <= VN_sign_out( 10925 downto 10920 );
    VN1821_data_out <= VN_data_out( 10931 downto 10926 );
    VN1821_sign_out <= VN_sign_out( 10931 downto 10926 );
    VN1822_data_out <= VN_data_out( 10937 downto 10932 );
    VN1822_sign_out <= VN_sign_out( 10937 downto 10932 );
    VN1823_data_out <= VN_data_out( 10943 downto 10938 );
    VN1823_sign_out <= VN_sign_out( 10943 downto 10938 );
    VN1824_data_out <= VN_data_out( 10949 downto 10944 );
    VN1824_sign_out <= VN_sign_out( 10949 downto 10944 );
    VN1825_data_out <= VN_data_out( 10955 downto 10950 );
    VN1825_sign_out <= VN_sign_out( 10955 downto 10950 );
    VN1826_data_out <= VN_data_out( 10961 downto 10956 );
    VN1826_sign_out <= VN_sign_out( 10961 downto 10956 );
    VN1827_data_out <= VN_data_out( 10967 downto 10962 );
    VN1827_sign_out <= VN_sign_out( 10967 downto 10962 );
    VN1828_data_out <= VN_data_out( 10973 downto 10968 );
    VN1828_sign_out <= VN_sign_out( 10973 downto 10968 );
    VN1829_data_out <= VN_data_out( 10979 downto 10974 );
    VN1829_sign_out <= VN_sign_out( 10979 downto 10974 );
    VN1830_data_out <= VN_data_out( 10985 downto 10980 );
    VN1830_sign_out <= VN_sign_out( 10985 downto 10980 );
    VN1831_data_out <= VN_data_out( 10991 downto 10986 );
    VN1831_sign_out <= VN_sign_out( 10991 downto 10986 );
    VN1832_data_out <= VN_data_out( 10997 downto 10992 );
    VN1832_sign_out <= VN_sign_out( 10997 downto 10992 );
    VN1833_data_out <= VN_data_out( 11003 downto 10998 );
    VN1833_sign_out <= VN_sign_out( 11003 downto 10998 );
    VN1834_data_out <= VN_data_out( 11009 downto 11004 );
    VN1834_sign_out <= VN_sign_out( 11009 downto 11004 );
    VN1835_data_out <= VN_data_out( 11015 downto 11010 );
    VN1835_sign_out <= VN_sign_out( 11015 downto 11010 );
    VN1836_data_out <= VN_data_out( 11021 downto 11016 );
    VN1836_sign_out <= VN_sign_out( 11021 downto 11016 );
    VN1837_data_out <= VN_data_out( 11027 downto 11022 );
    VN1837_sign_out <= VN_sign_out( 11027 downto 11022 );
    VN1838_data_out <= VN_data_out( 11033 downto 11028 );
    VN1838_sign_out <= VN_sign_out( 11033 downto 11028 );
    VN1839_data_out <= VN_data_out( 11039 downto 11034 );
    VN1839_sign_out <= VN_sign_out( 11039 downto 11034 );
    VN1840_data_out <= VN_data_out( 11045 downto 11040 );
    VN1840_sign_out <= VN_sign_out( 11045 downto 11040 );
    VN1841_data_out <= VN_data_out( 11051 downto 11046 );
    VN1841_sign_out <= VN_sign_out( 11051 downto 11046 );
    VN1842_data_out <= VN_data_out( 11057 downto 11052 );
    VN1842_sign_out <= VN_sign_out( 11057 downto 11052 );
    VN1843_data_out <= VN_data_out( 11063 downto 11058 );
    VN1843_sign_out <= VN_sign_out( 11063 downto 11058 );
    VN1844_data_out <= VN_data_out( 11069 downto 11064 );
    VN1844_sign_out <= VN_sign_out( 11069 downto 11064 );
    VN1845_data_out <= VN_data_out( 11075 downto 11070 );
    VN1845_sign_out <= VN_sign_out( 11075 downto 11070 );
    VN1846_data_out <= VN_data_out( 11081 downto 11076 );
    VN1846_sign_out <= VN_sign_out( 11081 downto 11076 );
    VN1847_data_out <= VN_data_out( 11087 downto 11082 );
    VN1847_sign_out <= VN_sign_out( 11087 downto 11082 );
    VN1848_data_out <= VN_data_out( 11093 downto 11088 );
    VN1848_sign_out <= VN_sign_out( 11093 downto 11088 );
    VN1849_data_out <= VN_data_out( 11099 downto 11094 );
    VN1849_sign_out <= VN_sign_out( 11099 downto 11094 );
    VN1850_data_out <= VN_data_out( 11105 downto 11100 );
    VN1850_sign_out <= VN_sign_out( 11105 downto 11100 );
    VN1851_data_out <= VN_data_out( 11111 downto 11106 );
    VN1851_sign_out <= VN_sign_out( 11111 downto 11106 );
    VN1852_data_out <= VN_data_out( 11117 downto 11112 );
    VN1852_sign_out <= VN_sign_out( 11117 downto 11112 );
    VN1853_data_out <= VN_data_out( 11123 downto 11118 );
    VN1853_sign_out <= VN_sign_out( 11123 downto 11118 );
    VN1854_data_out <= VN_data_out( 11129 downto 11124 );
    VN1854_sign_out <= VN_sign_out( 11129 downto 11124 );
    VN1855_data_out <= VN_data_out( 11135 downto 11130 );
    VN1855_sign_out <= VN_sign_out( 11135 downto 11130 );
    VN1856_data_out <= VN_data_out( 11141 downto 11136 );
    VN1856_sign_out <= VN_sign_out( 11141 downto 11136 );
    VN1857_data_out <= VN_data_out( 11147 downto 11142 );
    VN1857_sign_out <= VN_sign_out( 11147 downto 11142 );
    VN1858_data_out <= VN_data_out( 11153 downto 11148 );
    VN1858_sign_out <= VN_sign_out( 11153 downto 11148 );
    VN1859_data_out <= VN_data_out( 11159 downto 11154 );
    VN1859_sign_out <= VN_sign_out( 11159 downto 11154 );
    VN1860_data_out <= VN_data_out( 11165 downto 11160 );
    VN1860_sign_out <= VN_sign_out( 11165 downto 11160 );
    VN1861_data_out <= VN_data_out( 11171 downto 11166 );
    VN1861_sign_out <= VN_sign_out( 11171 downto 11166 );
    VN1862_data_out <= VN_data_out( 11177 downto 11172 );
    VN1862_sign_out <= VN_sign_out( 11177 downto 11172 );
    VN1863_data_out <= VN_data_out( 11183 downto 11178 );
    VN1863_sign_out <= VN_sign_out( 11183 downto 11178 );
    VN1864_data_out <= VN_data_out( 11189 downto 11184 );
    VN1864_sign_out <= VN_sign_out( 11189 downto 11184 );
    VN1865_data_out <= VN_data_out( 11195 downto 11190 );
    VN1865_sign_out <= VN_sign_out( 11195 downto 11190 );
    VN1866_data_out <= VN_data_out( 11201 downto 11196 );
    VN1866_sign_out <= VN_sign_out( 11201 downto 11196 );
    VN1867_data_out <= VN_data_out( 11207 downto 11202 );
    VN1867_sign_out <= VN_sign_out( 11207 downto 11202 );
    VN1868_data_out <= VN_data_out( 11213 downto 11208 );
    VN1868_sign_out <= VN_sign_out( 11213 downto 11208 );
    VN1869_data_out <= VN_data_out( 11219 downto 11214 );
    VN1869_sign_out <= VN_sign_out( 11219 downto 11214 );
    VN1870_data_out <= VN_data_out( 11225 downto 11220 );
    VN1870_sign_out <= VN_sign_out( 11225 downto 11220 );
    VN1871_data_out <= VN_data_out( 11231 downto 11226 );
    VN1871_sign_out <= VN_sign_out( 11231 downto 11226 );
    VN1872_data_out <= VN_data_out( 11237 downto 11232 );
    VN1872_sign_out <= VN_sign_out( 11237 downto 11232 );
    VN1873_data_out <= VN_data_out( 11243 downto 11238 );
    VN1873_sign_out <= VN_sign_out( 11243 downto 11238 );
    VN1874_data_out <= VN_data_out( 11249 downto 11244 );
    VN1874_sign_out <= VN_sign_out( 11249 downto 11244 );
    VN1875_data_out <= VN_data_out( 11255 downto 11250 );
    VN1875_sign_out <= VN_sign_out( 11255 downto 11250 );
    VN1876_data_out <= VN_data_out( 11261 downto 11256 );
    VN1876_sign_out <= VN_sign_out( 11261 downto 11256 );
    VN1877_data_out <= VN_data_out( 11267 downto 11262 );
    VN1877_sign_out <= VN_sign_out( 11267 downto 11262 );
    VN1878_data_out <= VN_data_out( 11273 downto 11268 );
    VN1878_sign_out <= VN_sign_out( 11273 downto 11268 );
    VN1879_data_out <= VN_data_out( 11279 downto 11274 );
    VN1879_sign_out <= VN_sign_out( 11279 downto 11274 );
    VN1880_data_out <= VN_data_out( 11285 downto 11280 );
    VN1880_sign_out <= VN_sign_out( 11285 downto 11280 );
    VN1881_data_out <= VN_data_out( 11291 downto 11286 );
    VN1881_sign_out <= VN_sign_out( 11291 downto 11286 );
    VN1882_data_out <= VN_data_out( 11297 downto 11292 );
    VN1882_sign_out <= VN_sign_out( 11297 downto 11292 );
    VN1883_data_out <= VN_data_out( 11303 downto 11298 );
    VN1883_sign_out <= VN_sign_out( 11303 downto 11298 );
    VN1884_data_out <= VN_data_out( 11309 downto 11304 );
    VN1884_sign_out <= VN_sign_out( 11309 downto 11304 );
    VN1885_data_out <= VN_data_out( 11315 downto 11310 );
    VN1885_sign_out <= VN_sign_out( 11315 downto 11310 );
    VN1886_data_out <= VN_data_out( 11321 downto 11316 );
    VN1886_sign_out <= VN_sign_out( 11321 downto 11316 );
    VN1887_data_out <= VN_data_out( 11327 downto 11322 );
    VN1887_sign_out <= VN_sign_out( 11327 downto 11322 );
    VN1888_data_out <= VN_data_out( 11333 downto 11328 );
    VN1888_sign_out <= VN_sign_out( 11333 downto 11328 );
    VN1889_data_out <= VN_data_out( 11339 downto 11334 );
    VN1889_sign_out <= VN_sign_out( 11339 downto 11334 );
    VN1890_data_out <= VN_data_out( 11345 downto 11340 );
    VN1890_sign_out <= VN_sign_out( 11345 downto 11340 );
    VN1891_data_out <= VN_data_out( 11351 downto 11346 );
    VN1891_sign_out <= VN_sign_out( 11351 downto 11346 );
    VN1892_data_out <= VN_data_out( 11357 downto 11352 );
    VN1892_sign_out <= VN_sign_out( 11357 downto 11352 );
    VN1893_data_out <= VN_data_out( 11363 downto 11358 );
    VN1893_sign_out <= VN_sign_out( 11363 downto 11358 );
    VN1894_data_out <= VN_data_out( 11369 downto 11364 );
    VN1894_sign_out <= VN_sign_out( 11369 downto 11364 );
    VN1895_data_out <= VN_data_out( 11375 downto 11370 );
    VN1895_sign_out <= VN_sign_out( 11375 downto 11370 );
    VN1896_data_out <= VN_data_out( 11381 downto 11376 );
    VN1896_sign_out <= VN_sign_out( 11381 downto 11376 );
    VN1897_data_out <= VN_data_out( 11387 downto 11382 );
    VN1897_sign_out <= VN_sign_out( 11387 downto 11382 );
    VN1898_data_out <= VN_data_out( 11393 downto 11388 );
    VN1898_sign_out <= VN_sign_out( 11393 downto 11388 );
    VN1899_data_out <= VN_data_out( 11399 downto 11394 );
    VN1899_sign_out <= VN_sign_out( 11399 downto 11394 );
    VN1900_data_out <= VN_data_out( 11405 downto 11400 );
    VN1900_sign_out <= VN_sign_out( 11405 downto 11400 );
    VN1901_data_out <= VN_data_out( 11411 downto 11406 );
    VN1901_sign_out <= VN_sign_out( 11411 downto 11406 );
    VN1902_data_out <= VN_data_out( 11417 downto 11412 );
    VN1902_sign_out <= VN_sign_out( 11417 downto 11412 );
    VN1903_data_out <= VN_data_out( 11423 downto 11418 );
    VN1903_sign_out <= VN_sign_out( 11423 downto 11418 );
    VN1904_data_out <= VN_data_out( 11429 downto 11424 );
    VN1904_sign_out <= VN_sign_out( 11429 downto 11424 );
    VN1905_data_out <= VN_data_out( 11435 downto 11430 );
    VN1905_sign_out <= VN_sign_out( 11435 downto 11430 );
    VN1906_data_out <= VN_data_out( 11441 downto 11436 );
    VN1906_sign_out <= VN_sign_out( 11441 downto 11436 );
    VN1907_data_out <= VN_data_out( 11447 downto 11442 );
    VN1907_sign_out <= VN_sign_out( 11447 downto 11442 );
    VN1908_data_out <= VN_data_out( 11453 downto 11448 );
    VN1908_sign_out <= VN_sign_out( 11453 downto 11448 );
    VN1909_data_out <= VN_data_out( 11459 downto 11454 );
    VN1909_sign_out <= VN_sign_out( 11459 downto 11454 );
    VN1910_data_out <= VN_data_out( 11465 downto 11460 );
    VN1910_sign_out <= VN_sign_out( 11465 downto 11460 );
    VN1911_data_out <= VN_data_out( 11471 downto 11466 );
    VN1911_sign_out <= VN_sign_out( 11471 downto 11466 );
    VN1912_data_out <= VN_data_out( 11477 downto 11472 );
    VN1912_sign_out <= VN_sign_out( 11477 downto 11472 );
    VN1913_data_out <= VN_data_out( 11483 downto 11478 );
    VN1913_sign_out <= VN_sign_out( 11483 downto 11478 );
    VN1914_data_out <= VN_data_out( 11489 downto 11484 );
    VN1914_sign_out <= VN_sign_out( 11489 downto 11484 );
    VN1915_data_out <= VN_data_out( 11495 downto 11490 );
    VN1915_sign_out <= VN_sign_out( 11495 downto 11490 );
    VN1916_data_out <= VN_data_out( 11501 downto 11496 );
    VN1916_sign_out <= VN_sign_out( 11501 downto 11496 );
    VN1917_data_out <= VN_data_out( 11507 downto 11502 );
    VN1917_sign_out <= VN_sign_out( 11507 downto 11502 );
    VN1918_data_out <= VN_data_out( 11513 downto 11508 );
    VN1918_sign_out <= VN_sign_out( 11513 downto 11508 );
    VN1919_data_out <= VN_data_out( 11519 downto 11514 );
    VN1919_sign_out <= VN_sign_out( 11519 downto 11514 );
    VN1920_data_out <= VN_data_out( 11525 downto 11520 );
    VN1920_sign_out <= VN_sign_out( 11525 downto 11520 );
    VN1921_data_out <= VN_data_out( 11531 downto 11526 );
    VN1921_sign_out <= VN_sign_out( 11531 downto 11526 );
    VN1922_data_out <= VN_data_out( 11537 downto 11532 );
    VN1922_sign_out <= VN_sign_out( 11537 downto 11532 );
    VN1923_data_out <= VN_data_out( 11543 downto 11538 );
    VN1923_sign_out <= VN_sign_out( 11543 downto 11538 );
    VN1924_data_out <= VN_data_out( 11549 downto 11544 );
    VN1924_sign_out <= VN_sign_out( 11549 downto 11544 );
    VN1925_data_out <= VN_data_out( 11555 downto 11550 );
    VN1925_sign_out <= VN_sign_out( 11555 downto 11550 );
    VN1926_data_out <= VN_data_out( 11561 downto 11556 );
    VN1926_sign_out <= VN_sign_out( 11561 downto 11556 );
    VN1927_data_out <= VN_data_out( 11567 downto 11562 );
    VN1927_sign_out <= VN_sign_out( 11567 downto 11562 );
    VN1928_data_out <= VN_data_out( 11573 downto 11568 );
    VN1928_sign_out <= VN_sign_out( 11573 downto 11568 );
    VN1929_data_out <= VN_data_out( 11579 downto 11574 );
    VN1929_sign_out <= VN_sign_out( 11579 downto 11574 );
    VN1930_data_out <= VN_data_out( 11585 downto 11580 );
    VN1930_sign_out <= VN_sign_out( 11585 downto 11580 );
    VN1931_data_out <= VN_data_out( 11591 downto 11586 );
    VN1931_sign_out <= VN_sign_out( 11591 downto 11586 );
    VN1932_data_out <= VN_data_out( 11597 downto 11592 );
    VN1932_sign_out <= VN_sign_out( 11597 downto 11592 );
    VN1933_data_out <= VN_data_out( 11603 downto 11598 );
    VN1933_sign_out <= VN_sign_out( 11603 downto 11598 );
    VN1934_data_out <= VN_data_out( 11609 downto 11604 );
    VN1934_sign_out <= VN_sign_out( 11609 downto 11604 );
    VN1935_data_out <= VN_data_out( 11615 downto 11610 );
    VN1935_sign_out <= VN_sign_out( 11615 downto 11610 );
    VN1936_data_out <= VN_data_out( 11621 downto 11616 );
    VN1936_sign_out <= VN_sign_out( 11621 downto 11616 );
    VN1937_data_out <= VN_data_out( 11627 downto 11622 );
    VN1937_sign_out <= VN_sign_out( 11627 downto 11622 );
    VN1938_data_out <= VN_data_out( 11633 downto 11628 );
    VN1938_sign_out <= VN_sign_out( 11633 downto 11628 );
    VN1939_data_out <= VN_data_out( 11639 downto 11634 );
    VN1939_sign_out <= VN_sign_out( 11639 downto 11634 );
    VN1940_data_out <= VN_data_out( 11645 downto 11640 );
    VN1940_sign_out <= VN_sign_out( 11645 downto 11640 );
    VN1941_data_out <= VN_data_out( 11651 downto 11646 );
    VN1941_sign_out <= VN_sign_out( 11651 downto 11646 );
    VN1942_data_out <= VN_data_out( 11657 downto 11652 );
    VN1942_sign_out <= VN_sign_out( 11657 downto 11652 );
    VN1943_data_out <= VN_data_out( 11663 downto 11658 );
    VN1943_sign_out <= VN_sign_out( 11663 downto 11658 );
    VN1944_data_out <= VN_data_out( 11669 downto 11664 );
    VN1944_sign_out <= VN_sign_out( 11669 downto 11664 );
    VN1945_data_out <= VN_data_out( 11675 downto 11670 );
    VN1945_sign_out <= VN_sign_out( 11675 downto 11670 );
    VN1946_data_out <= VN_data_out( 11681 downto 11676 );
    VN1946_sign_out <= VN_sign_out( 11681 downto 11676 );
    VN1947_data_out <= VN_data_out( 11687 downto 11682 );
    VN1947_sign_out <= VN_sign_out( 11687 downto 11682 );
    VN1948_data_out <= VN_data_out( 11693 downto 11688 );
    VN1948_sign_out <= VN_sign_out( 11693 downto 11688 );
    VN1949_data_out <= VN_data_out( 11699 downto 11694 );
    VN1949_sign_out <= VN_sign_out( 11699 downto 11694 );
    VN1950_data_out <= VN_data_out( 11705 downto 11700 );
    VN1950_sign_out <= VN_sign_out( 11705 downto 11700 );
    VN1951_data_out <= VN_data_out( 11711 downto 11706 );
    VN1951_sign_out <= VN_sign_out( 11711 downto 11706 );
    VN1952_data_out <= VN_data_out( 11717 downto 11712 );
    VN1952_sign_out <= VN_sign_out( 11717 downto 11712 );
    VN1953_data_out <= VN_data_out( 11723 downto 11718 );
    VN1953_sign_out <= VN_sign_out( 11723 downto 11718 );
    VN1954_data_out <= VN_data_out( 11729 downto 11724 );
    VN1954_sign_out <= VN_sign_out( 11729 downto 11724 );
    VN1955_data_out <= VN_data_out( 11735 downto 11730 );
    VN1955_sign_out <= VN_sign_out( 11735 downto 11730 );
    VN1956_data_out <= VN_data_out( 11741 downto 11736 );
    VN1956_sign_out <= VN_sign_out( 11741 downto 11736 );
    VN1957_data_out <= VN_data_out( 11747 downto 11742 );
    VN1957_sign_out <= VN_sign_out( 11747 downto 11742 );
    VN1958_data_out <= VN_data_out( 11753 downto 11748 );
    VN1958_sign_out <= VN_sign_out( 11753 downto 11748 );
    VN1959_data_out <= VN_data_out( 11759 downto 11754 );
    VN1959_sign_out <= VN_sign_out( 11759 downto 11754 );
    VN1960_data_out <= VN_data_out( 11765 downto 11760 );
    VN1960_sign_out <= VN_sign_out( 11765 downto 11760 );
    VN1961_data_out <= VN_data_out( 11771 downto 11766 );
    VN1961_sign_out <= VN_sign_out( 11771 downto 11766 );
    VN1962_data_out <= VN_data_out( 11777 downto 11772 );
    VN1962_sign_out <= VN_sign_out( 11777 downto 11772 );
    VN1963_data_out <= VN_data_out( 11783 downto 11778 );
    VN1963_sign_out <= VN_sign_out( 11783 downto 11778 );
    VN1964_data_out <= VN_data_out( 11789 downto 11784 );
    VN1964_sign_out <= VN_sign_out( 11789 downto 11784 );
    VN1965_data_out <= VN_data_out( 11795 downto 11790 );
    VN1965_sign_out <= VN_sign_out( 11795 downto 11790 );
    VN1966_data_out <= VN_data_out( 11801 downto 11796 );
    VN1966_sign_out <= VN_sign_out( 11801 downto 11796 );
    VN1967_data_out <= VN_data_out( 11807 downto 11802 );
    VN1967_sign_out <= VN_sign_out( 11807 downto 11802 );
    VN1968_data_out <= VN_data_out( 11813 downto 11808 );
    VN1968_sign_out <= VN_sign_out( 11813 downto 11808 );
    VN1969_data_out <= VN_data_out( 11819 downto 11814 );
    VN1969_sign_out <= VN_sign_out( 11819 downto 11814 );
    VN1970_data_out <= VN_data_out( 11825 downto 11820 );
    VN1970_sign_out <= VN_sign_out( 11825 downto 11820 );
    VN1971_data_out <= VN_data_out( 11831 downto 11826 );
    VN1971_sign_out <= VN_sign_out( 11831 downto 11826 );
    VN1972_data_out <= VN_data_out( 11837 downto 11832 );
    VN1972_sign_out <= VN_sign_out( 11837 downto 11832 );
    VN1973_data_out <= VN_data_out( 11843 downto 11838 );
    VN1973_sign_out <= VN_sign_out( 11843 downto 11838 );
    VN1974_data_out <= VN_data_out( 11849 downto 11844 );
    VN1974_sign_out <= VN_sign_out( 11849 downto 11844 );
    VN1975_data_out <= VN_data_out( 11855 downto 11850 );
    VN1975_sign_out <= VN_sign_out( 11855 downto 11850 );
    VN1976_data_out <= VN_data_out( 11861 downto 11856 );
    VN1976_sign_out <= VN_sign_out( 11861 downto 11856 );
    VN1977_data_out <= VN_data_out( 11867 downto 11862 );
    VN1977_sign_out <= VN_sign_out( 11867 downto 11862 );
    VN1978_data_out <= VN_data_out( 11873 downto 11868 );
    VN1978_sign_out <= VN_sign_out( 11873 downto 11868 );
    VN1979_data_out <= VN_data_out( 11879 downto 11874 );
    VN1979_sign_out <= VN_sign_out( 11879 downto 11874 );
    VN1980_data_out <= VN_data_out( 11885 downto 11880 );
    VN1980_sign_out <= VN_sign_out( 11885 downto 11880 );
    VN1981_data_out <= VN_data_out( 11891 downto 11886 );
    VN1981_sign_out <= VN_sign_out( 11891 downto 11886 );
    VN1982_data_out <= VN_data_out( 11897 downto 11892 );
    VN1982_sign_out <= VN_sign_out( 11897 downto 11892 );
    VN1983_data_out <= VN_data_out( 11903 downto 11898 );
    VN1983_sign_out <= VN_sign_out( 11903 downto 11898 );
    VN1984_data_out <= VN_data_out( 11909 downto 11904 );
    VN1984_sign_out <= VN_sign_out( 11909 downto 11904 );
    VN1985_data_out <= VN_data_out( 11915 downto 11910 );
    VN1985_sign_out <= VN_sign_out( 11915 downto 11910 );
    VN1986_data_out <= VN_data_out( 11921 downto 11916 );
    VN1986_sign_out <= VN_sign_out( 11921 downto 11916 );
    VN1987_data_out <= VN_data_out( 11927 downto 11922 );
    VN1987_sign_out <= VN_sign_out( 11927 downto 11922 );
    VN1988_data_out <= VN_data_out( 11933 downto 11928 );
    VN1988_sign_out <= VN_sign_out( 11933 downto 11928 );
    VN1989_data_out <= VN_data_out( 11939 downto 11934 );
    VN1989_sign_out <= VN_sign_out( 11939 downto 11934 );
    VN1990_data_out <= VN_data_out( 11945 downto 11940 );
    VN1990_sign_out <= VN_sign_out( 11945 downto 11940 );
    VN1991_data_out <= VN_data_out( 11951 downto 11946 );
    VN1991_sign_out <= VN_sign_out( 11951 downto 11946 );
    VN1992_data_out <= VN_data_out( 11957 downto 11952 );
    VN1992_sign_out <= VN_sign_out( 11957 downto 11952 );
    VN1993_data_out <= VN_data_out( 11963 downto 11958 );
    VN1993_sign_out <= VN_sign_out( 11963 downto 11958 );
    VN1994_data_out <= VN_data_out( 11969 downto 11964 );
    VN1994_sign_out <= VN_sign_out( 11969 downto 11964 );
    VN1995_data_out <= VN_data_out( 11975 downto 11970 );
    VN1995_sign_out <= VN_sign_out( 11975 downto 11970 );
    VN1996_data_out <= VN_data_out( 11981 downto 11976 );
    VN1996_sign_out <= VN_sign_out( 11981 downto 11976 );
    VN1997_data_out <= VN_data_out( 11987 downto 11982 );
    VN1997_sign_out <= VN_sign_out( 11987 downto 11982 );
    VN1998_data_out <= VN_data_out( 11993 downto 11988 );
    VN1998_sign_out <= VN_sign_out( 11993 downto 11988 );
    VN1999_data_out <= VN_data_out( 11999 downto 11994 );
    VN1999_sign_out <= VN_sign_out( 11999 downto 11994 );
    VN2000_data_out <= VN_data_out( 12005 downto 12000 );
    VN2000_sign_out <= VN_sign_out( 12005 downto 12000 );
    VN2001_data_out <= VN_data_out( 12011 downto 12006 );
    VN2001_sign_out <= VN_sign_out( 12011 downto 12006 );
    VN2002_data_out <= VN_data_out( 12017 downto 12012 );
    VN2002_sign_out <= VN_sign_out( 12017 downto 12012 );
    VN2003_data_out <= VN_data_out( 12023 downto 12018 );
    VN2003_sign_out <= VN_sign_out( 12023 downto 12018 );
    VN2004_data_out <= VN_data_out( 12029 downto 12024 );
    VN2004_sign_out <= VN_sign_out( 12029 downto 12024 );
    VN2005_data_out <= VN_data_out( 12035 downto 12030 );
    VN2005_sign_out <= VN_sign_out( 12035 downto 12030 );
    VN2006_data_out <= VN_data_out( 12041 downto 12036 );
    VN2006_sign_out <= VN_sign_out( 12041 downto 12036 );
    VN2007_data_out <= VN_data_out( 12047 downto 12042 );
    VN2007_sign_out <= VN_sign_out( 12047 downto 12042 );
    VN2008_data_out <= VN_data_out( 12053 downto 12048 );
    VN2008_sign_out <= VN_sign_out( 12053 downto 12048 );
    VN2009_data_out <= VN_data_out( 12059 downto 12054 );
    VN2009_sign_out <= VN_sign_out( 12059 downto 12054 );
    VN2010_data_out <= VN_data_out( 12065 downto 12060 );
    VN2010_sign_out <= VN_sign_out( 12065 downto 12060 );
    VN2011_data_out <= VN_data_out( 12071 downto 12066 );
    VN2011_sign_out <= VN_sign_out( 12071 downto 12066 );
    VN2012_data_out <= VN_data_out( 12077 downto 12072 );
    VN2012_sign_out <= VN_sign_out( 12077 downto 12072 );
    VN2013_data_out <= VN_data_out( 12083 downto 12078 );
    VN2013_sign_out <= VN_sign_out( 12083 downto 12078 );
    VN2014_data_out <= VN_data_out( 12089 downto 12084 );
    VN2014_sign_out <= VN_sign_out( 12089 downto 12084 );
    VN2015_data_out <= VN_data_out( 12095 downto 12090 );
    VN2015_sign_out <= VN_sign_out( 12095 downto 12090 );
    VN2016_data_out <= VN_data_out( 12101 downto 12096 );
    VN2016_sign_out <= VN_sign_out( 12101 downto 12096 );
    VN2017_data_out <= VN_data_out( 12107 downto 12102 );
    VN2017_sign_out <= VN_sign_out( 12107 downto 12102 );
    VN2018_data_out <= VN_data_out( 12113 downto 12108 );
    VN2018_sign_out <= VN_sign_out( 12113 downto 12108 );
    VN2019_data_out <= VN_data_out( 12119 downto 12114 );
    VN2019_sign_out <= VN_sign_out( 12119 downto 12114 );
    VN2020_data_out <= VN_data_out( 12125 downto 12120 );
    VN2020_sign_out <= VN_sign_out( 12125 downto 12120 );
    VN2021_data_out <= VN_data_out( 12131 downto 12126 );
    VN2021_sign_out <= VN_sign_out( 12131 downto 12126 );
    VN2022_data_out <= VN_data_out( 12137 downto 12132 );
    VN2022_sign_out <= VN_sign_out( 12137 downto 12132 );
    VN2023_data_out <= VN_data_out( 12143 downto 12138 );
    VN2023_sign_out <= VN_sign_out( 12143 downto 12138 );
    VN2024_data_out <= VN_data_out( 12149 downto 12144 );
    VN2024_sign_out <= VN_sign_out( 12149 downto 12144 );
    VN2025_data_out <= VN_data_out( 12155 downto 12150 );
    VN2025_sign_out <= VN_sign_out( 12155 downto 12150 );
    VN2026_data_out <= VN_data_out( 12161 downto 12156 );
    VN2026_sign_out <= VN_sign_out( 12161 downto 12156 );
    VN2027_data_out <= VN_data_out( 12167 downto 12162 );
    VN2027_sign_out <= VN_sign_out( 12167 downto 12162 );
    VN2028_data_out <= VN_data_out( 12173 downto 12168 );
    VN2028_sign_out <= VN_sign_out( 12173 downto 12168 );
    VN2029_data_out <= VN_data_out( 12179 downto 12174 );
    VN2029_sign_out <= VN_sign_out( 12179 downto 12174 );
    VN2030_data_out <= VN_data_out( 12185 downto 12180 );
    VN2030_sign_out <= VN_sign_out( 12185 downto 12180 );
    VN2031_data_out <= VN_data_out( 12191 downto 12186 );
    VN2031_sign_out <= VN_sign_out( 12191 downto 12186 );
    VN2032_data_out <= VN_data_out( 12197 downto 12192 );
    VN2032_sign_out <= VN_sign_out( 12197 downto 12192 );
    VN2033_data_out <= VN_data_out( 12203 downto 12198 );
    VN2033_sign_out <= VN_sign_out( 12203 downto 12198 );
    VN2034_data_out <= VN_data_out( 12209 downto 12204 );
    VN2034_sign_out <= VN_sign_out( 12209 downto 12204 );
    VN2035_data_out <= VN_data_out( 12215 downto 12210 );
    VN2035_sign_out <= VN_sign_out( 12215 downto 12210 );
    VN2036_data_out <= VN_data_out( 12221 downto 12216 );
    VN2036_sign_out <= VN_sign_out( 12221 downto 12216 );
    VN2037_data_out <= VN_data_out( 12227 downto 12222 );
    VN2037_sign_out <= VN_sign_out( 12227 downto 12222 );
    VN2038_data_out <= VN_data_out( 12233 downto 12228 );
    VN2038_sign_out <= VN_sign_out( 12233 downto 12228 );
    VN2039_data_out <= VN_data_out( 12239 downto 12234 );
    VN2039_sign_out <= VN_sign_out( 12239 downto 12234 );
    VN2040_data_out <= VN_data_out( 12245 downto 12240 );
    VN2040_sign_out <= VN_sign_out( 12245 downto 12240 );
    VN2041_data_out <= VN_data_out( 12251 downto 12246 );
    VN2041_sign_out <= VN_sign_out( 12251 downto 12246 );
    VN2042_data_out <= VN_data_out( 12257 downto 12252 );
    VN2042_sign_out <= VN_sign_out( 12257 downto 12252 );
    VN2043_data_out <= VN_data_out( 12263 downto 12258 );
    VN2043_sign_out <= VN_sign_out( 12263 downto 12258 );
    VN2044_data_out <= VN_data_out( 12269 downto 12264 );
    VN2044_sign_out <= VN_sign_out( 12269 downto 12264 );
    VN2045_data_out <= VN_data_out( 12275 downto 12270 );
    VN2045_sign_out <= VN_sign_out( 12275 downto 12270 );
    VN2046_data_out <= VN_data_out( 12281 downto 12276 );
    VN2046_sign_out <= VN_sign_out( 12281 downto 12276 );
    VN2047_data_out <= VN_data_out( 12287 downto 12282 );
    VN2047_sign_out <= VN_sign_out( 12287 downto 12282 );


    --CN0_data_in(0) <= VN53_data_out(0);
    CN0_data_in(0) <= VN53_data_out(0);
    CN0_sign_in(0) <= VN53_sign_out(0);
    CN0_data_in(1) <= VN110_data_out(0);
    CN0_sign_in(1) <= VN110_sign_out(0);
    CN0_data_in(2) <= VN170_data_out(0);
    CN0_sign_in(2) <= VN170_sign_out(0);
    CN0_data_in(3) <= VN224_data_out(0);
    CN0_sign_in(3) <= VN224_sign_out(0);
    CN0_data_in(4) <= VN279_data_out(0);
    CN0_sign_in(4) <= VN279_sign_out(0);
    CN0_data_in(5) <= VN332_data_out(0);
    CN0_sign_in(5) <= VN332_sign_out(0);
    CN0_data_in(6) <= VN447_data_out(0);
    CN0_sign_in(6) <= VN447_sign_out(0);
    CN0_data_in(7) <= VN505_data_out(0);
    CN0_sign_in(7) <= VN505_sign_out(0);
    CN0_data_in(8) <= VN616_data_out(0);
    CN0_sign_in(8) <= VN616_sign_out(0);
    CN0_data_in(9) <= VN668_data_out(0);
    CN0_sign_in(9) <= VN668_sign_out(0);
    CN0_data_in(10) <= VN1496_data_out(0);
    CN0_sign_in(10) <= VN1496_sign_out(0);
    CN0_data_in(11) <= VN1497_data_out(0);
    CN0_sign_in(11) <= VN1497_sign_out(0);
    CN0_data_in(12) <= VN1498_data_out(0);
    CN0_sign_in(12) <= VN1498_sign_out(0);
    CN0_data_in(13) <= VN1499_data_out(0);
    CN0_sign_in(13) <= VN1499_sign_out(0);
    CN0_data_in(14) <= VN1500_data_out(0);
    CN0_sign_in(14) <= VN1500_sign_out(0);
    CN0_data_in(15) <= VN1501_data_out(0);
    CN0_sign_in(15) <= VN1501_sign_out(0);
    CN0_data_in(16) <= VN1502_data_out(0);
    CN0_sign_in(16) <= VN1502_sign_out(0);
    CN0_data_in(17) <= VN1503_data_out(0);
    CN0_sign_in(17) <= VN1503_sign_out(0);
    CN0_data_in(18) <= VN1505_data_out(0);
    CN0_sign_in(18) <= VN1505_sign_out(0);
    CN0_data_in(19) <= VN1509_data_out(0);
    CN0_sign_in(19) <= VN1509_sign_out(0);
    CN0_data_in(20) <= VN1514_data_out(0);
    CN0_sign_in(20) <= VN1514_sign_out(0);
    CN0_data_in(21) <= VN1519_data_out(0);
    CN0_sign_in(21) <= VN1519_sign_out(0);
    CN0_data_in(22) <= VN1525_data_out(0);
    CN0_sign_in(22) <= VN1525_sign_out(0);
    CN0_data_in(23) <= VN1532_data_out(0);
    CN0_sign_in(23) <= VN1532_sign_out(0);
    CN0_data_in(24) <= VN1536_data_out(0);
    CN0_sign_in(24) <= VN1536_sign_out(0);
    CN0_data_in(25) <= VN1552_data_out(0);
    CN0_sign_in(25) <= VN1552_sign_out(0);
    CN0_data_in(26) <= VN1575_data_out(0);
    CN0_sign_in(26) <= VN1575_sign_out(0);
    CN0_data_in(27) <= VN1607_data_out(0);
    CN0_sign_in(27) <= VN1607_sign_out(0);
    CN0_data_in(28) <= VN1648_data_out(0);
    CN0_sign_in(28) <= VN1648_sign_out(0);
    CN0_data_in(29) <= VN1687_data_out(0);
    CN0_sign_in(29) <= VN1687_sign_out(0);
    CN0_data_in(30) <= VN1718_data_out(0);
    CN0_sign_in(30) <= VN1718_sign_out(0);
    CN0_data_in(31) <= VN1724_data_out(0);
    CN0_sign_in(31) <= VN1724_sign_out(0);
    CN1_data_in(0) <= VN51_data_out(0);
    CN1_sign_in(0) <= VN51_sign_out(0);
    CN1_data_in(1) <= VN139_data_out(0);
    CN1_sign_in(1) <= VN139_sign_out(0);
    CN1_data_in(2) <= VN223_data_out(0);
    CN1_sign_in(2) <= VN223_sign_out(0);
    CN1_data_in(3) <= VN241_data_out(0);
    CN1_sign_in(3) <= VN241_sign_out(0);
    CN1_data_in(4) <= VN307_data_out(0);
    CN1_sign_in(4) <= VN307_sign_out(0);
    CN1_data_in(5) <= VN356_data_out(0);
    CN1_sign_in(5) <= VN356_sign_out(0);
    CN1_data_in(6) <= VN408_data_out(0);
    CN1_sign_in(6) <= VN408_sign_out(0);
    CN1_data_in(7) <= VN476_data_out(0);
    CN1_sign_in(7) <= VN476_sign_out(0);
    CN1_data_in(8) <= VN515_data_out(0);
    CN1_sign_in(8) <= VN515_sign_out(0);
    CN1_data_in(9) <= VN600_data_out(0);
    CN1_sign_in(9) <= VN600_sign_out(0);
    CN1_data_in(10) <= VN617_data_out(0);
    CN1_sign_in(10) <= VN617_sign_out(0);
    CN1_data_in(11) <= VN689_data_out(0);
    CN1_sign_in(11) <= VN689_sign_out(0);
    CN1_data_in(12) <= VN762_data_out(0);
    CN1_sign_in(12) <= VN762_sign_out(0);
    CN1_data_in(13) <= VN797_data_out(0);
    CN1_sign_in(13) <= VN797_sign_out(0);
    CN1_data_in(14) <= VN854_data_out(0);
    CN1_sign_in(14) <= VN854_sign_out(0);
    CN1_data_in(15) <= VN927_data_out(0);
    CN1_sign_in(15) <= VN927_sign_out(0);
    CN1_data_in(16) <= VN990_data_out(0);
    CN1_sign_in(16) <= VN990_sign_out(0);
    CN1_data_in(17) <= VN1023_data_out(0);
    CN1_sign_in(17) <= VN1023_sign_out(0);
    CN1_data_in(18) <= VN1059_data_out(0);
    CN1_sign_in(18) <= VN1059_sign_out(0);
    CN1_data_in(19) <= VN1077_data_out(0);
    CN1_sign_in(19) <= VN1077_sign_out(0);
    CN1_data_in(20) <= VN1138_data_out(0);
    CN1_sign_in(20) <= VN1138_sign_out(0);
    CN1_data_in(21) <= VN1200_data_out(0);
    CN1_sign_in(21) <= VN1200_sign_out(0);
    CN1_data_in(22) <= VN1292_data_out(0);
    CN1_sign_in(22) <= VN1292_sign_out(0);
    CN1_data_in(23) <= VN1442_data_out(0);
    CN1_sign_in(23) <= VN1442_sign_out(0);
    CN1_data_in(24) <= VN1488_data_out(0);
    CN1_sign_in(24) <= VN1488_sign_out(0);
    CN1_data_in(25) <= VN1522_data_out(0);
    CN1_sign_in(25) <= VN1522_sign_out(0);
    CN1_data_in(26) <= VN1535_data_out(0);
    CN1_sign_in(26) <= VN1535_sign_out(0);
    CN1_data_in(27) <= VN1550_data_out(0);
    CN1_sign_in(27) <= VN1550_sign_out(0);
    CN1_data_in(28) <= VN1585_data_out(0);
    CN1_sign_in(28) <= VN1585_sign_out(0);
    CN1_data_in(29) <= VN1681_data_out(0);
    CN1_sign_in(29) <= VN1681_sign_out(0);
    CN1_data_in(30) <= VN1994_data_out(0);
    CN1_sign_in(30) <= VN1994_sign_out(0);
    CN1_data_in(31) <= VN1996_data_out(0);
    CN1_sign_in(31) <= VN1996_sign_out(0);
    CN2_data_in(0) <= VN50_data_out(0);
    CN2_sign_in(0) <= VN50_sign_out(0);
    CN2_data_in(1) <= VN92_data_out(0);
    CN2_sign_in(1) <= VN92_sign_out(0);
    CN2_data_in(2) <= VN138_data_out(0);
    CN2_sign_in(2) <= VN138_sign_out(0);
    CN2_data_in(3) <= VN222_data_out(0);
    CN2_sign_in(3) <= VN222_sign_out(0);
    CN2_data_in(4) <= VN240_data_out(0);
    CN2_sign_in(4) <= VN240_sign_out(0);
    CN2_data_in(5) <= VN306_data_out(0);
    CN2_sign_in(5) <= VN306_sign_out(0);
    CN2_data_in(6) <= VN355_data_out(0);
    CN2_sign_in(6) <= VN355_sign_out(0);
    CN2_data_in(7) <= VN407_data_out(0);
    CN2_sign_in(7) <= VN407_sign_out(0);
    CN2_data_in(8) <= VN475_data_out(0);
    CN2_sign_in(8) <= VN475_sign_out(0);
    CN2_data_in(9) <= VN599_data_out(0);
    CN2_sign_in(9) <= VN599_sign_out(0);
    CN2_data_in(10) <= VN688_data_out(0);
    CN2_sign_in(10) <= VN688_sign_out(0);
    CN2_data_in(11) <= VN761_data_out(0);
    CN2_sign_in(11) <= VN761_sign_out(0);
    CN2_data_in(12) <= VN853_data_out(0);
    CN2_sign_in(12) <= VN853_sign_out(0);
    CN2_data_in(13) <= VN989_data_out(0);
    CN2_sign_in(13) <= VN989_sign_out(0);
    CN2_data_in(14) <= VN1003_data_out(0);
    CN2_sign_in(14) <= VN1003_sign_out(0);
    CN2_data_in(15) <= VN1022_data_out(0);
    CN2_sign_in(15) <= VN1022_sign_out(0);
    CN2_data_in(16) <= VN1076_data_out(0);
    CN2_sign_in(16) <= VN1076_sign_out(0);
    CN2_data_in(17) <= VN1137_data_out(0);
    CN2_sign_in(17) <= VN1137_sign_out(0);
    CN2_data_in(18) <= VN1199_data_out(0);
    CN2_sign_in(18) <= VN1199_sign_out(0);
    CN2_data_in(19) <= VN1291_data_out(0);
    CN2_sign_in(19) <= VN1291_sign_out(0);
    CN2_data_in(20) <= VN1441_data_out(0);
    CN2_sign_in(20) <= VN1441_sign_out(0);
    CN2_data_in(21) <= VN1521_data_out(0);
    CN2_sign_in(21) <= VN1521_sign_out(0);
    CN2_data_in(22) <= VN1534_data_out(0);
    CN2_sign_in(22) <= VN1534_sign_out(0);
    CN2_data_in(23) <= VN1549_data_out(0);
    CN2_sign_in(23) <= VN1549_sign_out(0);
    CN2_data_in(24) <= VN1584_data_out(0);
    CN2_sign_in(24) <= VN1584_sign_out(0);
    CN2_data_in(25) <= VN1707_data_out(0);
    CN2_sign_in(25) <= VN1707_sign_out(0);
    CN2_data_in(26) <= VN1808_data_out(0);
    CN2_sign_in(26) <= VN1808_sign_out(0);
    CN2_data_in(27) <= VN1837_data_out(0);
    CN2_sign_in(27) <= VN1837_sign_out(0);
    CN2_data_in(28) <= VN1904_data_out(0);
    CN2_sign_in(28) <= VN1904_sign_out(0);
    CN2_data_in(29) <= VN1948_data_out(0);
    CN2_sign_in(29) <= VN1948_sign_out(0);
    CN2_data_in(30) <= VN2003_data_out(0);
    CN2_sign_in(30) <= VN2003_sign_out(0);
    CN2_data_in(31) <= VN2007_data_out(0);
    CN2_sign_in(31) <= VN2007_sign_out(0);
    CN3_data_in(0) <= VN91_data_out(0);
    CN3_sign_in(0) <= VN91_sign_out(0);
    CN3_data_in(1) <= VN137_data_out(0);
    CN3_sign_in(1) <= VN137_sign_out(0);
    CN3_data_in(2) <= VN221_data_out(0);
    CN3_sign_in(2) <= VN221_sign_out(0);
    CN3_data_in(3) <= VN239_data_out(0);
    CN3_sign_in(3) <= VN239_sign_out(0);
    CN3_data_in(4) <= VN305_data_out(0);
    CN3_sign_in(4) <= VN305_sign_out(0);
    CN3_data_in(5) <= VN474_data_out(0);
    CN3_sign_in(5) <= VN474_sign_out(0);
    CN3_data_in(6) <= VN514_data_out(0);
    CN3_sign_in(6) <= VN514_sign_out(0);
    CN3_data_in(7) <= VN598_data_out(0);
    CN3_sign_in(7) <= VN598_sign_out(0);
    CN3_data_in(8) <= VN687_data_out(0);
    CN3_sign_in(8) <= VN687_sign_out(0);
    CN3_data_in(9) <= VN760_data_out(0);
    CN3_sign_in(9) <= VN760_sign_out(0);
    CN3_data_in(10) <= VN796_data_out(0);
    CN3_sign_in(10) <= VN796_sign_out(0);
    CN3_data_in(11) <= VN852_data_out(0);
    CN3_sign_in(11) <= VN852_sign_out(0);
    CN3_data_in(12) <= VN926_data_out(0);
    CN3_sign_in(12) <= VN926_sign_out(0);
    CN3_data_in(13) <= VN988_data_out(0);
    CN3_sign_in(13) <= VN988_sign_out(0);
    CN3_data_in(14) <= VN1021_data_out(0);
    CN3_sign_in(14) <= VN1021_sign_out(0);
    CN3_data_in(15) <= VN1075_data_out(0);
    CN3_sign_in(15) <= VN1075_sign_out(0);
    CN3_data_in(16) <= VN1136_data_out(0);
    CN3_sign_in(16) <= VN1136_sign_out(0);
    CN3_data_in(17) <= VN1290_data_out(0);
    CN3_sign_in(17) <= VN1290_sign_out(0);
    CN3_data_in(18) <= VN1440_data_out(0);
    CN3_sign_in(18) <= VN1440_sign_out(0);
    CN3_data_in(19) <= VN1520_data_out(0);
    CN3_sign_in(19) <= VN1520_sign_out(0);
    CN3_data_in(20) <= VN1533_data_out(0);
    CN3_sign_in(20) <= VN1533_sign_out(0);
    CN3_data_in(21) <= VN1548_data_out(0);
    CN3_sign_in(21) <= VN1548_sign_out(0);
    CN3_data_in(22) <= VN1647_data_out(0);
    CN3_sign_in(22) <= VN1647_sign_out(0);
    CN3_data_in(23) <= VN1680_data_out(0);
    CN3_sign_in(23) <= VN1680_sign_out(0);
    CN3_data_in(24) <= VN1801_data_out(0);
    CN3_sign_in(24) <= VN1801_sign_out(0);
    CN3_data_in(25) <= VN1824_data_out(0);
    CN3_sign_in(25) <= VN1824_sign_out(0);
    CN3_data_in(26) <= VN1833_data_out(0);
    CN3_sign_in(26) <= VN1833_sign_out(0);
    CN3_data_in(27) <= VN1845_data_out(0);
    CN3_sign_in(27) <= VN1845_sign_out(0);
    CN3_data_in(28) <= VN1850_data_out(0);
    CN3_sign_in(28) <= VN1850_sign_out(0);
    CN3_data_in(29) <= VN1919_data_out(0);
    CN3_sign_in(29) <= VN1919_sign_out(0);
    CN3_data_in(30) <= VN1940_data_out(0);
    CN3_sign_in(30) <= VN1940_sign_out(0);
    CN3_data_in(31) <= VN1942_data_out(0);
    CN3_sign_in(31) <= VN1942_sign_out(0);
    CN4_data_in(0) <= VN49_data_out(0);
    CN4_sign_in(0) <= VN49_sign_out(0);
    CN4_data_in(1) <= VN90_data_out(0);
    CN4_sign_in(1) <= VN90_sign_out(0);
    CN4_data_in(2) <= VN220_data_out(0);
    CN4_sign_in(2) <= VN220_sign_out(0);
    CN4_data_in(3) <= VN238_data_out(0);
    CN4_sign_in(3) <= VN238_sign_out(0);
    CN4_data_in(4) <= VN304_data_out(0);
    CN4_sign_in(4) <= VN304_sign_out(0);
    CN4_data_in(5) <= VN354_data_out(0);
    CN4_sign_in(5) <= VN354_sign_out(0);
    CN4_data_in(6) <= VN406_data_out(0);
    CN4_sign_in(6) <= VN406_sign_out(0);
    CN4_data_in(7) <= VN473_data_out(0);
    CN4_sign_in(7) <= VN473_sign_out(0);
    CN4_data_in(8) <= VN513_data_out(0);
    CN4_sign_in(8) <= VN513_sign_out(0);
    CN4_data_in(9) <= VN597_data_out(0);
    CN4_sign_in(9) <= VN597_sign_out(0);
    CN4_data_in(10) <= VN667_data_out(0);
    CN4_sign_in(10) <= VN667_sign_out(0);
    CN4_data_in(11) <= VN686_data_out(0);
    CN4_sign_in(11) <= VN686_sign_out(0);
    CN4_data_in(12) <= VN759_data_out(0);
    CN4_sign_in(12) <= VN759_sign_out(0);
    CN4_data_in(13) <= VN795_data_out(0);
    CN4_sign_in(13) <= VN795_sign_out(0);
    CN4_data_in(14) <= VN851_data_out(0);
    CN4_sign_in(14) <= VN851_sign_out(0);
    CN4_data_in(15) <= VN887_data_out(0);
    CN4_sign_in(15) <= VN887_sign_out(0);
    CN4_data_in(16) <= VN925_data_out(0);
    CN4_sign_in(16) <= VN925_sign_out(0);
    CN4_data_in(17) <= VN987_data_out(0);
    CN4_sign_in(17) <= VN987_sign_out(0);
    CN4_data_in(18) <= VN1074_data_out(0);
    CN4_sign_in(18) <= VN1074_sign_out(0);
    CN4_data_in(19) <= VN1135_data_out(0);
    CN4_sign_in(19) <= VN1135_sign_out(0);
    CN4_data_in(20) <= VN1198_data_out(0);
    CN4_sign_in(20) <= VN1198_sign_out(0);
    CN4_data_in(21) <= VN1289_data_out(0);
    CN4_sign_in(21) <= VN1289_sign_out(0);
    CN4_data_in(22) <= VN1583_data_out(0);
    CN4_sign_in(22) <= VN1583_sign_out(0);
    CN4_data_in(23) <= VN1646_data_out(0);
    CN4_sign_in(23) <= VN1646_sign_out(0);
    CN4_data_in(24) <= VN1679_data_out(0);
    CN4_sign_in(24) <= VN1679_sign_out(0);
    CN4_data_in(25) <= VN1747_data_out(0);
    CN4_sign_in(25) <= VN1747_sign_out(0);
    CN4_data_in(26) <= VN1892_data_out(0);
    CN4_sign_in(26) <= VN1892_sign_out(0);
    CN4_data_in(27) <= VN1901_data_out(0);
    CN4_sign_in(27) <= VN1901_sign_out(0);
    CN4_data_in(28) <= VN1907_data_out(0);
    CN4_sign_in(28) <= VN1907_sign_out(0);
    CN4_data_in(29) <= VN1944_data_out(0);
    CN4_sign_in(29) <= VN1944_sign_out(0);
    CN4_data_in(30) <= VN1977_data_out(0);
    CN4_sign_in(30) <= VN1977_sign_out(0);
    CN4_data_in(31) <= VN1978_data_out(0);
    CN4_sign_in(31) <= VN1978_sign_out(0);
    CN5_data_in(0) <= VN48_data_out(0);
    CN5_sign_in(0) <= VN48_sign_out(0);
    CN5_data_in(1) <= VN89_data_out(0);
    CN5_sign_in(1) <= VN89_sign_out(0);
    CN5_data_in(2) <= VN136_data_out(0);
    CN5_sign_in(2) <= VN136_sign_out(0);
    CN5_data_in(3) <= VN219_data_out(0);
    CN5_sign_in(3) <= VN219_sign_out(0);
    CN5_data_in(4) <= VN237_data_out(0);
    CN5_sign_in(4) <= VN237_sign_out(0);
    CN5_data_in(5) <= VN303_data_out(0);
    CN5_sign_in(5) <= VN303_sign_out(0);
    CN5_data_in(6) <= VN353_data_out(0);
    CN5_sign_in(6) <= VN353_sign_out(0);
    CN5_data_in(7) <= VN405_data_out(0);
    CN5_sign_in(7) <= VN405_sign_out(0);
    CN5_data_in(8) <= VN472_data_out(0);
    CN5_sign_in(8) <= VN472_sign_out(0);
    CN5_data_in(9) <= VN512_data_out(0);
    CN5_sign_in(9) <= VN512_sign_out(0);
    CN5_data_in(10) <= VN596_data_out(0);
    CN5_sign_in(10) <= VN596_sign_out(0);
    CN5_data_in(11) <= VN666_data_out(0);
    CN5_sign_in(11) <= VN666_sign_out(0);
    CN5_data_in(12) <= VN685_data_out(0);
    CN5_sign_in(12) <= VN685_sign_out(0);
    CN5_data_in(13) <= VN758_data_out(0);
    CN5_sign_in(13) <= VN758_sign_out(0);
    CN5_data_in(14) <= VN794_data_out(0);
    CN5_sign_in(14) <= VN794_sign_out(0);
    CN5_data_in(15) <= VN830_data_out(0);
    CN5_sign_in(15) <= VN830_sign_out(0);
    CN5_data_in(16) <= VN850_data_out(0);
    CN5_sign_in(16) <= VN850_sign_out(0);
    CN5_data_in(17) <= VN924_data_out(0);
    CN5_sign_in(17) <= VN924_sign_out(0);
    CN5_data_in(18) <= VN986_data_out(0);
    CN5_sign_in(18) <= VN986_sign_out(0);
    CN5_data_in(19) <= VN1020_data_out(0);
    CN5_sign_in(19) <= VN1020_sign_out(0);
    CN5_data_in(20) <= VN1073_data_out(0);
    CN5_sign_in(20) <= VN1073_sign_out(0);
    CN5_data_in(21) <= VN1134_data_out(0);
    CN5_sign_in(21) <= VN1134_sign_out(0);
    CN5_data_in(22) <= VN1197_data_out(0);
    CN5_sign_in(22) <= VN1197_sign_out(0);
    CN5_data_in(23) <= VN1275_data_out(0);
    CN5_sign_in(23) <= VN1275_sign_out(0);
    CN5_data_in(24) <= VN1288_data_out(0);
    CN5_sign_in(24) <= VN1288_sign_out(0);
    CN5_data_in(25) <= VN1383_data_out(0);
    CN5_sign_in(25) <= VN1383_sign_out(0);
    CN5_data_in(26) <= VN1439_data_out(0);
    CN5_sign_in(26) <= VN1439_sign_out(0);
    CN5_data_in(27) <= VN1547_data_out(0);
    CN5_sign_in(27) <= VN1547_sign_out(0);
    CN5_data_in(28) <= VN1582_data_out(0);
    CN5_sign_in(28) <= VN1582_sign_out(0);
    CN5_data_in(29) <= VN1645_data_out(0);
    CN5_sign_in(29) <= VN1645_sign_out(0);
    CN5_data_in(30) <= VN1678_data_out(0);
    CN5_sign_in(30) <= VN1678_sign_out(0);
    CN5_data_in(31) <= VN1725_data_out(0);
    CN5_sign_in(31) <= VN1725_sign_out(0);
    CN6_data_in(0) <= VN47_data_out(0);
    CN6_sign_in(0) <= VN47_sign_out(0);
    CN6_data_in(1) <= VN88_data_out(0);
    CN6_sign_in(1) <= VN88_sign_out(0);
    CN6_data_in(2) <= VN135_data_out(0);
    CN6_sign_in(2) <= VN135_sign_out(0);
    CN6_data_in(3) <= VN218_data_out(0);
    CN6_sign_in(3) <= VN218_sign_out(0);
    CN6_data_in(4) <= VN236_data_out(0);
    CN6_sign_in(4) <= VN236_sign_out(0);
    CN6_data_in(5) <= VN302_data_out(0);
    CN6_sign_in(5) <= VN302_sign_out(0);
    CN6_data_in(6) <= VN352_data_out(0);
    CN6_sign_in(6) <= VN352_sign_out(0);
    CN6_data_in(7) <= VN404_data_out(0);
    CN6_sign_in(7) <= VN404_sign_out(0);
    CN6_data_in(8) <= VN471_data_out(0);
    CN6_sign_in(8) <= VN471_sign_out(0);
    CN6_data_in(9) <= VN511_data_out(0);
    CN6_sign_in(9) <= VN511_sign_out(0);
    CN6_data_in(10) <= VN595_data_out(0);
    CN6_sign_in(10) <= VN595_sign_out(0);
    CN6_data_in(11) <= VN665_data_out(0);
    CN6_sign_in(11) <= VN665_sign_out(0);
    CN6_data_in(12) <= VN684_data_out(0);
    CN6_sign_in(12) <= VN684_sign_out(0);
    CN6_data_in(13) <= VN757_data_out(0);
    CN6_sign_in(13) <= VN757_sign_out(0);
    CN6_data_in(14) <= VN777_data_out(0);
    CN6_sign_in(14) <= VN777_sign_out(0);
    CN6_data_in(15) <= VN793_data_out(0);
    CN6_sign_in(15) <= VN793_sign_out(0);
    CN6_data_in(16) <= VN849_data_out(0);
    CN6_sign_in(16) <= VN849_sign_out(0);
    CN6_data_in(17) <= VN923_data_out(0);
    CN6_sign_in(17) <= VN923_sign_out(0);
    CN6_data_in(18) <= VN985_data_out(0);
    CN6_sign_in(18) <= VN985_sign_out(0);
    CN6_data_in(19) <= VN1019_data_out(0);
    CN6_sign_in(19) <= VN1019_sign_out(0);
    CN6_data_in(20) <= VN1072_data_out(0);
    CN6_sign_in(20) <= VN1072_sign_out(0);
    CN6_data_in(21) <= VN1133_data_out(0);
    CN6_sign_in(21) <= VN1133_sign_out(0);
    CN6_data_in(22) <= VN1196_data_out(0);
    CN6_sign_in(22) <= VN1196_sign_out(0);
    CN6_data_in(23) <= VN1274_data_out(0);
    CN6_sign_in(23) <= VN1274_sign_out(0);
    CN6_data_in(24) <= VN1287_data_out(0);
    CN6_sign_in(24) <= VN1287_sign_out(0);
    CN6_data_in(25) <= VN1382_data_out(0);
    CN6_sign_in(25) <= VN1382_sign_out(0);
    CN6_data_in(26) <= VN1438_data_out(0);
    CN6_sign_in(26) <= VN1438_sign_out(0);
    CN6_data_in(27) <= VN1546_data_out(0);
    CN6_sign_in(27) <= VN1546_sign_out(0);
    CN6_data_in(28) <= VN1581_data_out(0);
    CN6_sign_in(28) <= VN1581_sign_out(0);
    CN6_data_in(29) <= VN1644_data_out(0);
    CN6_sign_in(29) <= VN1644_sign_out(0);
    CN6_data_in(30) <= VN1706_data_out(0);
    CN6_sign_in(30) <= VN1706_sign_out(0);
    CN6_data_in(31) <= VN1726_data_out(0);
    CN6_sign_in(31) <= VN1726_sign_out(0);
    CN7_data_in(0) <= VN46_data_out(0);
    CN7_sign_in(0) <= VN46_sign_out(0);
    CN7_data_in(1) <= VN87_data_out(0);
    CN7_sign_in(1) <= VN87_sign_out(0);
    CN7_data_in(2) <= VN134_data_out(0);
    CN7_sign_in(2) <= VN134_sign_out(0);
    CN7_data_in(3) <= VN217_data_out(0);
    CN7_sign_in(3) <= VN217_sign_out(0);
    CN7_data_in(4) <= VN235_data_out(0);
    CN7_sign_in(4) <= VN235_sign_out(0);
    CN7_data_in(5) <= VN301_data_out(0);
    CN7_sign_in(5) <= VN301_sign_out(0);
    CN7_data_in(6) <= VN351_data_out(0);
    CN7_sign_in(6) <= VN351_sign_out(0);
    CN7_data_in(7) <= VN403_data_out(0);
    CN7_sign_in(7) <= VN403_sign_out(0);
    CN7_data_in(8) <= VN470_data_out(0);
    CN7_sign_in(8) <= VN470_sign_out(0);
    CN7_data_in(9) <= VN510_data_out(0);
    CN7_sign_in(9) <= VN510_sign_out(0);
    CN7_data_in(10) <= VN594_data_out(0);
    CN7_sign_in(10) <= VN594_sign_out(0);
    CN7_data_in(11) <= VN664_data_out(0);
    CN7_sign_in(11) <= VN664_sign_out(0);
    CN7_data_in(12) <= VN683_data_out(0);
    CN7_sign_in(12) <= VN683_sign_out(0);
    CN7_data_in(13) <= VN722_data_out(0);
    CN7_sign_in(13) <= VN722_sign_out(0);
    CN7_data_in(14) <= VN756_data_out(0);
    CN7_sign_in(14) <= VN756_sign_out(0);
    CN7_data_in(15) <= VN792_data_out(0);
    CN7_sign_in(15) <= VN792_sign_out(0);
    CN7_data_in(16) <= VN848_data_out(0);
    CN7_sign_in(16) <= VN848_sign_out(0);
    CN7_data_in(17) <= VN922_data_out(0);
    CN7_sign_in(17) <= VN922_sign_out(0);
    CN7_data_in(18) <= VN984_data_out(0);
    CN7_sign_in(18) <= VN984_sign_out(0);
    CN7_data_in(19) <= VN1018_data_out(0);
    CN7_sign_in(19) <= VN1018_sign_out(0);
    CN7_data_in(20) <= VN1071_data_out(0);
    CN7_sign_in(20) <= VN1071_sign_out(0);
    CN7_data_in(21) <= VN1132_data_out(0);
    CN7_sign_in(21) <= VN1132_sign_out(0);
    CN7_data_in(22) <= VN1195_data_out(0);
    CN7_sign_in(22) <= VN1195_sign_out(0);
    CN7_data_in(23) <= VN1273_data_out(0);
    CN7_sign_in(23) <= VN1273_sign_out(0);
    CN7_data_in(24) <= VN1286_data_out(0);
    CN7_sign_in(24) <= VN1286_sign_out(0);
    CN7_data_in(25) <= VN1381_data_out(0);
    CN7_sign_in(25) <= VN1381_sign_out(0);
    CN7_data_in(26) <= VN1437_data_out(0);
    CN7_sign_in(26) <= VN1437_sign_out(0);
    CN7_data_in(27) <= VN1545_data_out(0);
    CN7_sign_in(27) <= VN1545_sign_out(0);
    CN7_data_in(28) <= VN1580_data_out(0);
    CN7_sign_in(28) <= VN1580_sign_out(0);
    CN7_data_in(29) <= VN1677_data_out(0);
    CN7_sign_in(29) <= VN1677_sign_out(0);
    CN7_data_in(30) <= VN1705_data_out(0);
    CN7_sign_in(30) <= VN1705_sign_out(0);
    CN7_data_in(31) <= VN1727_data_out(0);
    CN7_sign_in(31) <= VN1727_sign_out(0);
    CN8_data_in(0) <= VN45_data_out(0);
    CN8_sign_in(0) <= VN45_sign_out(0);
    CN8_data_in(1) <= VN133_data_out(0);
    CN8_sign_in(1) <= VN133_sign_out(0);
    CN8_data_in(2) <= VN216_data_out(0);
    CN8_sign_in(2) <= VN216_sign_out(0);
    CN8_data_in(3) <= VN402_data_out(0);
    CN8_sign_in(3) <= VN402_sign_out(0);
    CN8_data_in(4) <= VN469_data_out(0);
    CN8_sign_in(4) <= VN469_sign_out(0);
    CN8_data_in(5) <= VN593_data_out(0);
    CN8_sign_in(5) <= VN593_sign_out(0);
    CN8_data_in(6) <= VN682_data_out(0);
    CN8_sign_in(6) <= VN682_sign_out(0);
    CN8_data_in(7) <= VN755_data_out(0);
    CN8_sign_in(7) <= VN755_sign_out(0);
    CN8_data_in(8) <= VN847_data_out(0);
    CN8_sign_in(8) <= VN847_sign_out(0);
    CN8_data_in(9) <= VN983_data_out(0);
    CN8_sign_in(9) <= VN983_sign_out(0);
    CN8_data_in(10) <= VN1017_data_out(0);
    CN8_sign_in(10) <= VN1017_sign_out(0);
    CN8_data_in(11) <= VN1070_data_out(0);
    CN8_sign_in(11) <= VN1070_sign_out(0);
    CN8_data_in(12) <= VN1131_data_out(0);
    CN8_sign_in(12) <= VN1131_sign_out(0);
    CN8_data_in(13) <= VN1194_data_out(0);
    CN8_sign_in(13) <= VN1194_sign_out(0);
    CN8_data_in(14) <= VN1272_data_out(0);
    CN8_sign_in(14) <= VN1272_sign_out(0);
    CN8_data_in(15) <= VN1380_data_out(0);
    CN8_sign_in(15) <= VN1380_sign_out(0);
    CN8_data_in(16) <= VN1436_data_out(0);
    CN8_sign_in(16) <= VN1436_sign_out(0);
    CN8_data_in(17) <= VN1544_data_out(0);
    CN8_sign_in(17) <= VN1544_sign_out(0);
    CN8_data_in(18) <= VN1643_data_out(0);
    CN8_sign_in(18) <= VN1643_sign_out(0);
    CN8_data_in(19) <= VN1676_data_out(0);
    CN8_sign_in(19) <= VN1676_sign_out(0);
    CN8_data_in(20) <= VN1788_data_out(0);
    CN8_sign_in(20) <= VN1788_sign_out(0);
    CN8_data_in(21) <= VN1792_data_out(0);
    CN8_sign_in(21) <= VN1792_sign_out(0);
    CN8_data_in(22) <= VN1859_data_out(0);
    CN8_sign_in(22) <= VN1859_sign_out(0);
    CN8_data_in(23) <= VN1886_data_out(0);
    CN8_sign_in(23) <= VN1886_sign_out(0);
    CN8_data_in(24) <= VN1891_data_out(0);
    CN8_sign_in(24) <= VN1891_sign_out(0);
    CN8_data_in(25) <= VN1902_data_out(0);
    CN8_sign_in(25) <= VN1902_sign_out(0);
    CN8_data_in(26) <= VN1924_data_out(0);
    CN8_sign_in(26) <= VN1924_sign_out(0);
    CN8_data_in(27) <= VN1965_data_out(0);
    CN8_sign_in(27) <= VN1965_sign_out(0);
    CN8_data_in(28) <= VN1997_data_out(0);
    CN8_sign_in(28) <= VN1997_sign_out(0);
    CN8_data_in(29) <= VN2019_data_out(0);
    CN8_sign_in(29) <= VN2019_sign_out(0);
    CN8_data_in(30) <= VN2037_data_out(0);
    CN8_sign_in(30) <= VN2037_sign_out(0);
    CN8_data_in(31) <= VN2038_data_out(0);
    CN8_sign_in(31) <= VN2038_sign_out(0);
    CN9_data_in(0) <= VN44_data_out(0);
    CN9_sign_in(0) <= VN44_sign_out(0);
    CN9_data_in(1) <= VN86_data_out(0);
    CN9_sign_in(1) <= VN86_sign_out(0);
    CN9_data_in(2) <= VN132_data_out(0);
    CN9_sign_in(2) <= VN132_sign_out(0);
    CN9_data_in(3) <= VN215_data_out(0);
    CN9_sign_in(3) <= VN215_sign_out(0);
    CN9_data_in(4) <= VN234_data_out(0);
    CN9_sign_in(4) <= VN234_sign_out(0);
    CN9_data_in(5) <= VN300_data_out(0);
    CN9_sign_in(5) <= VN300_sign_out(0);
    CN9_data_in(6) <= VN350_data_out(0);
    CN9_sign_in(6) <= VN350_sign_out(0);
    CN9_data_in(7) <= VN391_data_out(0);
    CN9_sign_in(7) <= VN391_sign_out(0);
    CN9_data_in(8) <= VN401_data_out(0);
    CN9_sign_in(8) <= VN401_sign_out(0);
    CN9_data_in(9) <= VN468_data_out(0);
    CN9_sign_in(9) <= VN468_sign_out(0);
    CN9_data_in(10) <= VN509_data_out(0);
    CN9_sign_in(10) <= VN509_sign_out(0);
    CN9_data_in(11) <= VN592_data_out(0);
    CN9_sign_in(11) <= VN592_sign_out(0);
    CN9_data_in(12) <= VN663_data_out(0);
    CN9_sign_in(12) <= VN663_sign_out(0);
    CN9_data_in(13) <= VN681_data_out(0);
    CN9_sign_in(13) <= VN681_sign_out(0);
    CN9_data_in(14) <= VN754_data_out(0);
    CN9_sign_in(14) <= VN754_sign_out(0);
    CN9_data_in(15) <= VN791_data_out(0);
    CN9_sign_in(15) <= VN791_sign_out(0);
    CN9_data_in(16) <= VN846_data_out(0);
    CN9_sign_in(16) <= VN846_sign_out(0);
    CN9_data_in(17) <= VN921_data_out(0);
    CN9_sign_in(17) <= VN921_sign_out(0);
    CN9_data_in(18) <= VN982_data_out(0);
    CN9_sign_in(18) <= VN982_sign_out(0);
    CN9_data_in(19) <= VN1016_data_out(0);
    CN9_sign_in(19) <= VN1016_sign_out(0);
    CN9_data_in(20) <= VN1069_data_out(0);
    CN9_sign_in(20) <= VN1069_sign_out(0);
    CN9_data_in(21) <= VN1130_data_out(0);
    CN9_sign_in(21) <= VN1130_sign_out(0);
    CN9_data_in(22) <= VN1193_data_out(0);
    CN9_sign_in(22) <= VN1193_sign_out(0);
    CN9_data_in(23) <= VN1271_data_out(0);
    CN9_sign_in(23) <= VN1271_sign_out(0);
    CN9_data_in(24) <= VN1285_data_out(0);
    CN9_sign_in(24) <= VN1285_sign_out(0);
    CN9_data_in(25) <= VN1379_data_out(0);
    CN9_sign_in(25) <= VN1379_sign_out(0);
    CN9_data_in(26) <= VN1435_data_out(0);
    CN9_sign_in(26) <= VN1435_sign_out(0);
    CN9_data_in(27) <= VN1543_data_out(0);
    CN9_sign_in(27) <= VN1543_sign_out(0);
    CN9_data_in(28) <= VN1579_data_out(0);
    CN9_sign_in(28) <= VN1579_sign_out(0);
    CN9_data_in(29) <= VN1642_data_out(0);
    CN9_sign_in(29) <= VN1642_sign_out(0);
    CN9_data_in(30) <= VN1675_data_out(0);
    CN9_sign_in(30) <= VN1675_sign_out(0);
    CN9_data_in(31) <= VN1728_data_out(0);
    CN9_sign_in(31) <= VN1728_sign_out(0);
    CN10_data_in(0) <= VN43_data_out(0);
    CN10_sign_in(0) <= VN43_sign_out(0);
    CN10_data_in(1) <= VN85_data_out(0);
    CN10_sign_in(1) <= VN85_sign_out(0);
    CN10_data_in(2) <= VN131_data_out(0);
    CN10_sign_in(2) <= VN131_sign_out(0);
    CN10_data_in(3) <= VN233_data_out(0);
    CN10_sign_in(3) <= VN233_sign_out(0);
    CN10_data_in(4) <= VN349_data_out(0);
    CN10_sign_in(4) <= VN349_sign_out(0);
    CN10_data_in(5) <= VN467_data_out(0);
    CN10_sign_in(5) <= VN467_sign_out(0);
    CN10_data_in(6) <= VN508_data_out(0);
    CN10_sign_in(6) <= VN508_sign_out(0);
    CN10_data_in(7) <= VN662_data_out(0);
    CN10_sign_in(7) <= VN662_sign_out(0);
    CN10_data_in(8) <= VN753_data_out(0);
    CN10_sign_in(8) <= VN753_sign_out(0);
    CN10_data_in(9) <= VN790_data_out(0);
    CN10_sign_in(9) <= VN790_sign_out(0);
    CN10_data_in(10) <= VN845_data_out(0);
    CN10_sign_in(10) <= VN845_sign_out(0);
    CN10_data_in(11) <= VN920_data_out(0);
    CN10_sign_in(11) <= VN920_sign_out(0);
    CN10_data_in(12) <= VN981_data_out(0);
    CN10_sign_in(12) <= VN981_sign_out(0);
    CN10_data_in(13) <= VN1015_data_out(0);
    CN10_sign_in(13) <= VN1015_sign_out(0);
    CN10_data_in(14) <= VN1270_data_out(0);
    CN10_sign_in(14) <= VN1270_sign_out(0);
    CN10_data_in(15) <= VN1378_data_out(0);
    CN10_sign_in(15) <= VN1378_sign_out(0);
    CN10_data_in(16) <= VN1455_data_out(0);
    CN10_sign_in(16) <= VN1455_sign_out(0);
    CN10_data_in(17) <= VN1542_data_out(0);
    CN10_sign_in(17) <= VN1542_sign_out(0);
    CN10_data_in(18) <= VN1578_data_out(0);
    CN10_sign_in(18) <= VN1578_sign_out(0);
    CN10_data_in(19) <= VN1641_data_out(0);
    CN10_sign_in(19) <= VN1641_sign_out(0);
    CN10_data_in(20) <= VN1674_data_out(0);
    CN10_sign_in(20) <= VN1674_sign_out(0);
    CN10_data_in(21) <= VN1704_data_out(0);
    CN10_sign_in(21) <= VN1704_sign_out(0);
    CN10_data_in(22) <= VN1830_data_out(0);
    CN10_sign_in(22) <= VN1830_sign_out(0);
    CN10_data_in(23) <= VN1895_data_out(0);
    CN10_sign_in(23) <= VN1895_sign_out(0);
    CN10_data_in(24) <= VN1918_data_out(0);
    CN10_sign_in(24) <= VN1918_sign_out(0);
    CN10_data_in(25) <= VN1971_data_out(0);
    CN10_sign_in(25) <= VN1971_sign_out(0);
    CN10_data_in(26) <= VN1981_data_out(0);
    CN10_sign_in(26) <= VN1981_sign_out(0);
    CN10_data_in(27) <= VN1982_data_out(0);
    CN10_sign_in(27) <= VN1982_sign_out(0);
    CN10_data_in(28) <= VN1993_data_out(0);
    CN10_sign_in(28) <= VN1993_sign_out(0);
    CN10_data_in(29) <= VN2009_data_out(0);
    CN10_sign_in(29) <= VN2009_sign_out(0);
    CN10_data_in(30) <= VN2013_data_out(0);
    CN10_sign_in(30) <= VN2013_sign_out(0);
    CN10_data_in(31) <= VN2014_data_out(0);
    CN10_sign_in(31) <= VN2014_sign_out(0);
    CN11_data_in(0) <= VN42_data_out(0);
    CN11_sign_in(0) <= VN42_sign_out(0);
    CN11_data_in(1) <= VN84_data_out(0);
    CN11_sign_in(1) <= VN84_sign_out(0);
    CN11_data_in(2) <= VN130_data_out(0);
    CN11_sign_in(2) <= VN130_sign_out(0);
    CN11_data_in(3) <= VN214_data_out(0);
    CN11_sign_in(3) <= VN214_sign_out(0);
    CN11_data_in(4) <= VN232_data_out(0);
    CN11_sign_in(4) <= VN232_sign_out(0);
    CN11_data_in(5) <= VN348_data_out(0);
    CN11_sign_in(5) <= VN348_sign_out(0);
    CN11_data_in(6) <= VN400_data_out(0);
    CN11_sign_in(6) <= VN400_sign_out(0);
    CN11_data_in(7) <= VN591_data_out(0);
    CN11_sign_in(7) <= VN591_sign_out(0);
    CN11_data_in(8) <= VN661_data_out(0);
    CN11_sign_in(8) <= VN661_sign_out(0);
    CN11_data_in(9) <= VN680_data_out(0);
    CN11_sign_in(9) <= VN680_sign_out(0);
    CN11_data_in(10) <= VN752_data_out(0);
    CN11_sign_in(10) <= VN752_sign_out(0);
    CN11_data_in(11) <= VN789_data_out(0);
    CN11_sign_in(11) <= VN789_sign_out(0);
    CN11_data_in(12) <= VN844_data_out(0);
    CN11_sign_in(12) <= VN844_sign_out(0);
    CN11_data_in(13) <= VN919_data_out(0);
    CN11_sign_in(13) <= VN919_sign_out(0);
    CN11_data_in(14) <= VN1014_data_out(0);
    CN11_sign_in(14) <= VN1014_sign_out(0);
    CN11_data_in(15) <= VN1068_data_out(0);
    CN11_sign_in(15) <= VN1068_sign_out(0);
    CN11_data_in(16) <= VN1129_data_out(0);
    CN11_sign_in(16) <= VN1129_sign_out(0);
    CN11_data_in(17) <= VN1269_data_out(0);
    CN11_sign_in(17) <= VN1269_sign_out(0);
    CN11_data_in(18) <= VN1434_data_out(0);
    CN11_sign_in(18) <= VN1434_sign_out(0);
    CN11_data_in(19) <= VN1454_data_out(0);
    CN11_sign_in(19) <= VN1454_sign_out(0);
    CN11_data_in(20) <= VN1541_data_out(0);
    CN11_sign_in(20) <= VN1541_sign_out(0);
    CN11_data_in(21) <= VN1577_data_out(0);
    CN11_sign_in(21) <= VN1577_sign_out(0);
    CN11_data_in(22) <= VN1640_data_out(0);
    CN11_sign_in(22) <= VN1640_sign_out(0);
    CN11_data_in(23) <= VN1673_data_out(0);
    CN11_sign_in(23) <= VN1673_sign_out(0);
    CN11_data_in(24) <= VN1764_data_out(0);
    CN11_sign_in(24) <= VN1764_sign_out(0);
    CN11_data_in(25) <= VN1829_data_out(0);
    CN11_sign_in(25) <= VN1829_sign_out(0);
    CN11_data_in(26) <= VN1843_data_out(0);
    CN11_sign_in(26) <= VN1843_sign_out(0);
    CN11_data_in(27) <= VN1860_data_out(0);
    CN11_sign_in(27) <= VN1860_sign_out(0);
    CN11_data_in(28) <= VN1867_data_out(0);
    CN11_sign_in(28) <= VN1867_sign_out(0);
    CN11_data_in(29) <= VN1914_data_out(0);
    CN11_sign_in(29) <= VN1914_sign_out(0);
    CN11_data_in(30) <= VN1946_data_out(0);
    CN11_sign_in(30) <= VN1946_sign_out(0);
    CN11_data_in(31) <= VN1951_data_out(0);
    CN11_sign_in(31) <= VN1951_sign_out(0);
    CN12_data_in(0) <= VN41_data_out(0);
    CN12_sign_in(0) <= VN41_sign_out(0);
    CN12_data_in(1) <= VN83_data_out(0);
    CN12_sign_in(1) <= VN83_sign_out(0);
    CN12_data_in(2) <= VN129_data_out(0);
    CN12_sign_in(2) <= VN129_sign_out(0);
    CN12_data_in(3) <= VN213_data_out(0);
    CN12_sign_in(3) <= VN213_sign_out(0);
    CN12_data_in(4) <= VN231_data_out(0);
    CN12_sign_in(4) <= VN231_sign_out(0);
    CN12_data_in(5) <= VN299_data_out(0);
    CN12_sign_in(5) <= VN299_sign_out(0);
    CN12_data_in(6) <= VN347_data_out(0);
    CN12_sign_in(6) <= VN347_sign_out(0);
    CN12_data_in(7) <= VN399_data_out(0);
    CN12_sign_in(7) <= VN399_sign_out(0);
    CN12_data_in(8) <= VN466_data_out(0);
    CN12_sign_in(8) <= VN466_sign_out(0);
    CN12_data_in(9) <= VN507_data_out(0);
    CN12_sign_in(9) <= VN507_sign_out(0);
    CN12_data_in(10) <= VN590_data_out(0);
    CN12_sign_in(10) <= VN590_sign_out(0);
    CN12_data_in(11) <= VN660_data_out(0);
    CN12_sign_in(11) <= VN660_sign_out(0);
    CN12_data_in(12) <= VN679_data_out(0);
    CN12_sign_in(12) <= VN679_sign_out(0);
    CN12_data_in(13) <= VN751_data_out(0);
    CN12_sign_in(13) <= VN751_sign_out(0);
    CN12_data_in(14) <= VN788_data_out(0);
    CN12_sign_in(14) <= VN788_sign_out(0);
    CN12_data_in(15) <= VN843_data_out(0);
    CN12_sign_in(15) <= VN843_sign_out(0);
    CN12_data_in(16) <= VN918_data_out(0);
    CN12_sign_in(16) <= VN918_sign_out(0);
    CN12_data_in(17) <= VN980_data_out(0);
    CN12_sign_in(17) <= VN980_sign_out(0);
    CN12_data_in(18) <= VN1067_data_out(0);
    CN12_sign_in(18) <= VN1067_sign_out(0);
    CN12_data_in(19) <= VN1128_data_out(0);
    CN12_sign_in(19) <= VN1128_sign_out(0);
    CN12_data_in(20) <= VN1192_data_out(0);
    CN12_sign_in(20) <= VN1192_sign_out(0);
    CN12_data_in(21) <= VN1268_data_out(0);
    CN12_sign_in(21) <= VN1268_sign_out(0);
    CN12_data_in(22) <= VN1284_data_out(0);
    CN12_sign_in(22) <= VN1284_sign_out(0);
    CN12_data_in(23) <= VN1377_data_out(0);
    CN12_sign_in(23) <= VN1377_sign_out(0);
    CN12_data_in(24) <= VN1433_data_out(0);
    CN12_sign_in(24) <= VN1433_sign_out(0);
    CN12_data_in(25) <= VN1453_data_out(0);
    CN12_sign_in(25) <= VN1453_sign_out(0);
    CN12_data_in(26) <= VN1487_data_out(0);
    CN12_sign_in(26) <= VN1487_sign_out(0);
    CN12_data_in(27) <= VN1540_data_out(0);
    CN12_sign_in(27) <= VN1540_sign_out(0);
    CN12_data_in(28) <= VN1639_data_out(0);
    CN12_sign_in(28) <= VN1639_sign_out(0);
    CN12_data_in(29) <= VN1672_data_out(0);
    CN12_sign_in(29) <= VN1672_sign_out(0);
    CN12_data_in(30) <= VN1703_data_out(0);
    CN12_sign_in(30) <= VN1703_sign_out(0);
    CN12_data_in(31) <= VN1729_data_out(0);
    CN12_sign_in(31) <= VN1729_sign_out(0);
    CN13_data_in(0) <= VN82_data_out(0);
    CN13_sign_in(0) <= VN82_sign_out(0);
    CN13_data_in(1) <= VN128_data_out(0);
    CN13_sign_in(1) <= VN128_sign_out(0);
    CN13_data_in(2) <= VN212_data_out(0);
    CN13_sign_in(2) <= VN212_sign_out(0);
    CN13_data_in(3) <= VN230_data_out(0);
    CN13_sign_in(3) <= VN230_sign_out(0);
    CN13_data_in(4) <= VN298_data_out(0);
    CN13_sign_in(4) <= VN298_sign_out(0);
    CN13_data_in(5) <= VN346_data_out(0);
    CN13_sign_in(5) <= VN346_sign_out(0);
    CN13_data_in(6) <= VN398_data_out(0);
    CN13_sign_in(6) <= VN398_sign_out(0);
    CN13_data_in(7) <= VN465_data_out(0);
    CN13_sign_in(7) <= VN465_sign_out(0);
    CN13_data_in(8) <= VN506_data_out(0);
    CN13_sign_in(8) <= VN506_sign_out(0);
    CN13_data_in(9) <= VN589_data_out(0);
    CN13_sign_in(9) <= VN589_sign_out(0);
    CN13_data_in(10) <= VN659_data_out(0);
    CN13_sign_in(10) <= VN659_sign_out(0);
    CN13_data_in(11) <= VN678_data_out(0);
    CN13_sign_in(11) <= VN678_sign_out(0);
    CN13_data_in(12) <= VN750_data_out(0);
    CN13_sign_in(12) <= VN750_sign_out(0);
    CN13_data_in(13) <= VN787_data_out(0);
    CN13_sign_in(13) <= VN787_sign_out(0);
    CN13_data_in(14) <= VN842_data_out(0);
    CN13_sign_in(14) <= VN842_sign_out(0);
    CN13_data_in(15) <= VN917_data_out(0);
    CN13_sign_in(15) <= VN917_sign_out(0);
    CN13_data_in(16) <= VN979_data_out(0);
    CN13_sign_in(16) <= VN979_sign_out(0);
    CN13_data_in(17) <= VN1013_data_out(0);
    CN13_sign_in(17) <= VN1013_sign_out(0);
    CN13_data_in(18) <= VN1066_data_out(0);
    CN13_sign_in(18) <= VN1066_sign_out(0);
    CN13_data_in(19) <= VN1127_data_out(0);
    CN13_sign_in(19) <= VN1127_sign_out(0);
    CN13_data_in(20) <= VN1191_data_out(0);
    CN13_sign_in(20) <= VN1191_sign_out(0);
    CN13_data_in(21) <= VN1267_data_out(0);
    CN13_sign_in(21) <= VN1267_sign_out(0);
    CN13_data_in(22) <= VN1283_data_out(0);
    CN13_sign_in(22) <= VN1283_sign_out(0);
    CN13_data_in(23) <= VN1376_data_out(0);
    CN13_sign_in(23) <= VN1376_sign_out(0);
    CN13_data_in(24) <= VN1432_data_out(0);
    CN13_sign_in(24) <= VN1432_sign_out(0);
    CN13_data_in(25) <= VN1452_data_out(0);
    CN13_sign_in(25) <= VN1452_sign_out(0);
    CN13_data_in(26) <= VN1576_data_out(0);
    CN13_sign_in(26) <= VN1576_sign_out(0);
    CN13_data_in(27) <= VN1638_data_out(0);
    CN13_sign_in(27) <= VN1638_sign_out(0);
    CN13_data_in(28) <= VN1671_data_out(0);
    CN13_sign_in(28) <= VN1671_sign_out(0);
    CN13_data_in(29) <= VN1702_data_out(0);
    CN13_sign_in(29) <= VN1702_sign_out(0);
    CN13_data_in(30) <= VN1750_data_out(0);
    CN13_sign_in(30) <= VN1750_sign_out(0);
    CN13_data_in(31) <= VN1810_data_out(0);
    CN13_sign_in(31) <= VN1810_sign_out(0);
    CN14_data_in(0) <= VN40_data_out(0);
    CN14_sign_in(0) <= VN40_sign_out(0);
    CN14_data_in(1) <= VN81_data_out(0);
    CN14_sign_in(1) <= VN81_sign_out(0);
    CN14_data_in(2) <= VN127_data_out(0);
    CN14_sign_in(2) <= VN127_sign_out(0);
    CN14_data_in(3) <= VN211_data_out(0);
    CN14_sign_in(3) <= VN211_sign_out(0);
    CN14_data_in(4) <= VN229_data_out(0);
    CN14_sign_in(4) <= VN229_sign_out(0);
    CN14_data_in(5) <= VN297_data_out(0);
    CN14_sign_in(5) <= VN297_sign_out(0);
    CN14_data_in(6) <= VN345_data_out(0);
    CN14_sign_in(6) <= VN345_sign_out(0);
    CN14_data_in(7) <= VN397_data_out(0);
    CN14_sign_in(7) <= VN397_sign_out(0);
    CN14_data_in(8) <= VN464_data_out(0);
    CN14_sign_in(8) <= VN464_sign_out(0);
    CN14_data_in(9) <= VN560_data_out(0);
    CN14_sign_in(9) <= VN560_sign_out(0);
    CN14_data_in(10) <= VN588_data_out(0);
    CN14_sign_in(10) <= VN588_sign_out(0);
    CN14_data_in(11) <= VN658_data_out(0);
    CN14_sign_in(11) <= VN658_sign_out(0);
    CN14_data_in(12) <= VN677_data_out(0);
    CN14_sign_in(12) <= VN677_sign_out(0);
    CN14_data_in(13) <= VN749_data_out(0);
    CN14_sign_in(13) <= VN749_sign_out(0);
    CN14_data_in(14) <= VN786_data_out(0);
    CN14_sign_in(14) <= VN786_sign_out(0);
    CN14_data_in(15) <= VN841_data_out(0);
    CN14_sign_in(15) <= VN841_sign_out(0);
    CN14_data_in(16) <= VN916_data_out(0);
    CN14_sign_in(16) <= VN916_sign_out(0);
    CN14_data_in(17) <= VN978_data_out(0);
    CN14_sign_in(17) <= VN978_sign_out(0);
    CN14_data_in(18) <= VN1012_data_out(0);
    CN14_sign_in(18) <= VN1012_sign_out(0);
    CN14_data_in(19) <= VN1065_data_out(0);
    CN14_sign_in(19) <= VN1065_sign_out(0);
    CN14_data_in(20) <= VN1126_data_out(0);
    CN14_sign_in(20) <= VN1126_sign_out(0);
    CN14_data_in(21) <= VN1190_data_out(0);
    CN14_sign_in(21) <= VN1190_sign_out(0);
    CN14_data_in(22) <= VN1266_data_out(0);
    CN14_sign_in(22) <= VN1266_sign_out(0);
    CN14_data_in(23) <= VN1375_data_out(0);
    CN14_sign_in(23) <= VN1375_sign_out(0);
    CN14_data_in(24) <= VN1431_data_out(0);
    CN14_sign_in(24) <= VN1431_sign_out(0);
    CN14_data_in(25) <= VN1451_data_out(0);
    CN14_sign_in(25) <= VN1451_sign_out(0);
    CN14_data_in(26) <= VN1486_data_out(0);
    CN14_sign_in(26) <= VN1486_sign_out(0);
    CN14_data_in(27) <= VN1531_data_out(0);
    CN14_sign_in(27) <= VN1531_sign_out(0);
    CN14_data_in(28) <= VN1539_data_out(0);
    CN14_sign_in(28) <= VN1539_sign_out(0);
    CN14_data_in(29) <= VN1637_data_out(0);
    CN14_sign_in(29) <= VN1637_sign_out(0);
    CN14_data_in(30) <= VN1778_data_out(0);
    CN14_sign_in(30) <= VN1778_sign_out(0);
    CN14_data_in(31) <= VN1811_data_out(0);
    CN14_sign_in(31) <= VN1811_sign_out(0);
    CN15_data_in(0) <= VN39_data_out(0);
    CN15_sign_in(0) <= VN39_sign_out(0);
    CN15_data_in(1) <= VN80_data_out(0);
    CN15_sign_in(1) <= VN80_sign_out(0);
    CN15_data_in(2) <= VN126_data_out(0);
    CN15_sign_in(2) <= VN126_sign_out(0);
    CN15_data_in(3) <= VN210_data_out(0);
    CN15_sign_in(3) <= VN210_sign_out(0);
    CN15_data_in(4) <= VN228_data_out(0);
    CN15_sign_in(4) <= VN228_sign_out(0);
    CN15_data_in(5) <= VN296_data_out(0);
    CN15_sign_in(5) <= VN296_sign_out(0);
    CN15_data_in(6) <= VN344_data_out(0);
    CN15_sign_in(6) <= VN344_sign_out(0);
    CN15_data_in(7) <= VN396_data_out(0);
    CN15_sign_in(7) <= VN396_sign_out(0);
    CN15_data_in(8) <= VN559_data_out(0);
    CN15_sign_in(8) <= VN559_sign_out(0);
    CN15_data_in(9) <= VN657_data_out(0);
    CN15_sign_in(9) <= VN657_sign_out(0);
    CN15_data_in(10) <= VN785_data_out(0);
    CN15_sign_in(10) <= VN785_sign_out(0);
    CN15_data_in(11) <= VN840_data_out(0);
    CN15_sign_in(11) <= VN840_sign_out(0);
    CN15_data_in(12) <= VN915_data_out(0);
    CN15_sign_in(12) <= VN915_sign_out(0);
    CN15_data_in(13) <= VN977_data_out(0);
    CN15_sign_in(13) <= VN977_sign_out(0);
    CN15_data_in(14) <= VN1011_data_out(0);
    CN15_sign_in(14) <= VN1011_sign_out(0);
    CN15_data_in(15) <= VN1064_data_out(0);
    CN15_sign_in(15) <= VN1064_sign_out(0);
    CN15_data_in(16) <= VN1125_data_out(0);
    CN15_sign_in(16) <= VN1125_sign_out(0);
    CN15_data_in(17) <= VN1189_data_out(0);
    CN15_sign_in(17) <= VN1189_sign_out(0);
    CN15_data_in(18) <= VN1265_data_out(0);
    CN15_sign_in(18) <= VN1265_sign_out(0);
    CN15_data_in(19) <= VN1374_data_out(0);
    CN15_sign_in(19) <= VN1374_sign_out(0);
    CN15_data_in(20) <= VN1450_data_out(0);
    CN15_sign_in(20) <= VN1450_sign_out(0);
    CN15_data_in(21) <= VN1483_data_out(0);
    CN15_sign_in(21) <= VN1483_sign_out(0);
    CN15_data_in(22) <= VN1530_data_out(0);
    CN15_sign_in(22) <= VN1530_sign_out(0);
    CN15_data_in(23) <= VN1701_data_out(0);
    CN15_sign_in(23) <= VN1701_sign_out(0);
    CN15_data_in(24) <= VN1753_data_out(0);
    CN15_sign_in(24) <= VN1753_sign_out(0);
    CN15_data_in(25) <= VN1809_data_out(0);
    CN15_sign_in(25) <= VN1809_sign_out(0);
    CN15_data_in(26) <= VN1842_data_out(0);
    CN15_sign_in(26) <= VN1842_sign_out(0);
    CN15_data_in(27) <= VN1910_data_out(0);
    CN15_sign_in(27) <= VN1910_sign_out(0);
    CN15_data_in(28) <= VN1925_data_out(0);
    CN15_sign_in(28) <= VN1925_sign_out(0);
    CN15_data_in(29) <= VN1937_data_out(0);
    CN15_sign_in(29) <= VN1937_sign_out(0);
    CN15_data_in(30) <= VN1953_data_out(0);
    CN15_sign_in(30) <= VN1953_sign_out(0);
    CN15_data_in(31) <= VN1961_data_out(0);
    CN15_sign_in(31) <= VN1961_sign_out(0);
    CN16_data_in(0) <= VN38_data_out(0);
    CN16_sign_in(0) <= VN38_sign_out(0);
    CN16_data_in(1) <= VN125_data_out(0);
    CN16_sign_in(1) <= VN125_sign_out(0);
    CN16_data_in(2) <= VN209_data_out(0);
    CN16_sign_in(2) <= VN209_sign_out(0);
    CN16_data_in(3) <= VN227_data_out(0);
    CN16_sign_in(3) <= VN227_sign_out(0);
    CN16_data_in(4) <= VN295_data_out(0);
    CN16_sign_in(4) <= VN295_sign_out(0);
    CN16_data_in(5) <= VN343_data_out(0);
    CN16_sign_in(5) <= VN343_sign_out(0);
    CN16_data_in(6) <= VN395_data_out(0);
    CN16_sign_in(6) <= VN395_sign_out(0);
    CN16_data_in(7) <= VN463_data_out(0);
    CN16_sign_in(7) <= VN463_sign_out(0);
    CN16_data_in(8) <= VN587_data_out(0);
    CN16_sign_in(8) <= VN587_sign_out(0);
    CN16_data_in(9) <= VN656_data_out(0);
    CN16_sign_in(9) <= VN656_sign_out(0);
    CN16_data_in(10) <= VN676_data_out(0);
    CN16_sign_in(10) <= VN676_sign_out(0);
    CN16_data_in(11) <= VN748_data_out(0);
    CN16_sign_in(11) <= VN748_sign_out(0);
    CN16_data_in(12) <= VN839_data_out(0);
    CN16_sign_in(12) <= VN839_sign_out(0);
    CN16_data_in(13) <= VN976_data_out(0);
    CN16_sign_in(13) <= VN976_sign_out(0);
    CN16_data_in(14) <= VN1010_data_out(0);
    CN16_sign_in(14) <= VN1010_sign_out(0);
    CN16_data_in(15) <= VN1063_data_out(0);
    CN16_sign_in(15) <= VN1063_sign_out(0);
    CN16_data_in(16) <= VN1124_data_out(0);
    CN16_sign_in(16) <= VN1124_sign_out(0);
    CN16_data_in(17) <= VN1188_data_out(0);
    CN16_sign_in(17) <= VN1188_sign_out(0);
    CN16_data_in(18) <= VN1264_data_out(0);
    CN16_sign_in(18) <= VN1264_sign_out(0);
    CN16_data_in(19) <= VN1373_data_out(0);
    CN16_sign_in(19) <= VN1373_sign_out(0);
    CN16_data_in(20) <= VN1430_data_out(0);
    CN16_sign_in(20) <= VN1430_sign_out(0);
    CN16_data_in(21) <= VN1482_data_out(0);
    CN16_sign_in(21) <= VN1482_sign_out(0);
    CN16_data_in(22) <= VN1529_data_out(0);
    CN16_sign_in(22) <= VN1529_sign_out(0);
    CN16_data_in(23) <= VN1538_data_out(0);
    CN16_sign_in(23) <= VN1538_sign_out(0);
    CN16_data_in(24) <= VN1636_data_out(0);
    CN16_sign_in(24) <= VN1636_sign_out(0);
    CN16_data_in(25) <= VN1670_data_out(0);
    CN16_sign_in(25) <= VN1670_sign_out(0);
    CN16_data_in(26) <= VN1700_data_out(0);
    CN16_sign_in(26) <= VN1700_sign_out(0);
    CN16_data_in(27) <= VN1900_data_out(0);
    CN16_sign_in(27) <= VN1900_sign_out(0);
    CN16_data_in(28) <= VN2006_data_out(0);
    CN16_sign_in(28) <= VN2006_sign_out(0);
    CN16_data_in(29) <= VN2023_data_out(0);
    CN16_sign_in(29) <= VN2023_sign_out(0);
    CN16_data_in(30) <= VN2034_data_out(0);
    CN16_sign_in(30) <= VN2034_sign_out(0);
    CN16_data_in(31) <= VN2036_data_out(0);
    CN16_sign_in(31) <= VN2036_sign_out(0);
    CN17_data_in(0) <= VN37_data_out(0);
    CN17_sign_in(0) <= VN37_sign_out(0);
    CN17_data_in(1) <= VN79_data_out(0);
    CN17_sign_in(1) <= VN79_sign_out(0);
    CN17_data_in(2) <= VN124_data_out(0);
    CN17_sign_in(2) <= VN124_sign_out(0);
    CN17_data_in(3) <= VN208_data_out(0);
    CN17_sign_in(3) <= VN208_sign_out(0);
    CN17_data_in(4) <= VN226_data_out(0);
    CN17_sign_in(4) <= VN226_sign_out(0);
    CN17_data_in(5) <= VN294_data_out(0);
    CN17_sign_in(5) <= VN294_sign_out(0);
    CN17_data_in(6) <= VN342_data_out(0);
    CN17_sign_in(6) <= VN342_sign_out(0);
    CN17_data_in(7) <= VN394_data_out(0);
    CN17_sign_in(7) <= VN394_sign_out(0);
    CN17_data_in(8) <= VN462_data_out(0);
    CN17_sign_in(8) <= VN462_sign_out(0);
    CN17_data_in(9) <= VN558_data_out(0);
    CN17_sign_in(9) <= VN558_sign_out(0);
    CN17_data_in(10) <= VN586_data_out(0);
    CN17_sign_in(10) <= VN586_sign_out(0);
    CN17_data_in(11) <= VN655_data_out(0);
    CN17_sign_in(11) <= VN655_sign_out(0);
    CN17_data_in(12) <= VN675_data_out(0);
    CN17_sign_in(12) <= VN675_sign_out(0);
    CN17_data_in(13) <= VN747_data_out(0);
    CN17_sign_in(13) <= VN747_sign_out(0);
    CN17_data_in(14) <= VN784_data_out(0);
    CN17_sign_in(14) <= VN784_sign_out(0);
    CN17_data_in(15) <= VN838_data_out(0);
    CN17_sign_in(15) <= VN838_sign_out(0);
    CN17_data_in(16) <= VN914_data_out(0);
    CN17_sign_in(16) <= VN914_sign_out(0);
    CN17_data_in(17) <= VN975_data_out(0);
    CN17_sign_in(17) <= VN975_sign_out(0);
    CN17_data_in(18) <= VN1009_data_out(0);
    CN17_sign_in(18) <= VN1009_sign_out(0);
    CN17_data_in(19) <= VN1062_data_out(0);
    CN17_sign_in(19) <= VN1062_sign_out(0);
    CN17_data_in(20) <= VN1123_data_out(0);
    CN17_sign_in(20) <= VN1123_sign_out(0);
    CN17_data_in(21) <= VN1187_data_out(0);
    CN17_sign_in(21) <= VN1187_sign_out(0);
    CN17_data_in(22) <= VN1263_data_out(0);
    CN17_sign_in(22) <= VN1263_sign_out(0);
    CN17_data_in(23) <= VN1372_data_out(0);
    CN17_sign_in(23) <= VN1372_sign_out(0);
    CN17_data_in(24) <= VN1429_data_out(0);
    CN17_sign_in(24) <= VN1429_sign_out(0);
    CN17_data_in(25) <= VN1449_data_out(0);
    CN17_sign_in(25) <= VN1449_sign_out(0);
    CN17_data_in(26) <= VN1481_data_out(0);
    CN17_sign_in(26) <= VN1481_sign_out(0);
    CN17_data_in(27) <= VN1528_data_out(0);
    CN17_sign_in(27) <= VN1528_sign_out(0);
    CN17_data_in(28) <= VN1699_data_out(0);
    CN17_sign_in(28) <= VN1699_sign_out(0);
    CN17_data_in(29) <= VN1786_data_out(0);
    CN17_sign_in(29) <= VN1786_sign_out(0);
    CN17_data_in(30) <= VN1807_data_out(0);
    CN17_sign_in(30) <= VN1807_sign_out(0);
    CN17_data_in(31) <= VN1812_data_out(0);
    CN17_sign_in(31) <= VN1812_sign_out(0);
    CN18_data_in(0) <= VN36_data_out(0);
    CN18_sign_in(0) <= VN36_sign_out(0);
    CN18_data_in(1) <= VN78_data_out(0);
    CN18_sign_in(1) <= VN78_sign_out(0);
    CN18_data_in(2) <= VN123_data_out(0);
    CN18_sign_in(2) <= VN123_sign_out(0);
    CN18_data_in(3) <= VN207_data_out(0);
    CN18_sign_in(3) <= VN207_sign_out(0);
    CN18_data_in(4) <= VN225_data_out(0);
    CN18_sign_in(4) <= VN225_sign_out(0);
    CN18_data_in(5) <= VN293_data_out(0);
    CN18_sign_in(5) <= VN293_sign_out(0);
    CN18_data_in(6) <= VN341_data_out(0);
    CN18_sign_in(6) <= VN341_sign_out(0);
    CN18_data_in(7) <= VN393_data_out(0);
    CN18_sign_in(7) <= VN393_sign_out(0);
    CN18_data_in(8) <= VN461_data_out(0);
    CN18_sign_in(8) <= VN461_sign_out(0);
    CN18_data_in(9) <= VN557_data_out(0);
    CN18_sign_in(9) <= VN557_sign_out(0);
    CN18_data_in(10) <= VN585_data_out(0);
    CN18_sign_in(10) <= VN585_sign_out(0);
    CN18_data_in(11) <= VN654_data_out(0);
    CN18_sign_in(11) <= VN654_sign_out(0);
    CN18_data_in(12) <= VN674_data_out(0);
    CN18_sign_in(12) <= VN674_sign_out(0);
    CN18_data_in(13) <= VN746_data_out(0);
    CN18_sign_in(13) <= VN746_sign_out(0);
    CN18_data_in(14) <= VN783_data_out(0);
    CN18_sign_in(14) <= VN783_sign_out(0);
    CN18_data_in(15) <= VN837_data_out(0);
    CN18_sign_in(15) <= VN837_sign_out(0);
    CN18_data_in(16) <= VN913_data_out(0);
    CN18_sign_in(16) <= VN913_sign_out(0);
    CN18_data_in(17) <= VN974_data_out(0);
    CN18_sign_in(17) <= VN974_sign_out(0);
    CN18_data_in(18) <= VN1008_data_out(0);
    CN18_sign_in(18) <= VN1008_sign_out(0);
    CN18_data_in(19) <= VN1061_data_out(0);
    CN18_sign_in(19) <= VN1061_sign_out(0);
    CN18_data_in(20) <= VN1122_data_out(0);
    CN18_sign_in(20) <= VN1122_sign_out(0);
    CN18_data_in(21) <= VN1186_data_out(0);
    CN18_sign_in(21) <= VN1186_sign_out(0);
    CN18_data_in(22) <= VN1262_data_out(0);
    CN18_sign_in(22) <= VN1262_sign_out(0);
    CN18_data_in(23) <= VN1371_data_out(0);
    CN18_sign_in(23) <= VN1371_sign_out(0);
    CN18_data_in(24) <= VN1428_data_out(0);
    CN18_sign_in(24) <= VN1428_sign_out(0);
    CN18_data_in(25) <= VN1448_data_out(0);
    CN18_sign_in(25) <= VN1448_sign_out(0);
    CN18_data_in(26) <= VN1480_data_out(0);
    CN18_sign_in(26) <= VN1480_sign_out(0);
    CN18_data_in(27) <= VN1527_data_out(0);
    CN18_sign_in(27) <= VN1527_sign_out(0);
    CN18_data_in(28) <= VN1537_data_out(0);
    CN18_sign_in(28) <= VN1537_sign_out(0);
    CN18_data_in(29) <= VN1635_data_out(0);
    CN18_sign_in(29) <= VN1635_sign_out(0);
    CN18_data_in(30) <= VN1698_data_out(0);
    CN18_sign_in(30) <= VN1698_sign_out(0);
    CN18_data_in(31) <= VN1730_data_out(0);
    CN18_sign_in(31) <= VN1730_sign_out(0);
    CN19_data_in(0) <= VN35_data_out(0);
    CN19_sign_in(0) <= VN35_sign_out(0);
    CN19_data_in(1) <= VN77_data_out(0);
    CN19_sign_in(1) <= VN77_sign_out(0);
    CN19_data_in(2) <= VN122_data_out(0);
    CN19_sign_in(2) <= VN122_sign_out(0);
    CN19_data_in(3) <= VN278_data_out(0);
    CN19_sign_in(3) <= VN278_sign_out(0);
    CN19_data_in(4) <= VN340_data_out(0);
    CN19_sign_in(4) <= VN340_sign_out(0);
    CN19_data_in(5) <= VN460_data_out(0);
    CN19_sign_in(5) <= VN460_sign_out(0);
    CN19_data_in(6) <= VN556_data_out(0);
    CN19_sign_in(6) <= VN556_sign_out(0);
    CN19_data_in(7) <= VN584_data_out(0);
    CN19_sign_in(7) <= VN584_sign_out(0);
    CN19_data_in(8) <= VN745_data_out(0);
    CN19_sign_in(8) <= VN745_sign_out(0);
    CN19_data_in(9) <= VN782_data_out(0);
    CN19_sign_in(9) <= VN782_sign_out(0);
    CN19_data_in(10) <= VN836_data_out(0);
    CN19_sign_in(10) <= VN836_sign_out(0);
    CN19_data_in(11) <= VN912_data_out(0);
    CN19_sign_in(11) <= VN912_sign_out(0);
    CN19_data_in(12) <= VN973_data_out(0);
    CN19_sign_in(12) <= VN973_sign_out(0);
    CN19_data_in(13) <= VN1261_data_out(0);
    CN19_sign_in(13) <= VN1261_sign_out(0);
    CN19_data_in(14) <= VN1370_data_out(0);
    CN19_sign_in(14) <= VN1370_sign_out(0);
    CN19_data_in(15) <= VN1447_data_out(0);
    CN19_sign_in(15) <= VN1447_sign_out(0);
    CN19_data_in(16) <= VN1479_data_out(0);
    CN19_sign_in(16) <= VN1479_sign_out(0);
    CN19_data_in(17) <= VN1526_data_out(0);
    CN19_sign_in(17) <= VN1526_sign_out(0);
    CN19_data_in(18) <= VN1634_data_out(0);
    CN19_sign_in(18) <= VN1634_sign_out(0);
    CN19_data_in(19) <= VN1669_data_out(0);
    CN19_sign_in(19) <= VN1669_sign_out(0);
    CN19_data_in(20) <= VN1697_data_out(0);
    CN19_sign_in(20) <= VN1697_sign_out(0);
    CN19_data_in(21) <= VN1772_data_out(0);
    CN19_sign_in(21) <= VN1772_sign_out(0);
    CN19_data_in(22) <= VN1849_data_out(0);
    CN19_sign_in(22) <= VN1849_sign_out(0);
    CN19_data_in(23) <= VN1884_data_out(0);
    CN19_sign_in(23) <= VN1884_sign_out(0);
    CN19_data_in(24) <= VN1885_data_out(0);
    CN19_sign_in(24) <= VN1885_sign_out(0);
    CN19_data_in(25) <= VN1957_data_out(0);
    CN19_sign_in(25) <= VN1957_sign_out(0);
    CN19_data_in(26) <= VN1964_data_out(0);
    CN19_sign_in(26) <= VN1964_sign_out(0);
    CN19_data_in(27) <= VN1986_data_out(0);
    CN19_sign_in(27) <= VN1986_sign_out(0);
    CN19_data_in(28) <= VN1989_data_out(0);
    CN19_sign_in(28) <= VN1989_sign_out(0);
    CN19_data_in(29) <= VN2028_data_out(0);
    CN19_sign_in(29) <= VN2028_sign_out(0);
    CN19_data_in(30) <= VN2041_data_out(0);
    CN19_sign_in(30) <= VN2041_sign_out(0);
    CN19_data_in(31) <= VN2042_data_out(0);
    CN19_sign_in(31) <= VN2042_sign_out(0);
    CN20_data_in(0) <= VN34_data_out(0);
    CN20_sign_in(0) <= VN34_sign_out(0);
    CN20_data_in(1) <= VN76_data_out(0);
    CN20_sign_in(1) <= VN76_sign_out(0);
    CN20_data_in(2) <= VN277_data_out(0);
    CN20_sign_in(2) <= VN277_sign_out(0);
    CN20_data_in(3) <= VN292_data_out(0);
    CN20_sign_in(3) <= VN292_sign_out(0);
    CN20_data_in(4) <= VN339_data_out(0);
    CN20_sign_in(4) <= VN339_sign_out(0);
    CN20_data_in(5) <= VN459_data_out(0);
    CN20_sign_in(5) <= VN459_sign_out(0);
    CN20_data_in(6) <= VN555_data_out(0);
    CN20_sign_in(6) <= VN555_sign_out(0);
    CN20_data_in(7) <= VN583_data_out(0);
    CN20_sign_in(7) <= VN583_sign_out(0);
    CN20_data_in(8) <= VN673_data_out(0);
    CN20_sign_in(8) <= VN673_sign_out(0);
    CN20_data_in(9) <= VN781_data_out(0);
    CN20_sign_in(9) <= VN781_sign_out(0);
    CN20_data_in(10) <= VN911_data_out(0);
    CN20_sign_in(10) <= VN911_sign_out(0);
    CN20_data_in(11) <= VN972_data_out(0);
    CN20_sign_in(11) <= VN972_sign_out(0);
    CN20_data_in(12) <= VN1007_data_out(0);
    CN20_sign_in(12) <= VN1007_sign_out(0);
    CN20_data_in(13) <= VN1121_data_out(0);
    CN20_sign_in(13) <= VN1121_sign_out(0);
    CN20_data_in(14) <= VN1185_data_out(0);
    CN20_sign_in(14) <= VN1185_sign_out(0);
    CN20_data_in(15) <= VN1260_data_out(0);
    CN20_sign_in(15) <= VN1260_sign_out(0);
    CN20_data_in(16) <= VN1328_data_out(0);
    CN20_sign_in(16) <= VN1328_sign_out(0);
    CN20_data_in(17) <= VN1427_data_out(0);
    CN20_sign_in(17) <= VN1427_sign_out(0);
    CN20_data_in(18) <= VN1446_data_out(0);
    CN20_sign_in(18) <= VN1446_sign_out(0);
    CN20_data_in(19) <= VN1478_data_out(0);
    CN20_sign_in(19) <= VN1478_sign_out(0);
    CN20_data_in(20) <= VN1508_data_out(0);
    CN20_sign_in(20) <= VN1508_sign_out(0);
    CN20_data_in(21) <= VN1633_data_out(0);
    CN20_sign_in(21) <= VN1633_sign_out(0);
    CN20_data_in(22) <= VN1696_data_out(0);
    CN20_sign_in(22) <= VN1696_sign_out(0);
    CN20_data_in(23) <= VN1770_data_out(0);
    CN20_sign_in(23) <= VN1770_sign_out(0);
    CN20_data_in(24) <= VN1773_data_out(0);
    CN20_sign_in(24) <= VN1773_sign_out(0);
    CN20_data_in(25) <= VN1787_data_out(0);
    CN20_sign_in(25) <= VN1787_sign_out(0);
    CN20_data_in(26) <= VN1844_data_out(0);
    CN20_sign_in(26) <= VN1844_sign_out(0);
    CN20_data_in(27) <= VN1852_data_out(0);
    CN20_sign_in(27) <= VN1852_sign_out(0);
    CN20_data_in(28) <= VN1854_data_out(0);
    CN20_sign_in(28) <= VN1854_sign_out(0);
    CN20_data_in(29) <= VN1857_data_out(0);
    CN20_sign_in(29) <= VN1857_sign_out(0);
    CN20_data_in(30) <= VN1858_data_out(0);
    CN20_sign_in(30) <= VN1858_sign_out(0);
    CN20_data_in(31) <= VN1876_data_out(0);
    CN20_sign_in(31) <= VN1876_sign_out(0);
    CN21_data_in(0) <= VN33_data_out(0);
    CN21_sign_in(0) <= VN33_sign_out(0);
    CN21_data_in(1) <= VN75_data_out(0);
    CN21_sign_in(1) <= VN75_sign_out(0);
    CN21_data_in(2) <= VN121_data_out(0);
    CN21_sign_in(2) <= VN121_sign_out(0);
    CN21_data_in(3) <= VN206_data_out(0);
    CN21_sign_in(3) <= VN206_sign_out(0);
    CN21_data_in(4) <= VN276_data_out(0);
    CN21_sign_in(4) <= VN276_sign_out(0);
    CN21_data_in(5) <= VN291_data_out(0);
    CN21_sign_in(5) <= VN291_sign_out(0);
    CN21_data_in(6) <= VN338_data_out(0);
    CN21_sign_in(6) <= VN338_sign_out(0);
    CN21_data_in(7) <= VN392_data_out(0);
    CN21_sign_in(7) <= VN392_sign_out(0);
    CN21_data_in(8) <= VN458_data_out(0);
    CN21_sign_in(8) <= VN458_sign_out(0);
    CN21_data_in(9) <= VN554_data_out(0);
    CN21_sign_in(9) <= VN554_sign_out(0);
    CN21_data_in(10) <= VN653_data_out(0);
    CN21_sign_in(10) <= VN653_sign_out(0);
    CN21_data_in(11) <= VN672_data_out(0);
    CN21_sign_in(11) <= VN672_sign_out(0);
    CN21_data_in(12) <= VN744_data_out(0);
    CN21_sign_in(12) <= VN744_sign_out(0);
    CN21_data_in(13) <= VN780_data_out(0);
    CN21_sign_in(13) <= VN780_sign_out(0);
    CN21_data_in(14) <= VN835_data_out(0);
    CN21_sign_in(14) <= VN835_sign_out(0);
    CN21_data_in(15) <= VN910_data_out(0);
    CN21_sign_in(15) <= VN910_sign_out(0);
    CN21_data_in(16) <= VN971_data_out(0);
    CN21_sign_in(16) <= VN971_sign_out(0);
    CN21_data_in(17) <= VN1006_data_out(0);
    CN21_sign_in(17) <= VN1006_sign_out(0);
    CN21_data_in(18) <= VN1111_data_out(0);
    CN21_sign_in(18) <= VN1111_sign_out(0);
    CN21_data_in(19) <= VN1120_data_out(0);
    CN21_sign_in(19) <= VN1120_sign_out(0);
    CN21_data_in(20) <= VN1184_data_out(0);
    CN21_sign_in(20) <= VN1184_sign_out(0);
    CN21_data_in(21) <= VN1259_data_out(0);
    CN21_sign_in(21) <= VN1259_sign_out(0);
    CN21_data_in(22) <= VN1327_data_out(0);
    CN21_sign_in(22) <= VN1327_sign_out(0);
    CN21_data_in(23) <= VN1369_data_out(0);
    CN21_sign_in(23) <= VN1369_sign_out(0);
    CN21_data_in(24) <= VN1425_data_out(0);
    CN21_sign_in(24) <= VN1425_sign_out(0);
    CN21_data_in(25) <= VN1426_data_out(0);
    CN21_sign_in(25) <= VN1426_sign_out(0);
    CN21_data_in(26) <= VN1445_data_out(0);
    CN21_sign_in(26) <= VN1445_sign_out(0);
    CN21_data_in(27) <= VN1477_data_out(0);
    CN21_sign_in(27) <= VN1477_sign_out(0);
    CN21_data_in(28) <= VN1632_data_out(0);
    CN21_sign_in(28) <= VN1632_sign_out(0);
    CN21_data_in(29) <= VN1668_data_out(0);
    CN21_sign_in(29) <= VN1668_sign_out(0);
    CN21_data_in(30) <= VN1932_data_out(0);
    CN21_sign_in(30) <= VN1932_sign_out(0);
    CN21_data_in(31) <= VN1934_data_out(0);
    CN21_sign_in(31) <= VN1934_sign_out(0);
    CN22_data_in(0) <= VN32_data_out(0);
    CN22_sign_in(0) <= VN32_sign_out(0);
    CN22_data_in(1) <= VN74_data_out(0);
    CN22_sign_in(1) <= VN74_sign_out(0);
    CN22_data_in(2) <= VN120_data_out(0);
    CN22_sign_in(2) <= VN120_sign_out(0);
    CN22_data_in(3) <= VN205_data_out(0);
    CN22_sign_in(3) <= VN205_sign_out(0);
    CN22_data_in(4) <= VN275_data_out(0);
    CN22_sign_in(4) <= VN275_sign_out(0);
    CN22_data_in(5) <= VN290_data_out(0);
    CN22_sign_in(5) <= VN290_sign_out(0);
    CN22_data_in(6) <= VN337_data_out(0);
    CN22_sign_in(6) <= VN337_sign_out(0);
    CN22_data_in(7) <= VN446_data_out(0);
    CN22_sign_in(7) <= VN446_sign_out(0);
    CN22_data_in(8) <= VN457_data_out(0);
    CN22_sign_in(8) <= VN457_sign_out(0);
    CN22_data_in(9) <= VN582_data_out(0);
    CN22_sign_in(9) <= VN582_sign_out(0);
    CN22_data_in(10) <= VN671_data_out(0);
    CN22_sign_in(10) <= VN671_sign_out(0);
    CN22_data_in(11) <= VN743_data_out(0);
    CN22_sign_in(11) <= VN743_sign_out(0);
    CN22_data_in(12) <= VN834_data_out(0);
    CN22_sign_in(12) <= VN834_sign_out(0);
    CN22_data_in(13) <= VN970_data_out(0);
    CN22_sign_in(13) <= VN970_sign_out(0);
    CN22_data_in(14) <= VN1119_data_out(0);
    CN22_sign_in(14) <= VN1119_sign_out(0);
    CN22_data_in(15) <= VN1183_data_out(0);
    CN22_sign_in(15) <= VN1183_sign_out(0);
    CN22_data_in(16) <= VN1258_data_out(0);
    CN22_sign_in(16) <= VN1258_sign_out(0);
    CN22_data_in(17) <= VN1326_data_out(0);
    CN22_sign_in(17) <= VN1326_sign_out(0);
    CN22_data_in(18) <= VN1368_data_out(0);
    CN22_sign_in(18) <= VN1368_sign_out(0);
    CN22_data_in(19) <= VN1390_data_out(0);
    CN22_sign_in(19) <= VN1390_sign_out(0);
    CN22_data_in(20) <= VN1424_data_out(0);
    CN22_sign_in(20) <= VN1424_sign_out(0);
    CN22_data_in(21) <= VN1507_data_out(0);
    CN22_sign_in(21) <= VN1507_sign_out(0);
    CN22_data_in(22) <= VN1631_data_out(0);
    CN22_sign_in(22) <= VN1631_sign_out(0);
    CN22_data_in(23) <= VN1765_data_out(0);
    CN22_sign_in(23) <= VN1765_sign_out(0);
    CN22_data_in(24) <= VN1793_data_out(0);
    CN22_sign_in(24) <= VN1793_sign_out(0);
    CN22_data_in(25) <= VN1795_data_out(0);
    CN22_sign_in(25) <= VN1795_sign_out(0);
    CN22_data_in(26) <= VN1882_data_out(0);
    CN22_sign_in(26) <= VN1882_sign_out(0);
    CN22_data_in(27) <= VN1903_data_out(0);
    CN22_sign_in(27) <= VN1903_sign_out(0);
    CN22_data_in(28) <= VN1941_data_out(0);
    CN22_sign_in(28) <= VN1941_sign_out(0);
    CN22_data_in(29) <= VN1987_data_out(0);
    CN22_sign_in(29) <= VN1987_sign_out(0);
    CN22_data_in(30) <= VN2032_data_out(0);
    CN22_sign_in(30) <= VN2032_sign_out(0);
    CN22_data_in(31) <= VN2035_data_out(0);
    CN22_sign_in(31) <= VN2035_sign_out(0);
    CN23_data_in(0) <= VN31_data_out(0);
    CN23_sign_in(0) <= VN31_sign_out(0);
    CN23_data_in(1) <= VN73_data_out(0);
    CN23_sign_in(1) <= VN73_sign_out(0);
    CN23_data_in(2) <= VN119_data_out(0);
    CN23_sign_in(2) <= VN119_sign_out(0);
    CN23_data_in(3) <= VN204_data_out(0);
    CN23_sign_in(3) <= VN204_sign_out(0);
    CN23_data_in(4) <= VN274_data_out(0);
    CN23_sign_in(4) <= VN274_sign_out(0);
    CN23_data_in(5) <= VN289_data_out(0);
    CN23_sign_in(5) <= VN289_sign_out(0);
    CN23_data_in(6) <= VN336_data_out(0);
    CN23_sign_in(6) <= VN336_sign_out(0);
    CN23_data_in(7) <= VN445_data_out(0);
    CN23_sign_in(7) <= VN445_sign_out(0);
    CN23_data_in(8) <= VN456_data_out(0);
    CN23_sign_in(8) <= VN456_sign_out(0);
    CN23_data_in(9) <= VN553_data_out(0);
    CN23_sign_in(9) <= VN553_sign_out(0);
    CN23_data_in(10) <= VN581_data_out(0);
    CN23_sign_in(10) <= VN581_sign_out(0);
    CN23_data_in(11) <= VN652_data_out(0);
    CN23_sign_in(11) <= VN652_sign_out(0);
    CN23_data_in(12) <= VN742_data_out(0);
    CN23_sign_in(12) <= VN742_sign_out(0);
    CN23_data_in(13) <= VN779_data_out(0);
    CN23_sign_in(13) <= VN779_sign_out(0);
    CN23_data_in(14) <= VN833_data_out(0);
    CN23_sign_in(14) <= VN833_sign_out(0);
    CN23_data_in(15) <= VN909_data_out(0);
    CN23_sign_in(15) <= VN909_sign_out(0);
    CN23_data_in(16) <= VN969_data_out(0);
    CN23_sign_in(16) <= VN969_sign_out(0);
    CN23_data_in(17) <= VN1005_data_out(0);
    CN23_sign_in(17) <= VN1005_sign_out(0);
    CN23_data_in(18) <= VN1109_data_out(0);
    CN23_sign_in(18) <= VN1109_sign_out(0);
    CN23_data_in(19) <= VN1118_data_out(0);
    CN23_sign_in(19) <= VN1118_sign_out(0);
    CN23_data_in(20) <= VN1182_data_out(0);
    CN23_sign_in(20) <= VN1182_sign_out(0);
    CN23_data_in(21) <= VN1257_data_out(0);
    CN23_sign_in(21) <= VN1257_sign_out(0);
    CN23_data_in(22) <= VN1325_data_out(0);
    CN23_sign_in(22) <= VN1325_sign_out(0);
    CN23_data_in(23) <= VN1367_data_out(0);
    CN23_sign_in(23) <= VN1367_sign_out(0);
    CN23_data_in(24) <= VN1389_data_out(0);
    CN23_sign_in(24) <= VN1389_sign_out(0);
    CN23_data_in(25) <= VN1423_data_out(0);
    CN23_sign_in(25) <= VN1423_sign_out(0);
    CN23_data_in(26) <= VN1444_data_out(0);
    CN23_sign_in(26) <= VN1444_sign_out(0);
    CN23_data_in(27) <= VN1476_data_out(0);
    CN23_sign_in(27) <= VN1476_sign_out(0);
    CN23_data_in(28) <= VN1630_data_out(0);
    CN23_sign_in(28) <= VN1630_sign_out(0);
    CN23_data_in(29) <= VN1754_data_out(0);
    CN23_sign_in(29) <= VN1754_sign_out(0);
    CN23_data_in(30) <= VN1802_data_out(0);
    CN23_sign_in(30) <= VN1802_sign_out(0);
    CN23_data_in(31) <= VN1813_data_out(0);
    CN23_sign_in(31) <= VN1813_sign_out(0);
    CN24_data_in(0) <= VN30_data_out(0);
    CN24_sign_in(0) <= VN30_sign_out(0);
    CN24_data_in(1) <= VN72_data_out(0);
    CN24_sign_in(1) <= VN72_sign_out(0);
    CN24_data_in(2) <= VN118_data_out(0);
    CN24_sign_in(2) <= VN118_sign_out(0);
    CN24_data_in(3) <= VN203_data_out(0);
    CN24_sign_in(3) <= VN203_sign_out(0);
    CN24_data_in(4) <= VN273_data_out(0);
    CN24_sign_in(4) <= VN273_sign_out(0);
    CN24_data_in(5) <= VN288_data_out(0);
    CN24_sign_in(5) <= VN288_sign_out(0);
    CN24_data_in(6) <= VN335_data_out(0);
    CN24_sign_in(6) <= VN335_sign_out(0);
    CN24_data_in(7) <= VN444_data_out(0);
    CN24_sign_in(7) <= VN444_sign_out(0);
    CN24_data_in(8) <= VN455_data_out(0);
    CN24_sign_in(8) <= VN455_sign_out(0);
    CN24_data_in(9) <= VN552_data_out(0);
    CN24_sign_in(9) <= VN552_sign_out(0);
    CN24_data_in(10) <= VN580_data_out(0);
    CN24_sign_in(10) <= VN580_sign_out(0);
    CN24_data_in(11) <= VN651_data_out(0);
    CN24_sign_in(11) <= VN651_sign_out(0);
    CN24_data_in(12) <= VN670_data_out(0);
    CN24_sign_in(12) <= VN670_sign_out(0);
    CN24_data_in(13) <= VN741_data_out(0);
    CN24_sign_in(13) <= VN741_sign_out(0);
    CN24_data_in(14) <= VN778_data_out(0);
    CN24_sign_in(14) <= VN778_sign_out(0);
    CN24_data_in(15) <= VN832_data_out(0);
    CN24_sign_in(15) <= VN832_sign_out(0);
    CN24_data_in(16) <= VN908_data_out(0);
    CN24_sign_in(16) <= VN908_sign_out(0);
    CN24_data_in(17) <= VN968_data_out(0);
    CN24_sign_in(17) <= VN968_sign_out(0);
    CN24_data_in(18) <= VN1004_data_out(0);
    CN24_sign_in(18) <= VN1004_sign_out(0);
    CN24_data_in(19) <= VN1117_data_out(0);
    CN24_sign_in(19) <= VN1117_sign_out(0);
    CN24_data_in(20) <= VN1181_data_out(0);
    CN24_sign_in(20) <= VN1181_sign_out(0);
    CN24_data_in(21) <= VN1324_data_out(0);
    CN24_sign_in(21) <= VN1324_sign_out(0);
    CN24_data_in(22) <= VN1366_data_out(0);
    CN24_sign_in(22) <= VN1366_sign_out(0);
    CN24_data_in(23) <= VN1388_data_out(0);
    CN24_sign_in(23) <= VN1388_sign_out(0);
    CN24_data_in(24) <= VN1422_data_out(0);
    CN24_sign_in(24) <= VN1422_sign_out(0);
    CN24_data_in(25) <= VN1443_data_out(0);
    CN24_sign_in(25) <= VN1443_sign_out(0);
    CN24_data_in(26) <= VN1506_data_out(0);
    CN24_sign_in(26) <= VN1506_sign_out(0);
    CN24_data_in(27) <= VN1667_data_out(0);
    CN24_sign_in(27) <= VN1667_sign_out(0);
    CN24_data_in(28) <= VN1695_data_out(0);
    CN24_sign_in(28) <= VN1695_sign_out(0);
    CN24_data_in(29) <= VN1760_data_out(0);
    CN24_sign_in(29) <= VN1760_sign_out(0);
    CN24_data_in(30) <= VN1784_data_out(0);
    CN24_sign_in(30) <= VN1784_sign_out(0);
    CN24_data_in(31) <= VN1814_data_out(0);
    CN24_sign_in(31) <= VN1814_sign_out(0);
    CN25_data_in(0) <= VN29_data_out(0);
    CN25_sign_in(0) <= VN29_sign_out(0);
    CN25_data_in(1) <= VN71_data_out(0);
    CN25_sign_in(1) <= VN71_sign_out(0);
    CN25_data_in(2) <= VN117_data_out(0);
    CN25_sign_in(2) <= VN117_sign_out(0);
    CN25_data_in(3) <= VN202_data_out(0);
    CN25_sign_in(3) <= VN202_sign_out(0);
    CN25_data_in(4) <= VN287_data_out(0);
    CN25_sign_in(4) <= VN287_sign_out(0);
    CN25_data_in(5) <= VN443_data_out(0);
    CN25_sign_in(5) <= VN443_sign_out(0);
    CN25_data_in(6) <= VN454_data_out(0);
    CN25_sign_in(6) <= VN454_sign_out(0);
    CN25_data_in(7) <= VN551_data_out(0);
    CN25_sign_in(7) <= VN551_sign_out(0);
    CN25_data_in(8) <= VN579_data_out(0);
    CN25_sign_in(8) <= VN579_sign_out(0);
    CN25_data_in(9) <= VN650_data_out(0);
    CN25_sign_in(9) <= VN650_sign_out(0);
    CN25_data_in(10) <= VN669_data_out(0);
    CN25_sign_in(10) <= VN669_sign_out(0);
    CN25_data_in(11) <= VN740_data_out(0);
    CN25_sign_in(11) <= VN740_sign_out(0);
    CN25_data_in(12) <= VN831_data_out(0);
    CN25_sign_in(12) <= VN831_sign_out(0);
    CN25_data_in(13) <= VN907_data_out(0);
    CN25_sign_in(13) <= VN907_sign_out(0);
    CN25_data_in(14) <= VN967_data_out(0);
    CN25_sign_in(14) <= VN967_sign_out(0);
    CN25_data_in(15) <= VN1107_data_out(0);
    CN25_sign_in(15) <= VN1107_sign_out(0);
    CN25_data_in(16) <= VN1116_data_out(0);
    CN25_sign_in(16) <= VN1116_sign_out(0);
    CN25_data_in(17) <= VN1180_data_out(0);
    CN25_sign_in(17) <= VN1180_sign_out(0);
    CN25_data_in(18) <= VN1256_data_out(0);
    CN25_sign_in(18) <= VN1256_sign_out(0);
    CN25_data_in(19) <= VN1323_data_out(0);
    CN25_sign_in(19) <= VN1323_sign_out(0);
    CN25_data_in(20) <= VN1365_data_out(0);
    CN25_sign_in(20) <= VN1365_sign_out(0);
    CN25_data_in(21) <= VN1387_data_out(0);
    CN25_sign_in(21) <= VN1387_sign_out(0);
    CN25_data_in(22) <= VN1466_data_out(0);
    CN25_sign_in(22) <= VN1466_sign_out(0);
    CN25_data_in(23) <= VN1504_data_out(0);
    CN25_sign_in(23) <= VN1504_sign_out(0);
    CN25_data_in(24) <= VN1629_data_out(0);
    CN25_sign_in(24) <= VN1629_sign_out(0);
    CN25_data_in(25) <= VN1759_data_out(0);
    CN25_sign_in(25) <= VN1759_sign_out(0);
    CN25_data_in(26) <= VN1766_data_out(0);
    CN25_sign_in(26) <= VN1766_sign_out(0);
    CN25_data_in(27) <= VN1800_data_out(0);
    CN25_sign_in(27) <= VN1800_sign_out(0);
    CN25_data_in(28) <= VN1841_data_out(0);
    CN25_sign_in(28) <= VN1841_sign_out(0);
    CN25_data_in(29) <= VN1862_data_out(0);
    CN25_sign_in(29) <= VN1862_sign_out(0);
    CN25_data_in(30) <= VN1875_data_out(0);
    CN25_sign_in(30) <= VN1875_sign_out(0);
    CN25_data_in(31) <= VN1877_data_out(0);
    CN25_sign_in(31) <= VN1877_sign_out(0);
    CN26_data_in(0) <= VN28_data_out(0);
    CN26_sign_in(0) <= VN28_sign_out(0);
    CN26_data_in(1) <= VN70_data_out(0);
    CN26_sign_in(1) <= VN70_sign_out(0);
    CN26_data_in(2) <= VN116_data_out(0);
    CN26_sign_in(2) <= VN116_sign_out(0);
    CN26_data_in(3) <= VN201_data_out(0);
    CN26_sign_in(3) <= VN201_sign_out(0);
    CN26_data_in(4) <= VN272_data_out(0);
    CN26_sign_in(4) <= VN272_sign_out(0);
    CN26_data_in(5) <= VN286_data_out(0);
    CN26_sign_in(5) <= VN286_sign_out(0);
    CN26_data_in(6) <= VN334_data_out(0);
    CN26_sign_in(6) <= VN334_sign_out(0);
    CN26_data_in(7) <= VN442_data_out(0);
    CN26_sign_in(7) <= VN442_sign_out(0);
    CN26_data_in(8) <= VN453_data_out(0);
    CN26_sign_in(8) <= VN453_sign_out(0);
    CN26_data_in(9) <= VN550_data_out(0);
    CN26_sign_in(9) <= VN550_sign_out(0);
    CN26_data_in(10) <= VN578_data_out(0);
    CN26_sign_in(10) <= VN578_sign_out(0);
    CN26_data_in(11) <= VN649_data_out(0);
    CN26_sign_in(11) <= VN649_sign_out(0);
    CN26_data_in(12) <= VN721_data_out(0);
    CN26_sign_in(12) <= VN721_sign_out(0);
    CN26_data_in(13) <= VN739_data_out(0);
    CN26_sign_in(13) <= VN739_sign_out(0);
    CN26_data_in(14) <= VN829_data_out(0);
    CN26_sign_in(14) <= VN829_sign_out(0);
    CN26_data_in(15) <= VN886_data_out(0);
    CN26_sign_in(15) <= VN886_sign_out(0);
    CN26_data_in(16) <= VN906_data_out(0);
    CN26_sign_in(16) <= VN906_sign_out(0);
    CN26_data_in(17) <= VN966_data_out(0);
    CN26_sign_in(17) <= VN966_sign_out(0);
    CN26_data_in(18) <= VN1058_data_out(0);
    CN26_sign_in(18) <= VN1058_sign_out(0);
    CN26_data_in(19) <= VN1106_data_out(0);
    CN26_sign_in(19) <= VN1106_sign_out(0);
    CN26_data_in(20) <= VN1115_data_out(0);
    CN26_sign_in(20) <= VN1115_sign_out(0);
    CN26_data_in(21) <= VN1179_data_out(0);
    CN26_sign_in(21) <= VN1179_sign_out(0);
    CN26_data_in(22) <= VN1255_data_out(0);
    CN26_sign_in(22) <= VN1255_sign_out(0);
    CN26_data_in(23) <= VN1322_data_out(0);
    CN26_sign_in(23) <= VN1322_sign_out(0);
    CN26_data_in(24) <= VN1364_data_out(0);
    CN26_sign_in(24) <= VN1364_sign_out(0);
    CN26_data_in(25) <= VN1386_data_out(0);
    CN26_sign_in(25) <= VN1386_sign_out(0);
    CN26_data_in(26) <= VN1421_data_out(0);
    CN26_sign_in(26) <= VN1421_sign_out(0);
    CN26_data_in(27) <= VN1465_data_out(0);
    CN26_sign_in(27) <= VN1465_sign_out(0);
    CN26_data_in(28) <= VN1558_data_out(0);
    CN26_sign_in(28) <= VN1558_sign_out(0);
    CN26_data_in(29) <= VN1666_data_out(0);
    CN26_sign_in(29) <= VN1666_sign_out(0);
    CN26_data_in(30) <= VN1694_data_out(0);
    CN26_sign_in(30) <= VN1694_sign_out(0);
    CN26_data_in(31) <= VN1731_data_out(0);
    CN26_sign_in(31) <= VN1731_sign_out(0);
    CN27_data_in(0) <= VN27_data_out(0);
    CN27_sign_in(0) <= VN27_sign_out(0);
    CN27_data_in(1) <= VN69_data_out(0);
    CN27_sign_in(1) <= VN69_sign_out(0);
    CN27_data_in(2) <= VN115_data_out(0);
    CN27_sign_in(2) <= VN115_sign_out(0);
    CN27_data_in(3) <= VN200_data_out(0);
    CN27_sign_in(3) <= VN200_sign_out(0);
    CN27_data_in(4) <= VN285_data_out(0);
    CN27_sign_in(4) <= VN285_sign_out(0);
    CN27_data_in(5) <= VN441_data_out(0);
    CN27_sign_in(5) <= VN441_sign_out(0);
    CN27_data_in(6) <= VN452_data_out(0);
    CN27_sign_in(6) <= VN452_sign_out(0);
    CN27_data_in(7) <= VN549_data_out(0);
    CN27_sign_in(7) <= VN549_sign_out(0);
    CN27_data_in(8) <= VN648_data_out(0);
    CN27_sign_in(8) <= VN648_sign_out(0);
    CN27_data_in(9) <= VN720_data_out(0);
    CN27_sign_in(9) <= VN720_sign_out(0);
    CN27_data_in(10) <= VN738_data_out(0);
    CN27_sign_in(10) <= VN738_sign_out(0);
    CN27_data_in(11) <= VN828_data_out(0);
    CN27_sign_in(11) <= VN828_sign_out(0);
    CN27_data_in(12) <= VN885_data_out(0);
    CN27_sign_in(12) <= VN885_sign_out(0);
    CN27_data_in(13) <= VN905_data_out(0);
    CN27_sign_in(13) <= VN905_sign_out(0);
    CN27_data_in(14) <= VN965_data_out(0);
    CN27_sign_in(14) <= VN965_sign_out(0);
    CN27_data_in(15) <= VN1057_data_out(0);
    CN27_sign_in(15) <= VN1057_sign_out(0);
    CN27_data_in(16) <= VN1105_data_out(0);
    CN27_sign_in(16) <= VN1105_sign_out(0);
    CN27_data_in(17) <= VN1178_data_out(0);
    CN27_sign_in(17) <= VN1178_sign_out(0);
    CN27_data_in(18) <= VN1321_data_out(0);
    CN27_sign_in(18) <= VN1321_sign_out(0);
    CN27_data_in(19) <= VN1385_data_out(0);
    CN27_sign_in(19) <= VN1385_sign_out(0);
    CN27_data_in(20) <= VN1420_data_out(0);
    CN27_sign_in(20) <= VN1420_sign_out(0);
    CN27_data_in(21) <= VN1464_data_out(0);
    CN27_sign_in(21) <= VN1464_sign_out(0);
    CN27_data_in(22) <= VN1557_data_out(0);
    CN27_sign_in(22) <= VN1557_sign_out(0);
    CN27_data_in(23) <= VN1665_data_out(0);
    CN27_sign_in(23) <= VN1665_sign_out(0);
    CN27_data_in(24) <= VN1769_data_out(0);
    CN27_sign_in(24) <= VN1769_sign_out(0);
    CN27_data_in(25) <= VN1780_data_out(0);
    CN27_sign_in(25) <= VN1780_sign_out(0);
    CN27_data_in(26) <= VN1828_data_out(0);
    CN27_sign_in(26) <= VN1828_sign_out(0);
    CN27_data_in(27) <= VN1839_data_out(0);
    CN27_sign_in(27) <= VN1839_sign_out(0);
    CN27_data_in(28) <= VN1848_data_out(0);
    CN27_sign_in(28) <= VN1848_sign_out(0);
    CN27_data_in(29) <= VN1869_data_out(0);
    CN27_sign_in(29) <= VN1869_sign_out(0);
    CN27_data_in(30) <= VN1933_data_out(0);
    CN27_sign_in(30) <= VN1933_sign_out(0);
    CN27_data_in(31) <= VN1935_data_out(0);
    CN27_sign_in(31) <= VN1935_sign_out(0);
    CN28_data_in(0) <= VN26_data_out(0);
    CN28_sign_in(0) <= VN26_sign_out(0);
    CN28_data_in(1) <= VN68_data_out(0);
    CN28_sign_in(1) <= VN68_sign_out(0);
    CN28_data_in(2) <= VN114_data_out(0);
    CN28_sign_in(2) <= VN114_sign_out(0);
    CN28_data_in(3) <= VN199_data_out(0);
    CN28_sign_in(3) <= VN199_sign_out(0);
    CN28_data_in(4) <= VN271_data_out(0);
    CN28_sign_in(4) <= VN271_sign_out(0);
    CN28_data_in(5) <= VN333_data_out(0);
    CN28_sign_in(5) <= VN333_sign_out(0);
    CN28_data_in(6) <= VN440_data_out(0);
    CN28_sign_in(6) <= VN440_sign_out(0);
    CN28_data_in(7) <= VN451_data_out(0);
    CN28_sign_in(7) <= VN451_sign_out(0);
    CN28_data_in(8) <= VN548_data_out(0);
    CN28_sign_in(8) <= VN548_sign_out(0);
    CN28_data_in(9) <= VN577_data_out(0);
    CN28_sign_in(9) <= VN577_sign_out(0);
    CN28_data_in(10) <= VN647_data_out(0);
    CN28_sign_in(10) <= VN647_sign_out(0);
    CN28_data_in(11) <= VN719_data_out(0);
    CN28_sign_in(11) <= VN719_sign_out(0);
    CN28_data_in(12) <= VN737_data_out(0);
    CN28_sign_in(12) <= VN737_sign_out(0);
    CN28_data_in(13) <= VN827_data_out(0);
    CN28_sign_in(13) <= VN827_sign_out(0);
    CN28_data_in(14) <= VN884_data_out(0);
    CN28_sign_in(14) <= VN884_sign_out(0);
    CN28_data_in(15) <= VN904_data_out(0);
    CN28_sign_in(15) <= VN904_sign_out(0);
    CN28_data_in(16) <= VN964_data_out(0);
    CN28_sign_in(16) <= VN964_sign_out(0);
    CN28_data_in(17) <= VN1056_data_out(0);
    CN28_sign_in(17) <= VN1056_sign_out(0);
    CN28_data_in(18) <= VN1104_data_out(0);
    CN28_sign_in(18) <= VN1104_sign_out(0);
    CN28_data_in(19) <= VN1114_data_out(0);
    CN28_sign_in(19) <= VN1114_sign_out(0);
    CN28_data_in(20) <= VN1177_data_out(0);
    CN28_sign_in(20) <= VN1177_sign_out(0);
    CN28_data_in(21) <= VN1254_data_out(0);
    CN28_sign_in(21) <= VN1254_sign_out(0);
    CN28_data_in(22) <= VN1320_data_out(0);
    CN28_sign_in(22) <= VN1320_sign_out(0);
    CN28_data_in(23) <= VN1363_data_out(0);
    CN28_sign_in(23) <= VN1363_sign_out(0);
    CN28_data_in(24) <= VN1384_data_out(0);
    CN28_sign_in(24) <= VN1384_sign_out(0);
    CN28_data_in(25) <= VN1419_data_out(0);
    CN28_sign_in(25) <= VN1419_sign_out(0);
    CN28_data_in(26) <= VN1463_data_out(0);
    CN28_sign_in(26) <= VN1463_sign_out(0);
    CN28_data_in(27) <= VN1556_data_out(0);
    CN28_sign_in(27) <= VN1556_sign_out(0);
    CN28_data_in(28) <= VN1628_data_out(0);
    CN28_sign_in(28) <= VN1628_sign_out(0);
    CN28_data_in(29) <= VN1664_data_out(0);
    CN28_sign_in(29) <= VN1664_sign_out(0);
    CN28_data_in(30) <= VN1693_data_out(0);
    CN28_sign_in(30) <= VN1693_sign_out(0);
    CN28_data_in(31) <= VN1732_data_out(0);
    CN28_sign_in(31) <= VN1732_sign_out(0);
    CN29_data_in(0) <= VN25_data_out(0);
    CN29_sign_in(0) <= VN25_sign_out(0);
    CN29_data_in(1) <= VN67_data_out(0);
    CN29_sign_in(1) <= VN67_sign_out(0);
    CN29_data_in(2) <= VN113_data_out(0);
    CN29_sign_in(2) <= VN113_sign_out(0);
    CN29_data_in(3) <= VN270_data_out(0);
    CN29_sign_in(3) <= VN270_sign_out(0);
    CN29_data_in(4) <= VN450_data_out(0);
    CN29_sign_in(4) <= VN450_sign_out(0);
    CN29_data_in(5) <= VN547_data_out(0);
    CN29_sign_in(5) <= VN547_sign_out(0);
    CN29_data_in(6) <= VN576_data_out(0);
    CN29_sign_in(6) <= VN576_sign_out(0);
    CN29_data_in(7) <= VN646_data_out(0);
    CN29_sign_in(7) <= VN646_sign_out(0);
    CN29_data_in(8) <= VN883_data_out(0);
    CN29_sign_in(8) <= VN883_sign_out(0);
    CN29_data_in(9) <= VN903_data_out(0);
    CN29_sign_in(9) <= VN903_sign_out(0);
    CN29_data_in(10) <= VN1055_data_out(0);
    CN29_sign_in(10) <= VN1055_sign_out(0);
    CN29_data_in(11) <= VN1103_data_out(0);
    CN29_sign_in(11) <= VN1103_sign_out(0);
    CN29_data_in(12) <= VN1253_data_out(0);
    CN29_sign_in(12) <= VN1253_sign_out(0);
    CN29_data_in(13) <= VN1319_data_out(0);
    CN29_sign_in(13) <= VN1319_sign_out(0);
    CN29_data_in(14) <= VN1362_data_out(0);
    CN29_sign_in(14) <= VN1362_sign_out(0);
    CN29_data_in(15) <= VN1418_data_out(0);
    CN29_sign_in(15) <= VN1418_sign_out(0);
    CN29_data_in(16) <= VN1462_data_out(0);
    CN29_sign_in(16) <= VN1462_sign_out(0);
    CN29_data_in(17) <= VN1555_data_out(0);
    CN29_sign_in(17) <= VN1555_sign_out(0);
    CN29_data_in(18) <= VN1627_data_out(0);
    CN29_sign_in(18) <= VN1627_sign_out(0);
    CN29_data_in(19) <= VN1758_data_out(0);
    CN29_sign_in(19) <= VN1758_sign_out(0);
    CN29_data_in(20) <= VN1781_data_out(0);
    CN29_sign_in(20) <= VN1781_sign_out(0);
    CN29_data_in(21) <= VN1803_data_out(0);
    CN29_sign_in(21) <= VN1803_sign_out(0);
    CN29_data_in(22) <= VN1894_data_out(0);
    CN29_sign_in(22) <= VN1894_sign_out(0);
    CN29_data_in(23) <= VN1898_data_out(0);
    CN29_sign_in(23) <= VN1898_sign_out(0);
    CN29_data_in(24) <= VN1913_data_out(0);
    CN29_sign_in(24) <= VN1913_sign_out(0);
    CN29_data_in(25) <= VN1922_data_out(0);
    CN29_sign_in(25) <= VN1922_sign_out(0);
    CN29_data_in(26) <= VN1955_data_out(0);
    CN29_sign_in(26) <= VN1955_sign_out(0);
    CN29_data_in(27) <= VN1960_data_out(0);
    CN29_sign_in(27) <= VN1960_sign_out(0);
    CN29_data_in(28) <= VN1980_data_out(0);
    CN29_sign_in(28) <= VN1980_sign_out(0);
    CN29_data_in(29) <= VN1985_data_out(0);
    CN29_sign_in(29) <= VN1985_sign_out(0);
    CN29_data_in(30) <= VN1988_data_out(0);
    CN29_sign_in(30) <= VN1988_sign_out(0);
    CN29_data_in(31) <= VN1990_data_out(0);
    CN29_sign_in(31) <= VN1990_sign_out(0);
    CN30_data_in(0) <= VN24_data_out(0);
    CN30_sign_in(0) <= VN24_sign_out(0);
    CN30_data_in(1) <= VN66_data_out(0);
    CN30_sign_in(1) <= VN66_sign_out(0);
    CN30_data_in(2) <= VN112_data_out(0);
    CN30_sign_in(2) <= VN112_sign_out(0);
    CN30_data_in(3) <= VN198_data_out(0);
    CN30_sign_in(3) <= VN198_sign_out(0);
    CN30_data_in(4) <= VN269_data_out(0);
    CN30_sign_in(4) <= VN269_sign_out(0);
    CN30_data_in(5) <= VN284_data_out(0);
    CN30_sign_in(5) <= VN284_sign_out(0);
    CN30_data_in(6) <= VN390_data_out(0);
    CN30_sign_in(6) <= VN390_sign_out(0);
    CN30_data_in(7) <= VN439_data_out(0);
    CN30_sign_in(7) <= VN439_sign_out(0);
    CN30_data_in(8) <= VN449_data_out(0);
    CN30_sign_in(8) <= VN449_sign_out(0);
    CN30_data_in(9) <= VN546_data_out(0);
    CN30_sign_in(9) <= VN546_sign_out(0);
    CN30_data_in(10) <= VN575_data_out(0);
    CN30_sign_in(10) <= VN575_sign_out(0);
    CN30_data_in(11) <= VN645_data_out(0);
    CN30_sign_in(11) <= VN645_sign_out(0);
    CN30_data_in(12) <= VN718_data_out(0);
    CN30_sign_in(12) <= VN718_sign_out(0);
    CN30_data_in(13) <= VN736_data_out(0);
    CN30_sign_in(13) <= VN736_sign_out(0);
    CN30_data_in(14) <= VN882_data_out(0);
    CN30_sign_in(14) <= VN882_sign_out(0);
    CN30_data_in(15) <= VN902_data_out(0);
    CN30_sign_in(15) <= VN902_sign_out(0);
    CN30_data_in(16) <= VN963_data_out(0);
    CN30_sign_in(16) <= VN963_sign_out(0);
    CN30_data_in(17) <= VN1054_data_out(0);
    CN30_sign_in(17) <= VN1054_sign_out(0);
    CN30_data_in(18) <= VN1102_data_out(0);
    CN30_sign_in(18) <= VN1102_sign_out(0);
    CN30_data_in(19) <= VN1176_data_out(0);
    CN30_sign_in(19) <= VN1176_sign_out(0);
    CN30_data_in(20) <= VN1252_data_out(0);
    CN30_sign_in(20) <= VN1252_sign_out(0);
    CN30_data_in(21) <= VN1318_data_out(0);
    CN30_sign_in(21) <= VN1318_sign_out(0);
    CN30_data_in(22) <= VN1334_data_out(0);
    CN30_sign_in(22) <= VN1334_sign_out(0);
    CN30_data_in(23) <= VN1361_data_out(0);
    CN30_sign_in(23) <= VN1361_sign_out(0);
    CN30_data_in(24) <= VN1417_data_out(0);
    CN30_sign_in(24) <= VN1417_sign_out(0);
    CN30_data_in(25) <= VN1461_data_out(0);
    CN30_sign_in(25) <= VN1461_sign_out(0);
    CN30_data_in(26) <= VN1513_data_out(0);
    CN30_sign_in(26) <= VN1513_sign_out(0);
    CN30_data_in(27) <= VN1663_data_out(0);
    CN30_sign_in(27) <= VN1663_sign_out(0);
    CN30_data_in(28) <= VN1692_data_out(0);
    CN30_sign_in(28) <= VN1692_sign_out(0);
    CN30_data_in(29) <= VN1771_data_out(0);
    CN30_sign_in(29) <= VN1771_sign_out(0);
    CN30_data_in(30) <= VN1806_data_out(0);
    CN30_sign_in(30) <= VN1806_sign_out(0);
    CN30_data_in(31) <= VN1815_data_out(0);
    CN30_sign_in(31) <= VN1815_sign_out(0);
    CN31_data_in(0) <= VN23_data_out(0);
    CN31_sign_in(0) <= VN23_sign_out(0);
    CN31_data_in(1) <= VN65_data_out(0);
    CN31_sign_in(1) <= VN65_sign_out(0);
    CN31_data_in(2) <= VN197_data_out(0);
    CN31_sign_in(2) <= VN197_sign_out(0);
    CN31_data_in(3) <= VN283_data_out(0);
    CN31_sign_in(3) <= VN283_sign_out(0);
    CN31_data_in(4) <= VN389_data_out(0);
    CN31_sign_in(4) <= VN389_sign_out(0);
    CN31_data_in(5) <= VN438_data_out(0);
    CN31_sign_in(5) <= VN438_sign_out(0);
    CN31_data_in(6) <= VN448_data_out(0);
    CN31_sign_in(6) <= VN448_sign_out(0);
    CN31_data_in(7) <= VN545_data_out(0);
    CN31_sign_in(7) <= VN545_sign_out(0);
    CN31_data_in(8) <= VN574_data_out(0);
    CN31_sign_in(8) <= VN574_sign_out(0);
    CN31_data_in(9) <= VN644_data_out(0);
    CN31_sign_in(9) <= VN644_sign_out(0);
    CN31_data_in(10) <= VN717_data_out(0);
    CN31_sign_in(10) <= VN717_sign_out(0);
    CN31_data_in(11) <= VN735_data_out(0);
    CN31_sign_in(11) <= VN735_sign_out(0);
    CN31_data_in(12) <= VN826_data_out(0);
    CN31_sign_in(12) <= VN826_sign_out(0);
    CN31_data_in(13) <= VN881_data_out(0);
    CN31_sign_in(13) <= VN881_sign_out(0);
    CN31_data_in(14) <= VN901_data_out(0);
    CN31_sign_in(14) <= VN901_sign_out(0);
    CN31_data_in(15) <= VN962_data_out(0);
    CN31_sign_in(15) <= VN962_sign_out(0);
    CN31_data_in(16) <= VN1053_data_out(0);
    CN31_sign_in(16) <= VN1053_sign_out(0);
    CN31_data_in(17) <= VN1101_data_out(0);
    CN31_sign_in(17) <= VN1101_sign_out(0);
    CN31_data_in(18) <= VN1175_data_out(0);
    CN31_sign_in(18) <= VN1175_sign_out(0);
    CN31_data_in(19) <= VN1251_data_out(0);
    CN31_sign_in(19) <= VN1251_sign_out(0);
    CN31_data_in(20) <= VN1317_data_out(0);
    CN31_sign_in(20) <= VN1317_sign_out(0);
    CN31_data_in(21) <= VN1333_data_out(0);
    CN31_sign_in(21) <= VN1333_sign_out(0);
    CN31_data_in(22) <= VN1360_data_out(0);
    CN31_sign_in(22) <= VN1360_sign_out(0);
    CN31_data_in(23) <= VN1416_data_out(0);
    CN31_sign_in(23) <= VN1416_sign_out(0);
    CN31_data_in(24) <= VN1460_data_out(0);
    CN31_sign_in(24) <= VN1460_sign_out(0);
    CN31_data_in(25) <= VN1554_data_out(0);
    CN31_sign_in(25) <= VN1554_sign_out(0);
    CN31_data_in(26) <= VN1626_data_out(0);
    CN31_sign_in(26) <= VN1626_sign_out(0);
    CN31_data_in(27) <= VN1782_data_out(0);
    CN31_sign_in(27) <= VN1782_sign_out(0);
    CN31_data_in(28) <= VN1790_data_out(0);
    CN31_sign_in(28) <= VN1790_sign_out(0);
    CN31_data_in(29) <= VN1921_data_out(0);
    CN31_sign_in(29) <= VN1921_sign_out(0);
    CN31_data_in(30) <= VN1952_data_out(0);
    CN31_sign_in(30) <= VN1952_sign_out(0);
    CN31_data_in(31) <= VN1962_data_out(0);
    CN31_sign_in(31) <= VN1962_sign_out(0);
    CN32_data_in(0) <= VN22_data_out(0);
    CN32_sign_in(0) <= VN22_sign_out(0);
    CN32_data_in(1) <= VN64_data_out(0);
    CN32_sign_in(1) <= VN64_sign_out(0);
    CN32_data_in(2) <= VN111_data_out(0);
    CN32_sign_in(2) <= VN111_sign_out(0);
    CN32_data_in(3) <= VN268_data_out(0);
    CN32_sign_in(3) <= VN268_sign_out(0);
    CN32_data_in(4) <= VN388_data_out(0);
    CN32_sign_in(4) <= VN388_sign_out(0);
    CN32_data_in(5) <= VN504_data_out(0);
    CN32_sign_in(5) <= VN504_sign_out(0);
    CN32_data_in(6) <= VN544_data_out(0);
    CN32_sign_in(6) <= VN544_sign_out(0);
    CN32_data_in(7) <= VN573_data_out(0);
    CN32_sign_in(7) <= VN573_sign_out(0);
    CN32_data_in(8) <= VN643_data_out(0);
    CN32_sign_in(8) <= VN643_sign_out(0);
    CN32_data_in(9) <= VN734_data_out(0);
    CN32_sign_in(9) <= VN734_sign_out(0);
    CN32_data_in(10) <= VN825_data_out(0);
    CN32_sign_in(10) <= VN825_sign_out(0);
    CN32_data_in(11) <= VN880_data_out(0);
    CN32_sign_in(11) <= VN880_sign_out(0);
    CN32_data_in(12) <= VN900_data_out(0);
    CN32_sign_in(12) <= VN900_sign_out(0);
    CN32_data_in(13) <= VN961_data_out(0);
    CN32_sign_in(13) <= VN961_sign_out(0);
    CN32_data_in(14) <= VN1052_data_out(0);
    CN32_sign_in(14) <= VN1052_sign_out(0);
    CN32_data_in(15) <= VN1250_data_out(0);
    CN32_sign_in(15) <= VN1250_sign_out(0);
    CN32_data_in(16) <= VN1316_data_out(0);
    CN32_sign_in(16) <= VN1316_sign_out(0);
    CN32_data_in(17) <= VN1359_data_out(0);
    CN32_sign_in(17) <= VN1359_sign_out(0);
    CN32_data_in(18) <= VN1459_data_out(0);
    CN32_sign_in(18) <= VN1459_sign_out(0);
    CN32_data_in(19) <= VN1662_data_out(0);
    CN32_sign_in(19) <= VN1662_sign_out(0);
    CN32_data_in(20) <= VN1691_data_out(0);
    CN32_sign_in(20) <= VN1691_sign_out(0);
    CN32_data_in(21) <= VN1742_data_out(0);
    CN32_sign_in(21) <= VN1742_sign_out(0);
    CN32_data_in(22) <= VN1826_data_out(0);
    CN32_sign_in(22) <= VN1826_sign_out(0);
    CN32_data_in(23) <= VN1831_data_out(0);
    CN32_sign_in(23) <= VN1831_sign_out(0);
    CN32_data_in(24) <= VN1943_data_out(0);
    CN32_sign_in(24) <= VN1943_sign_out(0);
    CN32_data_in(25) <= VN1958_data_out(0);
    CN32_sign_in(25) <= VN1958_sign_out(0);
    CN32_data_in(26) <= VN1959_data_out(0);
    CN32_sign_in(26) <= VN1959_sign_out(0);
    CN32_data_in(27) <= VN1973_data_out(0);
    CN32_sign_in(27) <= VN1973_sign_out(0);
    CN32_data_in(28) <= VN1999_data_out(0);
    CN32_sign_in(28) <= VN1999_sign_out(0);
    CN32_data_in(29) <= VN2008_data_out(0);
    CN32_sign_in(29) <= VN2008_sign_out(0);
    CN32_data_in(30) <= VN2027_data_out(0);
    CN32_sign_in(30) <= VN2027_sign_out(0);
    CN32_data_in(31) <= VN2029_data_out(0);
    CN32_sign_in(31) <= VN2029_sign_out(0);
    CN33_data_in(0) <= VN21_data_out(0);
    CN33_sign_in(0) <= VN21_sign_out(0);
    CN33_data_in(1) <= VN63_data_out(0);
    CN33_sign_in(1) <= VN63_sign_out(0);
    CN33_data_in(2) <= VN169_data_out(0);
    CN33_sign_in(2) <= VN169_sign_out(0);
    CN33_data_in(3) <= VN196_data_out(0);
    CN33_sign_in(3) <= VN196_sign_out(0);
    CN33_data_in(4) <= VN267_data_out(0);
    CN33_sign_in(4) <= VN267_sign_out(0);
    CN33_data_in(5) <= VN282_data_out(0);
    CN33_sign_in(5) <= VN282_sign_out(0);
    CN33_data_in(6) <= VN387_data_out(0);
    CN33_sign_in(6) <= VN387_sign_out(0);
    CN33_data_in(7) <= VN437_data_out(0);
    CN33_sign_in(7) <= VN437_sign_out(0);
    CN33_data_in(8) <= VN503_data_out(0);
    CN33_sign_in(8) <= VN503_sign_out(0);
    CN33_data_in(9) <= VN543_data_out(0);
    CN33_sign_in(9) <= VN543_sign_out(0);
    CN33_data_in(10) <= VN572_data_out(0);
    CN33_sign_in(10) <= VN572_sign_out(0);
    CN33_data_in(11) <= VN642_data_out(0);
    CN33_sign_in(11) <= VN642_sign_out(0);
    CN33_data_in(12) <= VN716_data_out(0);
    CN33_sign_in(12) <= VN716_sign_out(0);
    CN33_data_in(13) <= VN733_data_out(0);
    CN33_sign_in(13) <= VN733_sign_out(0);
    CN33_data_in(14) <= VN824_data_out(0);
    CN33_sign_in(14) <= VN824_sign_out(0);
    CN33_data_in(15) <= VN879_data_out(0);
    CN33_sign_in(15) <= VN879_sign_out(0);
    CN33_data_in(16) <= VN899_data_out(0);
    CN33_sign_in(16) <= VN899_sign_out(0);
    CN33_data_in(17) <= VN960_data_out(0);
    CN33_sign_in(17) <= VN960_sign_out(0);
    CN33_data_in(18) <= VN1051_data_out(0);
    CN33_sign_in(18) <= VN1051_sign_out(0);
    CN33_data_in(19) <= VN1100_data_out(0);
    CN33_sign_in(19) <= VN1100_sign_out(0);
    CN33_data_in(20) <= VN1174_data_out(0);
    CN33_sign_in(20) <= VN1174_sign_out(0);
    CN33_data_in(21) <= VN1249_data_out(0);
    CN33_sign_in(21) <= VN1249_sign_out(0);
    CN33_data_in(22) <= VN1315_data_out(0);
    CN33_sign_in(22) <= VN1315_sign_out(0);
    CN33_data_in(23) <= VN1332_data_out(0);
    CN33_sign_in(23) <= VN1332_sign_out(0);
    CN33_data_in(24) <= VN1358_data_out(0);
    CN33_sign_in(24) <= VN1358_sign_out(0);
    CN33_data_in(25) <= VN1415_data_out(0);
    CN33_sign_in(25) <= VN1415_sign_out(0);
    CN33_data_in(26) <= VN1458_data_out(0);
    CN33_sign_in(26) <= VN1458_sign_out(0);
    CN33_data_in(27) <= VN1512_data_out(0);
    CN33_sign_in(27) <= VN1512_sign_out(0);
    CN33_data_in(28) <= VN1574_data_out(0);
    CN33_sign_in(28) <= VN1574_sign_out(0);
    CN33_data_in(29) <= VN1625_data_out(0);
    CN33_sign_in(29) <= VN1625_sign_out(0);
    CN33_data_in(30) <= VN1690_data_out(0);
    CN33_sign_in(30) <= VN1690_sign_out(0);
    CN33_data_in(31) <= VN1733_data_out(0);
    CN33_sign_in(31) <= VN1733_sign_out(0);
    CN34_data_in(0) <= VN20_data_out(0);
    CN34_sign_in(0) <= VN20_sign_out(0);
    CN34_data_in(1) <= VN62_data_out(0);
    CN34_sign_in(1) <= VN62_sign_out(0);
    CN34_data_in(2) <= VN168_data_out(0);
    CN34_sign_in(2) <= VN168_sign_out(0);
    CN34_data_in(3) <= VN195_data_out(0);
    CN34_sign_in(3) <= VN195_sign_out(0);
    CN34_data_in(4) <= VN266_data_out(0);
    CN34_sign_in(4) <= VN266_sign_out(0);
    CN34_data_in(5) <= VN281_data_out(0);
    CN34_sign_in(5) <= VN281_sign_out(0);
    CN34_data_in(6) <= VN386_data_out(0);
    CN34_sign_in(6) <= VN386_sign_out(0);
    CN34_data_in(7) <= VN436_data_out(0);
    CN34_sign_in(7) <= VN436_sign_out(0);
    CN34_data_in(8) <= VN502_data_out(0);
    CN34_sign_in(8) <= VN502_sign_out(0);
    CN34_data_in(9) <= VN542_data_out(0);
    CN34_sign_in(9) <= VN542_sign_out(0);
    CN34_data_in(10) <= VN571_data_out(0);
    CN34_sign_in(10) <= VN571_sign_out(0);
    CN34_data_in(11) <= VN641_data_out(0);
    CN34_sign_in(11) <= VN641_sign_out(0);
    CN34_data_in(12) <= VN715_data_out(0);
    CN34_sign_in(12) <= VN715_sign_out(0);
    CN34_data_in(13) <= VN732_data_out(0);
    CN34_sign_in(13) <= VN732_sign_out(0);
    CN34_data_in(14) <= VN823_data_out(0);
    CN34_sign_in(14) <= VN823_sign_out(0);
    CN34_data_in(15) <= VN878_data_out(0);
    CN34_sign_in(15) <= VN878_sign_out(0);
    CN34_data_in(16) <= VN898_data_out(0);
    CN34_sign_in(16) <= VN898_sign_out(0);
    CN34_data_in(17) <= VN959_data_out(0);
    CN34_sign_in(17) <= VN959_sign_out(0);
    CN34_data_in(18) <= VN1050_data_out(0);
    CN34_sign_in(18) <= VN1050_sign_out(0);
    CN34_data_in(19) <= VN1099_data_out(0);
    CN34_sign_in(19) <= VN1099_sign_out(0);
    CN34_data_in(20) <= VN1173_data_out(0);
    CN34_sign_in(20) <= VN1173_sign_out(0);
    CN34_data_in(21) <= VN1248_data_out(0);
    CN34_sign_in(21) <= VN1248_sign_out(0);
    CN34_data_in(22) <= VN1314_data_out(0);
    CN34_sign_in(22) <= VN1314_sign_out(0);
    CN34_data_in(23) <= VN1331_data_out(0);
    CN34_sign_in(23) <= VN1331_sign_out(0);
    CN34_data_in(24) <= VN1414_data_out(0);
    CN34_sign_in(24) <= VN1414_sign_out(0);
    CN34_data_in(25) <= VN1511_data_out(0);
    CN34_sign_in(25) <= VN1511_sign_out(0);
    CN34_data_in(26) <= VN1573_data_out(0);
    CN34_sign_in(26) <= VN1573_sign_out(0);
    CN34_data_in(27) <= VN1606_data_out(0);
    CN34_sign_in(27) <= VN1606_sign_out(0);
    CN34_data_in(28) <= VN1624_data_out(0);
    CN34_sign_in(28) <= VN1624_sign_out(0);
    CN34_data_in(29) <= VN1661_data_out(0);
    CN34_sign_in(29) <= VN1661_sign_out(0);
    CN34_data_in(30) <= VN1822_data_out(0);
    CN34_sign_in(30) <= VN1822_sign_out(0);
    CN34_data_in(31) <= VN1878_data_out(0);
    CN34_sign_in(31) <= VN1878_sign_out(0);
    CN35_data_in(0) <= VN19_data_out(0);
    CN35_sign_in(0) <= VN19_sign_out(0);
    CN35_data_in(1) <= VN61_data_out(0);
    CN35_sign_in(1) <= VN61_sign_out(0);
    CN35_data_in(2) <= VN167_data_out(0);
    CN35_sign_in(2) <= VN167_sign_out(0);
    CN35_data_in(3) <= VN194_data_out(0);
    CN35_sign_in(3) <= VN194_sign_out(0);
    CN35_data_in(4) <= VN265_data_out(0);
    CN35_sign_in(4) <= VN265_sign_out(0);
    CN35_data_in(5) <= VN280_data_out(0);
    CN35_sign_in(5) <= VN280_sign_out(0);
    CN35_data_in(6) <= VN385_data_out(0);
    CN35_sign_in(6) <= VN385_sign_out(0);
    CN35_data_in(7) <= VN435_data_out(0);
    CN35_sign_in(7) <= VN435_sign_out(0);
    CN35_data_in(8) <= VN501_data_out(0);
    CN35_sign_in(8) <= VN501_sign_out(0);
    CN35_data_in(9) <= VN541_data_out(0);
    CN35_sign_in(9) <= VN541_sign_out(0);
    CN35_data_in(10) <= VN570_data_out(0);
    CN35_sign_in(10) <= VN570_sign_out(0);
    CN35_data_in(11) <= VN640_data_out(0);
    CN35_sign_in(11) <= VN640_sign_out(0);
    CN35_data_in(12) <= VN714_data_out(0);
    CN35_sign_in(12) <= VN714_sign_out(0);
    CN35_data_in(13) <= VN731_data_out(0);
    CN35_sign_in(13) <= VN731_sign_out(0);
    CN35_data_in(14) <= VN822_data_out(0);
    CN35_sign_in(14) <= VN822_sign_out(0);
    CN35_data_in(15) <= VN877_data_out(0);
    CN35_sign_in(15) <= VN877_sign_out(0);
    CN35_data_in(16) <= VN897_data_out(0);
    CN35_sign_in(16) <= VN897_sign_out(0);
    CN35_data_in(17) <= VN958_data_out(0);
    CN35_sign_in(17) <= VN958_sign_out(0);
    CN35_data_in(18) <= VN1049_data_out(0);
    CN35_sign_in(18) <= VN1049_sign_out(0);
    CN35_data_in(19) <= VN1098_data_out(0);
    CN35_sign_in(19) <= VN1098_sign_out(0);
    CN35_data_in(20) <= VN1172_data_out(0);
    CN35_sign_in(20) <= VN1172_sign_out(0);
    CN35_data_in(21) <= VN1247_data_out(0);
    CN35_sign_in(21) <= VN1247_sign_out(0);
    CN35_data_in(22) <= VN1313_data_out(0);
    CN35_sign_in(22) <= VN1313_sign_out(0);
    CN35_data_in(23) <= VN1330_data_out(0);
    CN35_sign_in(23) <= VN1330_sign_out(0);
    CN35_data_in(24) <= VN1357_data_out(0);
    CN35_sign_in(24) <= VN1357_sign_out(0);
    CN35_data_in(25) <= VN1413_data_out(0);
    CN35_sign_in(25) <= VN1413_sign_out(0);
    CN35_data_in(26) <= VN1510_data_out(0);
    CN35_sign_in(26) <= VN1510_sign_out(0);
    CN35_data_in(27) <= VN1605_data_out(0);
    CN35_sign_in(27) <= VN1605_sign_out(0);
    CN35_data_in(28) <= VN1623_data_out(0);
    CN35_sign_in(28) <= VN1623_sign_out(0);
    CN35_data_in(29) <= VN1660_data_out(0);
    CN35_sign_in(29) <= VN1660_sign_out(0);
    CN35_data_in(30) <= VN1689_data_out(0);
    CN35_sign_in(30) <= VN1689_sign_out(0);
    CN35_data_in(31) <= VN1734_data_out(0);
    CN35_sign_in(31) <= VN1734_sign_out(0);
    CN36_data_in(0) <= VN18_data_out(0);
    CN36_sign_in(0) <= VN18_sign_out(0);
    CN36_data_in(1) <= VN60_data_out(0);
    CN36_sign_in(1) <= VN60_sign_out(0);
    CN36_data_in(2) <= VN166_data_out(0);
    CN36_sign_in(2) <= VN166_sign_out(0);
    CN36_data_in(3) <= VN264_data_out(0);
    CN36_sign_in(3) <= VN264_sign_out(0);
    CN36_data_in(4) <= VN384_data_out(0);
    CN36_sign_in(4) <= VN384_sign_out(0);
    CN36_data_in(5) <= VN434_data_out(0);
    CN36_sign_in(5) <= VN434_sign_out(0);
    CN36_data_in(6) <= VN500_data_out(0);
    CN36_sign_in(6) <= VN500_sign_out(0);
    CN36_data_in(7) <= VN540_data_out(0);
    CN36_sign_in(7) <= VN540_sign_out(0);
    CN36_data_in(8) <= VN639_data_out(0);
    CN36_sign_in(8) <= VN639_sign_out(0);
    CN36_data_in(9) <= VN821_data_out(0);
    CN36_sign_in(9) <= VN821_sign_out(0);
    CN36_data_in(10) <= VN896_data_out(0);
    CN36_sign_in(10) <= VN896_sign_out(0);
    CN36_data_in(11) <= VN957_data_out(0);
    CN36_sign_in(11) <= VN957_sign_out(0);
    CN36_data_in(12) <= VN1048_data_out(0);
    CN36_sign_in(12) <= VN1048_sign_out(0);
    CN36_data_in(13) <= VN1171_data_out(0);
    CN36_sign_in(13) <= VN1171_sign_out(0);
    CN36_data_in(14) <= VN1246_data_out(0);
    CN36_sign_in(14) <= VN1246_sign_out(0);
    CN36_data_in(15) <= VN1329_data_out(0);
    CN36_sign_in(15) <= VN1329_sign_out(0);
    CN36_data_in(16) <= VN1356_data_out(0);
    CN36_sign_in(16) <= VN1356_sign_out(0);
    CN36_data_in(17) <= VN1412_data_out(0);
    CN36_sign_in(17) <= VN1412_sign_out(0);
    CN36_data_in(18) <= VN1604_data_out(0);
    CN36_sign_in(18) <= VN1604_sign_out(0);
    CN36_data_in(19) <= VN1622_data_out(0);
    CN36_sign_in(19) <= VN1622_sign_out(0);
    CN36_data_in(20) <= VN1659_data_out(0);
    CN36_sign_in(20) <= VN1659_sign_out(0);
    CN36_data_in(21) <= VN1743_data_out(0);
    CN36_sign_in(21) <= VN1743_sign_out(0);
    CN36_data_in(22) <= VN1873_data_out(0);
    CN36_sign_in(22) <= VN1873_sign_out(0);
    CN36_data_in(23) <= VN1888_data_out(0);
    CN36_sign_in(23) <= VN1888_sign_out(0);
    CN36_data_in(24) <= VN1947_data_out(0);
    CN36_sign_in(24) <= VN1947_sign_out(0);
    CN36_data_in(25) <= VN1950_data_out(0);
    CN36_sign_in(25) <= VN1950_sign_out(0);
    CN36_data_in(26) <= VN1969_data_out(0);
    CN36_sign_in(26) <= VN1969_sign_out(0);
    CN36_data_in(27) <= VN1976_data_out(0);
    CN36_sign_in(27) <= VN1976_sign_out(0);
    CN36_data_in(28) <= VN1995_data_out(0);
    CN36_sign_in(28) <= VN1995_sign_out(0);
    CN36_data_in(29) <= VN2002_data_out(0);
    CN36_sign_in(29) <= VN2002_sign_out(0);
    CN36_data_in(30) <= VN2022_data_out(0);
    CN36_sign_in(30) <= VN2022_sign_out(0);
    CN36_data_in(31) <= VN2030_data_out(0);
    CN36_sign_in(31) <= VN2030_sign_out(0);
    CN37_data_in(0) <= VN17_data_out(0);
    CN37_sign_in(0) <= VN17_sign_out(0);
    CN37_data_in(1) <= VN59_data_out(0);
    CN37_sign_in(1) <= VN59_sign_out(0);
    CN37_data_in(2) <= VN165_data_out(0);
    CN37_sign_in(2) <= VN165_sign_out(0);
    CN37_data_in(3) <= VN193_data_out(0);
    CN37_sign_in(3) <= VN193_sign_out(0);
    CN37_data_in(4) <= VN263_data_out(0);
    CN37_sign_in(4) <= VN263_sign_out(0);
    CN37_data_in(5) <= VN331_data_out(0);
    CN37_sign_in(5) <= VN331_sign_out(0);
    CN37_data_in(6) <= VN383_data_out(0);
    CN37_sign_in(6) <= VN383_sign_out(0);
    CN37_data_in(7) <= VN433_data_out(0);
    CN37_sign_in(7) <= VN433_sign_out(0);
    CN37_data_in(8) <= VN499_data_out(0);
    CN37_sign_in(8) <= VN499_sign_out(0);
    CN37_data_in(9) <= VN539_data_out(0);
    CN37_sign_in(9) <= VN539_sign_out(0);
    CN37_data_in(10) <= VN569_data_out(0);
    CN37_sign_in(10) <= VN569_sign_out(0);
    CN37_data_in(11) <= VN638_data_out(0);
    CN37_sign_in(11) <= VN638_sign_out(0);
    CN37_data_in(12) <= VN713_data_out(0);
    CN37_sign_in(12) <= VN713_sign_out(0);
    CN37_data_in(13) <= VN730_data_out(0);
    CN37_sign_in(13) <= VN730_sign_out(0);
    CN37_data_in(14) <= VN820_data_out(0);
    CN37_sign_in(14) <= VN820_sign_out(0);
    CN37_data_in(15) <= VN876_data_out(0);
    CN37_sign_in(15) <= VN876_sign_out(0);
    CN37_data_in(16) <= VN895_data_out(0);
    CN37_sign_in(16) <= VN895_sign_out(0);
    CN37_data_in(17) <= VN956_data_out(0);
    CN37_sign_in(17) <= VN956_sign_out(0);
    CN37_data_in(18) <= VN1047_data_out(0);
    CN37_sign_in(18) <= VN1047_sign_out(0);
    CN37_data_in(19) <= VN1097_data_out(0);
    CN37_sign_in(19) <= VN1097_sign_out(0);
    CN37_data_in(20) <= VN1163_data_out(0);
    CN37_sign_in(20) <= VN1163_sign_out(0);
    CN37_data_in(21) <= VN1170_data_out(0);
    CN37_sign_in(21) <= VN1170_sign_out(0);
    CN37_data_in(22) <= VN1245_data_out(0);
    CN37_sign_in(22) <= VN1245_sign_out(0);
    CN37_data_in(23) <= VN1282_data_out(0);
    CN37_sign_in(23) <= VN1282_sign_out(0);
    CN37_data_in(24) <= VN1312_data_out(0);
    CN37_sign_in(24) <= VN1312_sign_out(0);
    CN37_data_in(25) <= VN1355_data_out(0);
    CN37_sign_in(25) <= VN1355_sign_out(0);
    CN37_data_in(26) <= VN1572_data_out(0);
    CN37_sign_in(26) <= VN1572_sign_out(0);
    CN37_data_in(27) <= VN1603_data_out(0);
    CN37_sign_in(27) <= VN1603_sign_out(0);
    CN37_data_in(28) <= VN1621_data_out(0);
    CN37_sign_in(28) <= VN1621_sign_out(0);
    CN37_data_in(29) <= VN1658_data_out(0);
    CN37_sign_in(29) <= VN1658_sign_out(0);
    CN37_data_in(30) <= VN1688_data_out(0);
    CN37_sign_in(30) <= VN1688_sign_out(0);
    CN37_data_in(31) <= VN1735_data_out(0);
    CN37_sign_in(31) <= VN1735_sign_out(0);
    CN38_data_in(0) <= VN16_data_out(0);
    CN38_sign_in(0) <= VN16_sign_out(0);
    CN38_data_in(1) <= VN58_data_out(0);
    CN38_sign_in(1) <= VN58_sign_out(0);
    CN38_data_in(2) <= VN164_data_out(0);
    CN38_sign_in(2) <= VN164_sign_out(0);
    CN38_data_in(3) <= VN192_data_out(0);
    CN38_sign_in(3) <= VN192_sign_out(0);
    CN38_data_in(4) <= VN262_data_out(0);
    CN38_sign_in(4) <= VN262_sign_out(0);
    CN38_data_in(5) <= VN330_data_out(0);
    CN38_sign_in(5) <= VN330_sign_out(0);
    CN38_data_in(6) <= VN382_data_out(0);
    CN38_sign_in(6) <= VN382_sign_out(0);
    CN38_data_in(7) <= VN432_data_out(0);
    CN38_sign_in(7) <= VN432_sign_out(0);
    CN38_data_in(8) <= VN498_data_out(0);
    CN38_sign_in(8) <= VN498_sign_out(0);
    CN38_data_in(9) <= VN538_data_out(0);
    CN38_sign_in(9) <= VN538_sign_out(0);
    CN38_data_in(10) <= VN568_data_out(0);
    CN38_sign_in(10) <= VN568_sign_out(0);
    CN38_data_in(11) <= VN637_data_out(0);
    CN38_sign_in(11) <= VN637_sign_out(0);
    CN38_data_in(12) <= VN712_data_out(0);
    CN38_sign_in(12) <= VN712_sign_out(0);
    CN38_data_in(13) <= VN729_data_out(0);
    CN38_sign_in(13) <= VN729_sign_out(0);
    CN38_data_in(14) <= VN875_data_out(0);
    CN38_sign_in(14) <= VN875_sign_out(0);
    CN38_data_in(15) <= VN894_data_out(0);
    CN38_sign_in(15) <= VN894_sign_out(0);
    CN38_data_in(16) <= VN955_data_out(0);
    CN38_sign_in(16) <= VN955_sign_out(0);
    CN38_data_in(17) <= VN1046_data_out(0);
    CN38_sign_in(17) <= VN1046_sign_out(0);
    CN38_data_in(18) <= VN1096_data_out(0);
    CN38_sign_in(18) <= VN1096_sign_out(0);
    CN38_data_in(19) <= VN1162_data_out(0);
    CN38_sign_in(19) <= VN1162_sign_out(0);
    CN38_data_in(20) <= VN1244_data_out(0);
    CN38_sign_in(20) <= VN1244_sign_out(0);
    CN38_data_in(21) <= VN1281_data_out(0);
    CN38_sign_in(21) <= VN1281_sign_out(0);
    CN38_data_in(22) <= VN1311_data_out(0);
    CN38_sign_in(22) <= VN1311_sign_out(0);
    CN38_data_in(23) <= VN1411_data_out(0);
    CN38_sign_in(23) <= VN1411_sign_out(0);
    CN38_data_in(24) <= VN1518_data_out(0);
    CN38_sign_in(24) <= VN1518_sign_out(0);
    CN38_data_in(25) <= VN1571_data_out(0);
    CN38_sign_in(25) <= VN1571_sign_out(0);
    CN38_data_in(26) <= VN1620_data_out(0);
    CN38_sign_in(26) <= VN1620_sign_out(0);
    CN38_data_in(27) <= VN1767_data_out(0);
    CN38_sign_in(27) <= VN1767_sign_out(0);
    CN38_data_in(28) <= VN1881_data_out(0);
    CN38_sign_in(28) <= VN1881_sign_out(0);
    CN38_data_in(29) <= VN1897_data_out(0);
    CN38_sign_in(29) <= VN1897_sign_out(0);
    CN38_data_in(30) <= VN1909_data_out(0);
    CN38_sign_in(30) <= VN1909_sign_out(0);
    CN38_data_in(31) <= VN1915_data_out(0);
    CN38_sign_in(31) <= VN1915_sign_out(0);
    CN39_data_in(0) <= VN15_data_out(0);
    CN39_sign_in(0) <= VN15_sign_out(0);
    CN39_data_in(1) <= VN57_data_out(0);
    CN39_sign_in(1) <= VN57_sign_out(0);
    CN39_data_in(2) <= VN163_data_out(0);
    CN39_sign_in(2) <= VN163_sign_out(0);
    CN39_data_in(3) <= VN191_data_out(0);
    CN39_sign_in(3) <= VN191_sign_out(0);
    CN39_data_in(4) <= VN261_data_out(0);
    CN39_sign_in(4) <= VN261_sign_out(0);
    CN39_data_in(5) <= VN329_data_out(0);
    CN39_sign_in(5) <= VN329_sign_out(0);
    CN39_data_in(6) <= VN381_data_out(0);
    CN39_sign_in(6) <= VN381_sign_out(0);
    CN39_data_in(7) <= VN431_data_out(0);
    CN39_sign_in(7) <= VN431_sign_out(0);
    CN39_data_in(8) <= VN497_data_out(0);
    CN39_sign_in(8) <= VN497_sign_out(0);
    CN39_data_in(9) <= VN537_data_out(0);
    CN39_sign_in(9) <= VN537_sign_out(0);
    CN39_data_in(10) <= VN567_data_out(0);
    CN39_sign_in(10) <= VN567_sign_out(0);
    CN39_data_in(11) <= VN636_data_out(0);
    CN39_sign_in(11) <= VN636_sign_out(0);
    CN39_data_in(12) <= VN711_data_out(0);
    CN39_sign_in(12) <= VN711_sign_out(0);
    CN39_data_in(13) <= VN728_data_out(0);
    CN39_sign_in(13) <= VN728_sign_out(0);
    CN39_data_in(14) <= VN819_data_out(0);
    CN39_sign_in(14) <= VN819_sign_out(0);
    CN39_data_in(15) <= VN874_data_out(0);
    CN39_sign_in(15) <= VN874_sign_out(0);
    CN39_data_in(16) <= VN893_data_out(0);
    CN39_sign_in(16) <= VN893_sign_out(0);
    CN39_data_in(17) <= VN954_data_out(0);
    CN39_sign_in(17) <= VN954_sign_out(0);
    CN39_data_in(18) <= VN1045_data_out(0);
    CN39_sign_in(18) <= VN1045_sign_out(0);
    CN39_data_in(19) <= VN1095_data_out(0);
    CN39_sign_in(19) <= VN1095_sign_out(0);
    CN39_data_in(20) <= VN1161_data_out(0);
    CN39_sign_in(20) <= VN1161_sign_out(0);
    CN39_data_in(21) <= VN1243_data_out(0);
    CN39_sign_in(21) <= VN1243_sign_out(0);
    CN39_data_in(22) <= VN1280_data_out(0);
    CN39_sign_in(22) <= VN1280_sign_out(0);
    CN39_data_in(23) <= VN1310_data_out(0);
    CN39_sign_in(23) <= VN1310_sign_out(0);
    CN39_data_in(24) <= VN1354_data_out(0);
    CN39_sign_in(24) <= VN1354_sign_out(0);
    CN39_data_in(25) <= VN1410_data_out(0);
    CN39_sign_in(25) <= VN1410_sign_out(0);
    CN39_data_in(26) <= VN1517_data_out(0);
    CN39_sign_in(26) <= VN1517_sign_out(0);
    CN39_data_in(27) <= VN1570_data_out(0);
    CN39_sign_in(27) <= VN1570_sign_out(0);
    CN39_data_in(28) <= VN1602_data_out(0);
    CN39_sign_in(28) <= VN1602_sign_out(0);
    CN39_data_in(29) <= VN1619_data_out(0);
    CN39_sign_in(29) <= VN1619_sign_out(0);
    CN39_data_in(30) <= VN1657_data_out(0);
    CN39_sign_in(30) <= VN1657_sign_out(0);
    CN39_data_in(31) <= VN1736_data_out(0);
    CN39_sign_in(31) <= VN1736_sign_out(0);
    CN40_data_in(0) <= VN14_data_out(0);
    CN40_sign_in(0) <= VN14_sign_out(0);
    CN40_data_in(1) <= VN56_data_out(0);
    CN40_sign_in(1) <= VN56_sign_out(0);
    CN40_data_in(2) <= VN162_data_out(0);
    CN40_sign_in(2) <= VN162_sign_out(0);
    CN40_data_in(3) <= VN260_data_out(0);
    CN40_sign_in(3) <= VN260_sign_out(0);
    CN40_data_in(4) <= VN380_data_out(0);
    CN40_sign_in(4) <= VN380_sign_out(0);
    CN40_data_in(5) <= VN430_data_out(0);
    CN40_sign_in(5) <= VN430_sign_out(0);
    CN40_data_in(6) <= VN496_data_out(0);
    CN40_sign_in(6) <= VN496_sign_out(0);
    CN40_data_in(7) <= VN536_data_out(0);
    CN40_sign_in(7) <= VN536_sign_out(0);
    CN40_data_in(8) <= VN566_data_out(0);
    CN40_sign_in(8) <= VN566_sign_out(0);
    CN40_data_in(9) <= VN635_data_out(0);
    CN40_sign_in(9) <= VN635_sign_out(0);
    CN40_data_in(10) <= VN727_data_out(0);
    CN40_sign_in(10) <= VN727_sign_out(0);
    CN40_data_in(11) <= VN818_data_out(0);
    CN40_sign_in(11) <= VN818_sign_out(0);
    CN40_data_in(12) <= VN873_data_out(0);
    CN40_sign_in(12) <= VN873_sign_out(0);
    CN40_data_in(13) <= VN892_data_out(0);
    CN40_sign_in(13) <= VN892_sign_out(0);
    CN40_data_in(14) <= VN953_data_out(0);
    CN40_sign_in(14) <= VN953_sign_out(0);
    CN40_data_in(15) <= VN1044_data_out(0);
    CN40_sign_in(15) <= VN1044_sign_out(0);
    CN40_data_in(16) <= VN1160_data_out(0);
    CN40_sign_in(16) <= VN1160_sign_out(0);
    CN40_data_in(17) <= VN1242_data_out(0);
    CN40_sign_in(17) <= VN1242_sign_out(0);
    CN40_data_in(18) <= VN1279_data_out(0);
    CN40_sign_in(18) <= VN1279_sign_out(0);
    CN40_data_in(19) <= VN1353_data_out(0);
    CN40_sign_in(19) <= VN1353_sign_out(0);
    CN40_data_in(20) <= VN1409_data_out(0);
    CN40_sign_in(20) <= VN1409_sign_out(0);
    CN40_data_in(21) <= VN1569_data_out(0);
    CN40_sign_in(21) <= VN1569_sign_out(0);
    CN40_data_in(22) <= VN1601_data_out(0);
    CN40_sign_in(22) <= VN1601_sign_out(0);
    CN40_data_in(23) <= VN1618_data_out(0);
    CN40_sign_in(23) <= VN1618_sign_out(0);
    CN40_data_in(24) <= VN1656_data_out(0);
    CN40_sign_in(24) <= VN1656_sign_out(0);
    CN40_data_in(25) <= VN1717_data_out(0);
    CN40_sign_in(25) <= VN1717_sign_out(0);
    CN40_data_in(26) <= VN1856_data_out(0);
    CN40_sign_in(26) <= VN1856_sign_out(0);
    CN40_data_in(27) <= VN1912_data_out(0);
    CN40_sign_in(27) <= VN1912_sign_out(0);
    CN40_data_in(28) <= VN1974_data_out(0);
    CN40_sign_in(28) <= VN1974_sign_out(0);
    CN40_data_in(29) <= VN1984_data_out(0);
    CN40_sign_in(29) <= VN1984_sign_out(0);
    CN40_data_in(30) <= VN1991_data_out(0);
    CN40_sign_in(30) <= VN1991_sign_out(0);
    CN40_data_in(31) <= VN1992_data_out(0);
    CN40_sign_in(31) <= VN1992_sign_out(0);
    CN41_data_in(0) <= VN13_data_out(0);
    CN41_sign_in(0) <= VN13_sign_out(0);
    CN41_data_in(1) <= VN55_data_out(0);
    CN41_sign_in(1) <= VN55_sign_out(0);
    CN41_data_in(2) <= VN161_data_out(0);
    CN41_sign_in(2) <= VN161_sign_out(0);
    CN41_data_in(3) <= VN190_data_out(0);
    CN41_sign_in(3) <= VN190_sign_out(0);
    CN41_data_in(4) <= VN259_data_out(0);
    CN41_sign_in(4) <= VN259_sign_out(0);
    CN41_data_in(5) <= VN328_data_out(0);
    CN41_sign_in(5) <= VN328_sign_out(0);
    CN41_data_in(6) <= VN379_data_out(0);
    CN41_sign_in(6) <= VN379_sign_out(0);
    CN41_data_in(7) <= VN429_data_out(0);
    CN41_sign_in(7) <= VN429_sign_out(0);
    CN41_data_in(8) <= VN495_data_out(0);
    CN41_sign_in(8) <= VN495_sign_out(0);
    CN41_data_in(9) <= VN535_data_out(0);
    CN41_sign_in(9) <= VN535_sign_out(0);
    CN41_data_in(10) <= VN565_data_out(0);
    CN41_sign_in(10) <= VN565_sign_out(0);
    CN41_data_in(11) <= VN634_data_out(0);
    CN41_sign_in(11) <= VN634_sign_out(0);
    CN41_data_in(12) <= VN710_data_out(0);
    CN41_sign_in(12) <= VN710_sign_out(0);
    CN41_data_in(13) <= VN726_data_out(0);
    CN41_sign_in(13) <= VN726_sign_out(0);
    CN41_data_in(14) <= VN817_data_out(0);
    CN41_sign_in(14) <= VN817_sign_out(0);
    CN41_data_in(15) <= VN872_data_out(0);
    CN41_sign_in(15) <= VN872_sign_out(0);
    CN41_data_in(16) <= VN891_data_out(0);
    CN41_sign_in(16) <= VN891_sign_out(0);
    CN41_data_in(17) <= VN952_data_out(0);
    CN41_sign_in(17) <= VN952_sign_out(0);
    CN41_data_in(18) <= VN1043_data_out(0);
    CN41_sign_in(18) <= VN1043_sign_out(0);
    CN41_data_in(19) <= VN1094_data_out(0);
    CN41_sign_in(19) <= VN1094_sign_out(0);
    CN41_data_in(20) <= VN1159_data_out(0);
    CN41_sign_in(20) <= VN1159_sign_out(0);
    CN41_data_in(21) <= VN1278_data_out(0);
    CN41_sign_in(21) <= VN1278_sign_out(0);
    CN41_data_in(22) <= VN1309_data_out(0);
    CN41_sign_in(22) <= VN1309_sign_out(0);
    CN41_data_in(23) <= VN1352_data_out(0);
    CN41_sign_in(23) <= VN1352_sign_out(0);
    CN41_data_in(24) <= VN1408_data_out(0);
    CN41_sign_in(24) <= VN1408_sign_out(0);
    CN41_data_in(25) <= VN1568_data_out(0);
    CN41_sign_in(25) <= VN1568_sign_out(0);
    CN41_data_in(26) <= VN1600_data_out(0);
    CN41_sign_in(26) <= VN1600_sign_out(0);
    CN41_data_in(27) <= VN1617_data_out(0);
    CN41_sign_in(27) <= VN1617_sign_out(0);
    CN41_data_in(28) <= VN1716_data_out(0);
    CN41_sign_in(28) <= VN1716_sign_out(0);
    CN41_data_in(29) <= VN1748_data_out(0);
    CN41_sign_in(29) <= VN1748_sign_out(0);
    CN41_data_in(30) <= VN1755_data_out(0);
    CN41_sign_in(30) <= VN1755_sign_out(0);
    CN41_data_in(31) <= VN1816_data_out(0);
    CN41_sign_in(31) <= VN1816_sign_out(0);
    CN42_data_in(0) <= VN12_data_out(0);
    CN42_sign_in(0) <= VN12_sign_out(0);
    CN42_data_in(1) <= VN54_data_out(0);
    CN42_sign_in(1) <= VN54_sign_out(0);
    CN42_data_in(2) <= VN160_data_out(0);
    CN42_sign_in(2) <= VN160_sign_out(0);
    CN42_data_in(3) <= VN189_data_out(0);
    CN42_sign_in(3) <= VN189_sign_out(0);
    CN42_data_in(4) <= VN258_data_out(0);
    CN42_sign_in(4) <= VN258_sign_out(0);
    CN42_data_in(5) <= VN327_data_out(0);
    CN42_sign_in(5) <= VN327_sign_out(0);
    CN42_data_in(6) <= VN378_data_out(0);
    CN42_sign_in(6) <= VN378_sign_out(0);
    CN42_data_in(7) <= VN428_data_out(0);
    CN42_sign_in(7) <= VN428_sign_out(0);
    CN42_data_in(8) <= VN494_data_out(0);
    CN42_sign_in(8) <= VN494_sign_out(0);
    CN42_data_in(9) <= VN534_data_out(0);
    CN42_sign_in(9) <= VN534_sign_out(0);
    CN42_data_in(10) <= VN564_data_out(0);
    CN42_sign_in(10) <= VN564_sign_out(0);
    CN42_data_in(11) <= VN633_data_out(0);
    CN42_sign_in(11) <= VN633_sign_out(0);
    CN42_data_in(12) <= VN709_data_out(0);
    CN42_sign_in(12) <= VN709_sign_out(0);
    CN42_data_in(13) <= VN725_data_out(0);
    CN42_sign_in(13) <= VN725_sign_out(0);
    CN42_data_in(14) <= VN816_data_out(0);
    CN42_sign_in(14) <= VN816_sign_out(0);
    CN42_data_in(15) <= VN871_data_out(0);
    CN42_sign_in(15) <= VN871_sign_out(0);
    CN42_data_in(16) <= VN890_data_out(0);
    CN42_sign_in(16) <= VN890_sign_out(0);
    CN42_data_in(17) <= VN951_data_out(0);
    CN42_sign_in(17) <= VN951_sign_out(0);
    CN42_data_in(18) <= VN1042_data_out(0);
    CN42_sign_in(18) <= VN1042_sign_out(0);
    CN42_data_in(19) <= VN1093_data_out(0);
    CN42_sign_in(19) <= VN1093_sign_out(0);
    CN42_data_in(20) <= VN1158_data_out(0);
    CN42_sign_in(20) <= VN1158_sign_out(0);
    CN42_data_in(21) <= VN1241_data_out(0);
    CN42_sign_in(21) <= VN1241_sign_out(0);
    CN42_data_in(22) <= VN1308_data_out(0);
    CN42_sign_in(22) <= VN1308_sign_out(0);
    CN42_data_in(23) <= VN1351_data_out(0);
    CN42_sign_in(23) <= VN1351_sign_out(0);
    CN42_data_in(24) <= VN1407_data_out(0);
    CN42_sign_in(24) <= VN1407_sign_out(0);
    CN42_data_in(25) <= VN1516_data_out(0);
    CN42_sign_in(25) <= VN1516_sign_out(0);
    CN42_data_in(26) <= VN1553_data_out(0);
    CN42_sign_in(26) <= VN1553_sign_out(0);
    CN42_data_in(27) <= VN1567_data_out(0);
    CN42_sign_in(27) <= VN1567_sign_out(0);
    CN42_data_in(28) <= VN1616_data_out(0);
    CN42_sign_in(28) <= VN1616_sign_out(0);
    CN42_data_in(29) <= VN1655_data_out(0);
    CN42_sign_in(29) <= VN1655_sign_out(0);
    CN42_data_in(30) <= VN1715_data_out(0);
    CN42_sign_in(30) <= VN1715_sign_out(0);
    CN42_data_in(31) <= VN1737_data_out(0);
    CN42_sign_in(31) <= VN1737_sign_out(0);
    CN43_data_in(0) <= VN109_data_out(0);
    CN43_sign_in(0) <= VN109_sign_out(0);
    CN43_data_in(1) <= VN159_data_out(0);
    CN43_sign_in(1) <= VN159_sign_out(0);
    CN43_data_in(2) <= VN188_data_out(0);
    CN43_sign_in(2) <= VN188_sign_out(0);
    CN43_data_in(3) <= VN257_data_out(0);
    CN43_sign_in(3) <= VN257_sign_out(0);
    CN43_data_in(4) <= VN326_data_out(0);
    CN43_sign_in(4) <= VN326_sign_out(0);
    CN43_data_in(5) <= VN377_data_out(0);
    CN43_sign_in(5) <= VN377_sign_out(0);
    CN43_data_in(6) <= VN427_data_out(0);
    CN43_sign_in(6) <= VN427_sign_out(0);
    CN43_data_in(7) <= VN493_data_out(0);
    CN43_sign_in(7) <= VN493_sign_out(0);
    CN43_data_in(8) <= VN533_data_out(0);
    CN43_sign_in(8) <= VN533_sign_out(0);
    CN43_data_in(9) <= VN563_data_out(0);
    CN43_sign_in(9) <= VN563_sign_out(0);
    CN43_data_in(10) <= VN632_data_out(0);
    CN43_sign_in(10) <= VN632_sign_out(0);
    CN43_data_in(11) <= VN708_data_out(0);
    CN43_sign_in(11) <= VN708_sign_out(0);
    CN43_data_in(12) <= VN815_data_out(0);
    CN43_sign_in(12) <= VN815_sign_out(0);
    CN43_data_in(13) <= VN870_data_out(0);
    CN43_sign_in(13) <= VN870_sign_out(0);
    CN43_data_in(14) <= VN889_data_out(0);
    CN43_sign_in(14) <= VN889_sign_out(0);
    CN43_data_in(15) <= VN950_data_out(0);
    CN43_sign_in(15) <= VN950_sign_out(0);
    CN43_data_in(16) <= VN1041_data_out(0);
    CN43_sign_in(16) <= VN1041_sign_out(0);
    CN43_data_in(17) <= VN1092_data_out(0);
    CN43_sign_in(17) <= VN1092_sign_out(0);
    CN43_data_in(18) <= VN1157_data_out(0);
    CN43_sign_in(18) <= VN1157_sign_out(0);
    CN43_data_in(19) <= VN1277_data_out(0);
    CN43_sign_in(19) <= VN1277_sign_out(0);
    CN43_data_in(20) <= VN1307_data_out(0);
    CN43_sign_in(20) <= VN1307_sign_out(0);
    CN43_data_in(21) <= VN1350_data_out(0);
    CN43_sign_in(21) <= VN1350_sign_out(0);
    CN43_data_in(22) <= VN1406_data_out(0);
    CN43_sign_in(22) <= VN1406_sign_out(0);
    CN43_data_in(23) <= VN1515_data_out(0);
    CN43_sign_in(23) <= VN1515_sign_out(0);
    CN43_data_in(24) <= VN1566_data_out(0);
    CN43_sign_in(24) <= VN1566_sign_out(0);
    CN43_data_in(25) <= VN1599_data_out(0);
    CN43_sign_in(25) <= VN1599_sign_out(0);
    CN43_data_in(26) <= VN1615_data_out(0);
    CN43_sign_in(26) <= VN1615_sign_out(0);
    CN43_data_in(27) <= VN1654_data_out(0);
    CN43_sign_in(27) <= VN1654_sign_out(0);
    CN43_data_in(28) <= VN1749_data_out(0);
    CN43_sign_in(28) <= VN1749_sign_out(0);
    CN43_data_in(29) <= VN1762_data_out(0);
    CN43_sign_in(29) <= VN1762_sign_out(0);
    CN43_data_in(30) <= VN1889_data_out(0);
    CN43_sign_in(30) <= VN1889_sign_out(0);
    CN43_data_in(31) <= VN1906_data_out(0);
    CN43_sign_in(31) <= VN1906_sign_out(0);
    CN44_data_in(0) <= VN11_data_out(0);
    CN44_sign_in(0) <= VN11_sign_out(0);
    CN44_data_in(1) <= VN108_data_out(0);
    CN44_sign_in(1) <= VN108_sign_out(0);
    CN44_data_in(2) <= VN158_data_out(0);
    CN44_sign_in(2) <= VN158_sign_out(0);
    CN44_data_in(3) <= VN187_data_out(0);
    CN44_sign_in(3) <= VN187_sign_out(0);
    CN44_data_in(4) <= VN256_data_out(0);
    CN44_sign_in(4) <= VN256_sign_out(0);
    CN44_data_in(5) <= VN325_data_out(0);
    CN44_sign_in(5) <= VN325_sign_out(0);
    CN44_data_in(6) <= VN376_data_out(0);
    CN44_sign_in(6) <= VN376_sign_out(0);
    CN44_data_in(7) <= VN426_data_out(0);
    CN44_sign_in(7) <= VN426_sign_out(0);
    CN44_data_in(8) <= VN492_data_out(0);
    CN44_sign_in(8) <= VN492_sign_out(0);
    CN44_data_in(9) <= VN532_data_out(0);
    CN44_sign_in(9) <= VN532_sign_out(0);
    CN44_data_in(10) <= VN562_data_out(0);
    CN44_sign_in(10) <= VN562_sign_out(0);
    CN44_data_in(11) <= VN631_data_out(0);
    CN44_sign_in(11) <= VN631_sign_out(0);
    CN44_data_in(12) <= VN707_data_out(0);
    CN44_sign_in(12) <= VN707_sign_out(0);
    CN44_data_in(13) <= VN724_data_out(0);
    CN44_sign_in(13) <= VN724_sign_out(0);
    CN44_data_in(14) <= VN814_data_out(0);
    CN44_sign_in(14) <= VN814_sign_out(0);
    CN44_data_in(15) <= VN869_data_out(0);
    CN44_sign_in(15) <= VN869_sign_out(0);
    CN44_data_in(16) <= VN888_data_out(0);
    CN44_sign_in(16) <= VN888_sign_out(0);
    CN44_data_in(17) <= VN949_data_out(0);
    CN44_sign_in(17) <= VN949_sign_out(0);
    CN44_data_in(18) <= VN1040_data_out(0);
    CN44_sign_in(18) <= VN1040_sign_out(0);
    CN44_data_in(19) <= VN1091_data_out(0);
    CN44_sign_in(19) <= VN1091_sign_out(0);
    CN44_data_in(20) <= VN1156_data_out(0);
    CN44_sign_in(20) <= VN1156_sign_out(0);
    CN44_data_in(21) <= VN1217_data_out(0);
    CN44_sign_in(21) <= VN1217_sign_out(0);
    CN44_data_in(22) <= VN1240_data_out(0);
    CN44_sign_in(22) <= VN1240_sign_out(0);
    CN44_data_in(23) <= VN1276_data_out(0);
    CN44_sign_in(23) <= VN1276_sign_out(0);
    CN44_data_in(24) <= VN1306_data_out(0);
    CN44_sign_in(24) <= VN1306_sign_out(0);
    CN44_data_in(25) <= VN1349_data_out(0);
    CN44_sign_in(25) <= VN1349_sign_out(0);
    CN44_data_in(26) <= VN1405_data_out(0);
    CN44_sign_in(26) <= VN1405_sign_out(0);
    CN44_data_in(27) <= VN1565_data_out(0);
    CN44_sign_in(27) <= VN1565_sign_out(0);
    CN44_data_in(28) <= VN1598_data_out(0);
    CN44_sign_in(28) <= VN1598_sign_out(0);
    CN44_data_in(29) <= VN1614_data_out(0);
    CN44_sign_in(29) <= VN1614_sign_out(0);
    CN44_data_in(30) <= VN1714_data_out(0);
    CN44_sign_in(30) <= VN1714_sign_out(0);
    CN44_data_in(31) <= VN1738_data_out(0);
    CN44_sign_in(31) <= VN1738_sign_out(0);
    CN45_data_in(0) <= VN10_data_out(0);
    CN45_sign_in(0) <= VN10_sign_out(0);
    CN45_data_in(1) <= VN107_data_out(0);
    CN45_sign_in(1) <= VN107_sign_out(0);
    CN45_data_in(2) <= VN157_data_out(0);
    CN45_sign_in(2) <= VN157_sign_out(0);
    CN45_data_in(3) <= VN186_data_out(0);
    CN45_sign_in(3) <= VN186_sign_out(0);
    CN45_data_in(4) <= VN255_data_out(0);
    CN45_sign_in(4) <= VN255_sign_out(0);
    CN45_data_in(5) <= VN324_data_out(0);
    CN45_sign_in(5) <= VN324_sign_out(0);
    CN45_data_in(6) <= VN375_data_out(0);
    CN45_sign_in(6) <= VN375_sign_out(0);
    CN45_data_in(7) <= VN425_data_out(0);
    CN45_sign_in(7) <= VN425_sign_out(0);
    CN45_data_in(8) <= VN491_data_out(0);
    CN45_sign_in(8) <= VN491_sign_out(0);
    CN45_data_in(9) <= VN531_data_out(0);
    CN45_sign_in(9) <= VN531_sign_out(0);
    CN45_data_in(10) <= VN561_data_out(0);
    CN45_sign_in(10) <= VN561_sign_out(0);
    CN45_data_in(11) <= VN630_data_out(0);
    CN45_sign_in(11) <= VN630_sign_out(0);
    CN45_data_in(12) <= VN706_data_out(0);
    CN45_sign_in(12) <= VN706_sign_out(0);
    CN45_data_in(13) <= VN723_data_out(0);
    CN45_sign_in(13) <= VN723_sign_out(0);
    CN45_data_in(14) <= VN813_data_out(0);
    CN45_sign_in(14) <= VN813_sign_out(0);
    CN45_data_in(15) <= VN868_data_out(0);
    CN45_sign_in(15) <= VN868_sign_out(0);
    CN45_data_in(16) <= VN943_data_out(0);
    CN45_sign_in(16) <= VN943_sign_out(0);
    CN45_data_in(17) <= VN948_data_out(0);
    CN45_sign_in(17) <= VN948_sign_out(0);
    CN45_data_in(18) <= VN1039_data_out(0);
    CN45_sign_in(18) <= VN1039_sign_out(0);
    CN45_data_in(19) <= VN1090_data_out(0);
    CN45_sign_in(19) <= VN1090_sign_out(0);
    CN45_data_in(20) <= VN1155_data_out(0);
    CN45_sign_in(20) <= VN1155_sign_out(0);
    CN45_data_in(21) <= VN1216_data_out(0);
    CN45_sign_in(21) <= VN1216_sign_out(0);
    CN45_data_in(22) <= VN1224_data_out(0);
    CN45_sign_in(22) <= VN1224_sign_out(0);
    CN45_data_in(23) <= VN1305_data_out(0);
    CN45_sign_in(23) <= VN1305_sign_out(0);
    CN45_data_in(24) <= VN1348_data_out(0);
    CN45_sign_in(24) <= VN1348_sign_out(0);
    CN45_data_in(25) <= VN1404_data_out(0);
    CN45_sign_in(25) <= VN1404_sign_out(0);
    CN45_data_in(26) <= VN1564_data_out(0);
    CN45_sign_in(26) <= VN1564_sign_out(0);
    CN45_data_in(27) <= VN1597_data_out(0);
    CN45_sign_in(27) <= VN1597_sign_out(0);
    CN45_data_in(28) <= VN1653_data_out(0);
    CN45_sign_in(28) <= VN1653_sign_out(0);
    CN45_data_in(29) <= VN1713_data_out(0);
    CN45_sign_in(29) <= VN1713_sign_out(0);
    CN45_data_in(30) <= VN1756_data_out(0);
    CN45_sign_in(30) <= VN1756_sign_out(0);
    CN45_data_in(31) <= VN1817_data_out(0);
    CN45_sign_in(31) <= VN1817_sign_out(0);
    CN46_data_in(0) <= VN9_data_out(0);
    CN46_sign_in(0) <= VN9_sign_out(0);
    CN46_data_in(1) <= VN106_data_out(0);
    CN46_sign_in(1) <= VN106_sign_out(0);
    CN46_data_in(2) <= VN156_data_out(0);
    CN46_sign_in(2) <= VN156_sign_out(0);
    CN46_data_in(3) <= VN185_data_out(0);
    CN46_sign_in(3) <= VN185_sign_out(0);
    CN46_data_in(4) <= VN254_data_out(0);
    CN46_sign_in(4) <= VN254_sign_out(0);
    CN46_data_in(5) <= VN323_data_out(0);
    CN46_sign_in(5) <= VN323_sign_out(0);
    CN46_data_in(6) <= VN374_data_out(0);
    CN46_sign_in(6) <= VN374_sign_out(0);
    CN46_data_in(7) <= VN424_data_out(0);
    CN46_sign_in(7) <= VN424_sign_out(0);
    CN46_data_in(8) <= VN490_data_out(0);
    CN46_sign_in(8) <= VN490_sign_out(0);
    CN46_data_in(9) <= VN530_data_out(0);
    CN46_sign_in(9) <= VN530_sign_out(0);
    CN46_data_in(10) <= VN615_data_out(0);
    CN46_sign_in(10) <= VN615_sign_out(0);
    CN46_data_in(11) <= VN705_data_out(0);
    CN46_sign_in(11) <= VN705_sign_out(0);
    CN46_data_in(12) <= VN776_data_out(0);
    CN46_sign_in(12) <= VN776_sign_out(0);
    CN46_data_in(13) <= VN812_data_out(0);
    CN46_sign_in(13) <= VN812_sign_out(0);
    CN46_data_in(14) <= VN867_data_out(0);
    CN46_sign_in(14) <= VN867_sign_out(0);
    CN46_data_in(15) <= VN947_data_out(0);
    CN46_sign_in(15) <= VN947_sign_out(0);
    CN46_data_in(16) <= VN1038_data_out(0);
    CN46_sign_in(16) <= VN1038_sign_out(0);
    CN46_data_in(17) <= VN1154_data_out(0);
    CN46_sign_in(17) <= VN1154_sign_out(0);
    CN46_data_in(18) <= VN1215_data_out(0);
    CN46_sign_in(18) <= VN1215_sign_out(0);
    CN46_data_in(19) <= VN1223_data_out(0);
    CN46_sign_in(19) <= VN1223_sign_out(0);
    CN46_data_in(20) <= VN1239_data_out(0);
    CN46_sign_in(20) <= VN1239_sign_out(0);
    CN46_data_in(21) <= VN1304_data_out(0);
    CN46_sign_in(21) <= VN1304_sign_out(0);
    CN46_data_in(22) <= VN1347_data_out(0);
    CN46_sign_in(22) <= VN1347_sign_out(0);
    CN46_data_in(23) <= VN1403_data_out(0);
    CN46_sign_in(23) <= VN1403_sign_out(0);
    CN46_data_in(24) <= VN1563_data_out(0);
    CN46_sign_in(24) <= VN1563_sign_out(0);
    CN46_data_in(25) <= VN1596_data_out(0);
    CN46_sign_in(25) <= VN1596_sign_out(0);
    CN46_data_in(26) <= VN1613_data_out(0);
    CN46_sign_in(26) <= VN1613_sign_out(0);
    CN46_data_in(27) <= VN1791_data_out(0);
    CN46_sign_in(27) <= VN1791_sign_out(0);
    CN46_data_in(28) <= VN1825_data_out(0);
    CN46_sign_in(28) <= VN1825_sign_out(0);
    CN46_data_in(29) <= VN1832_data_out(0);
    CN46_sign_in(29) <= VN1832_sign_out(0);
    CN46_data_in(30) <= VN1861_data_out(0);
    CN46_sign_in(30) <= VN1861_sign_out(0);
    CN46_data_in(31) <= VN1879_data_out(0);
    CN46_sign_in(31) <= VN1879_sign_out(0);
    CN47_data_in(0) <= VN8_data_out(0);
    CN47_sign_in(0) <= VN8_sign_out(0);
    CN47_data_in(1) <= VN155_data_out(0);
    CN47_sign_in(1) <= VN155_sign_out(0);
    CN47_data_in(2) <= VN253_data_out(0);
    CN47_sign_in(2) <= VN253_sign_out(0);
    CN47_data_in(3) <= VN373_data_out(0);
    CN47_sign_in(3) <= VN373_sign_out(0);
    CN47_data_in(4) <= VN489_data_out(0);
    CN47_sign_in(4) <= VN489_sign_out(0);
    CN47_data_in(5) <= VN529_data_out(0);
    CN47_sign_in(5) <= VN529_sign_out(0);
    CN47_data_in(6) <= VN614_data_out(0);
    CN47_sign_in(6) <= VN614_sign_out(0);
    CN47_data_in(7) <= VN629_data_out(0);
    CN47_sign_in(7) <= VN629_sign_out(0);
    CN47_data_in(8) <= VN811_data_out(0);
    CN47_sign_in(8) <= VN811_sign_out(0);
    CN47_data_in(9) <= VN942_data_out(0);
    CN47_sign_in(9) <= VN942_sign_out(0);
    CN47_data_in(10) <= VN946_data_out(0);
    CN47_sign_in(10) <= VN946_sign_out(0);
    CN47_data_in(11) <= VN1037_data_out(0);
    CN47_sign_in(11) <= VN1037_sign_out(0);
    CN47_data_in(12) <= VN1222_data_out(0);
    CN47_sign_in(12) <= VN1222_sign_out(0);
    CN47_data_in(13) <= VN1238_data_out(0);
    CN47_sign_in(13) <= VN1238_sign_out(0);
    CN47_data_in(14) <= VN1346_data_out(0);
    CN47_sign_in(14) <= VN1346_sign_out(0);
    CN47_data_in(15) <= VN1402_data_out(0);
    CN47_sign_in(15) <= VN1402_sign_out(0);
    CN47_data_in(16) <= VN1612_data_out(0);
    CN47_sign_in(16) <= VN1612_sign_out(0);
    CN47_data_in(17) <= VN1652_data_out(0);
    CN47_sign_in(17) <= VN1652_sign_out(0);
    CN47_data_in(18) <= VN1741_data_out(0);
    CN47_sign_in(18) <= VN1741_sign_out(0);
    CN47_data_in(19) <= VN1746_data_out(0);
    CN47_sign_in(19) <= VN1746_sign_out(0);
    CN47_data_in(20) <= VN1893_data_out(0);
    CN47_sign_in(20) <= VN1893_sign_out(0);
    CN47_data_in(21) <= VN1896_data_out(0);
    CN47_sign_in(21) <= VN1896_sign_out(0);
    CN47_data_in(22) <= VN1899_data_out(0);
    CN47_sign_in(22) <= VN1899_sign_out(0);
    CN47_data_in(23) <= VN1923_data_out(0);
    CN47_sign_in(23) <= VN1923_sign_out(0);
    CN47_data_in(24) <= VN1956_data_out(0);
    CN47_sign_in(24) <= VN1956_sign_out(0);
    CN47_data_in(25) <= VN1968_data_out(0);
    CN47_sign_in(25) <= VN1968_sign_out(0);
    CN47_data_in(26) <= VN2001_data_out(0);
    CN47_sign_in(26) <= VN2001_sign_out(0);
    CN47_data_in(27) <= VN2020_data_out(0);
    CN47_sign_in(27) <= VN2020_sign_out(0);
    CN47_data_in(28) <= VN2021_data_out(0);
    CN47_sign_in(28) <= VN2021_sign_out(0);
    CN47_data_in(29) <= VN2033_data_out(0);
    CN47_sign_in(29) <= VN2033_sign_out(0);
    CN47_data_in(30) <= VN2044_data_out(0);
    CN47_sign_in(30) <= VN2044_sign_out(0);
    CN47_data_in(31) <= VN2045_data_out(0);
    CN47_sign_in(31) <= VN2045_sign_out(0);
    CN48_data_in(0) <= VN7_data_out(0);
    CN48_sign_in(0) <= VN7_sign_out(0);
    CN48_data_in(1) <= VN154_data_out(0);
    CN48_sign_in(1) <= VN154_sign_out(0);
    CN48_data_in(2) <= VN322_data_out(0);
    CN48_sign_in(2) <= VN322_sign_out(0);
    CN48_data_in(3) <= VN372_data_out(0);
    CN48_sign_in(3) <= VN372_sign_out(0);
    CN48_data_in(4) <= VN423_data_out(0);
    CN48_sign_in(4) <= VN423_sign_out(0);
    CN48_data_in(5) <= VN488_data_out(0);
    CN48_sign_in(5) <= VN488_sign_out(0);
    CN48_data_in(6) <= VN528_data_out(0);
    CN48_sign_in(6) <= VN528_sign_out(0);
    CN48_data_in(7) <= VN613_data_out(0);
    CN48_sign_in(7) <= VN613_sign_out(0);
    CN48_data_in(8) <= VN704_data_out(0);
    CN48_sign_in(8) <= VN704_sign_out(0);
    CN48_data_in(9) <= VN775_data_out(0);
    CN48_sign_in(9) <= VN775_sign_out(0);
    CN48_data_in(10) <= VN810_data_out(0);
    CN48_sign_in(10) <= VN810_sign_out(0);
    CN48_data_in(11) <= VN941_data_out(0);
    CN48_sign_in(11) <= VN941_sign_out(0);
    CN48_data_in(12) <= VN945_data_out(0);
    CN48_sign_in(12) <= VN945_sign_out(0);
    CN48_data_in(13) <= VN1036_data_out(0);
    CN48_sign_in(13) <= VN1036_sign_out(0);
    CN48_data_in(14) <= VN1089_data_out(0);
    CN48_sign_in(14) <= VN1089_sign_out(0);
    CN48_data_in(15) <= VN1153_data_out(0);
    CN48_sign_in(15) <= VN1153_sign_out(0);
    CN48_data_in(16) <= VN1221_data_out(0);
    CN48_sign_in(16) <= VN1221_sign_out(0);
    CN48_data_in(17) <= VN1237_data_out(0);
    CN48_sign_in(17) <= VN1237_sign_out(0);
    CN48_data_in(18) <= VN1345_data_out(0);
    CN48_sign_in(18) <= VN1345_sign_out(0);
    CN48_data_in(19) <= VN1401_data_out(0);
    CN48_sign_in(19) <= VN1401_sign_out(0);
    CN48_data_in(20) <= VN1562_data_out(0);
    CN48_sign_in(20) <= VN1562_sign_out(0);
    CN48_data_in(21) <= VN1595_data_out(0);
    CN48_sign_in(21) <= VN1595_sign_out(0);
    CN48_data_in(22) <= VN1763_data_out(0);
    CN48_sign_in(22) <= VN1763_sign_out(0);
    CN48_data_in(23) <= VN1796_data_out(0);
    CN48_sign_in(23) <= VN1796_sign_out(0);
    CN48_data_in(24) <= VN1823_data_out(0);
    CN48_sign_in(24) <= VN1823_sign_out(0);
    CN48_data_in(25) <= VN1887_data_out(0);
    CN48_sign_in(25) <= VN1887_sign_out(0);
    CN48_data_in(26) <= VN1911_data_out(0);
    CN48_sign_in(26) <= VN1911_sign_out(0);
    CN48_data_in(27) <= VN1938_data_out(0);
    CN48_sign_in(27) <= VN1938_sign_out(0);
    CN48_data_in(28) <= VN1954_data_out(0);
    CN48_sign_in(28) <= VN1954_sign_out(0);
    CN48_data_in(29) <= VN1979_data_out(0);
    CN48_sign_in(29) <= VN1979_sign_out(0);
    CN48_data_in(30) <= VN2004_data_out(0);
    CN48_sign_in(30) <= VN2004_sign_out(0);
    CN48_data_in(31) <= VN2005_data_out(0);
    CN48_sign_in(31) <= VN2005_sign_out(0);
    CN49_data_in(0) <= VN6_data_out(0);
    CN49_sign_in(0) <= VN6_sign_out(0);
    CN49_data_in(1) <= VN105_data_out(0);
    CN49_sign_in(1) <= VN105_sign_out(0);
    CN49_data_in(2) <= VN153_data_out(0);
    CN49_sign_in(2) <= VN153_sign_out(0);
    CN49_data_in(3) <= VN184_data_out(0);
    CN49_sign_in(3) <= VN184_sign_out(0);
    CN49_data_in(4) <= VN252_data_out(0);
    CN49_sign_in(4) <= VN252_sign_out(0);
    CN49_data_in(5) <= VN321_data_out(0);
    CN49_sign_in(5) <= VN321_sign_out(0);
    CN49_data_in(6) <= VN371_data_out(0);
    CN49_sign_in(6) <= VN371_sign_out(0);
    CN49_data_in(7) <= VN422_data_out(0);
    CN49_sign_in(7) <= VN422_sign_out(0);
    CN49_data_in(8) <= VN487_data_out(0);
    CN49_sign_in(8) <= VN487_sign_out(0);
    CN49_data_in(9) <= VN527_data_out(0);
    CN49_sign_in(9) <= VN527_sign_out(0);
    CN49_data_in(10) <= VN612_data_out(0);
    CN49_sign_in(10) <= VN612_sign_out(0);
    CN49_data_in(11) <= VN628_data_out(0);
    CN49_sign_in(11) <= VN628_sign_out(0);
    CN49_data_in(12) <= VN703_data_out(0);
    CN49_sign_in(12) <= VN703_sign_out(0);
    CN49_data_in(13) <= VN774_data_out(0);
    CN49_sign_in(13) <= VN774_sign_out(0);
    CN49_data_in(14) <= VN809_data_out(0);
    CN49_sign_in(14) <= VN809_sign_out(0);
    CN49_data_in(15) <= VN866_data_out(0);
    CN49_sign_in(15) <= VN866_sign_out(0);
    CN49_data_in(16) <= VN940_data_out(0);
    CN49_sign_in(16) <= VN940_sign_out(0);
    CN49_data_in(17) <= VN944_data_out(0);
    CN49_sign_in(17) <= VN944_sign_out(0);
    CN49_data_in(18) <= VN1035_data_out(0);
    CN49_sign_in(18) <= VN1035_sign_out(0);
    CN49_data_in(19) <= VN1088_data_out(0);
    CN49_sign_in(19) <= VN1088_sign_out(0);
    CN49_data_in(20) <= VN1152_data_out(0);
    CN49_sign_in(20) <= VN1152_sign_out(0);
    CN49_data_in(21) <= VN1214_data_out(0);
    CN49_sign_in(21) <= VN1214_sign_out(0);
    CN49_data_in(22) <= VN1220_data_out(0);
    CN49_sign_in(22) <= VN1220_sign_out(0);
    CN49_data_in(23) <= VN1236_data_out(0);
    CN49_sign_in(23) <= VN1236_sign_out(0);
    CN49_data_in(24) <= VN1303_data_out(0);
    CN49_sign_in(24) <= VN1303_sign_out(0);
    CN49_data_in(25) <= VN1344_data_out(0);
    CN49_sign_in(25) <= VN1344_sign_out(0);
    CN49_data_in(26) <= VN1400_data_out(0);
    CN49_sign_in(26) <= VN1400_sign_out(0);
    CN49_data_in(27) <= VN1561_data_out(0);
    CN49_sign_in(27) <= VN1561_sign_out(0);
    CN49_data_in(28) <= VN1594_data_out(0);
    CN49_sign_in(28) <= VN1594_sign_out(0);
    CN49_data_in(29) <= VN1611_data_out(0);
    CN49_sign_in(29) <= VN1611_sign_out(0);
    CN49_data_in(30) <= VN1651_data_out(0);
    CN49_sign_in(30) <= VN1651_sign_out(0);
    CN49_data_in(31) <= VN1739_data_out(0);
    CN49_sign_in(31) <= VN1739_sign_out(0);
    CN50_data_in(0) <= VN5_data_out(0);
    CN50_sign_in(0) <= VN5_sign_out(0);
    CN50_data_in(1) <= VN104_data_out(0);
    CN50_sign_in(1) <= VN104_sign_out(0);
    CN50_data_in(2) <= VN152_data_out(0);
    CN50_sign_in(2) <= VN152_sign_out(0);
    CN50_data_in(3) <= VN183_data_out(0);
    CN50_sign_in(3) <= VN183_sign_out(0);
    CN50_data_in(4) <= VN251_data_out(0);
    CN50_sign_in(4) <= VN251_sign_out(0);
    CN50_data_in(5) <= VN320_data_out(0);
    CN50_sign_in(5) <= VN320_sign_out(0);
    CN50_data_in(6) <= VN370_data_out(0);
    CN50_sign_in(6) <= VN370_sign_out(0);
    CN50_data_in(7) <= VN421_data_out(0);
    CN50_sign_in(7) <= VN421_sign_out(0);
    CN50_data_in(8) <= VN486_data_out(0);
    CN50_sign_in(8) <= VN486_sign_out(0);
    CN50_data_in(9) <= VN526_data_out(0);
    CN50_sign_in(9) <= VN526_sign_out(0);
    CN50_data_in(10) <= VN611_data_out(0);
    CN50_sign_in(10) <= VN611_sign_out(0);
    CN50_data_in(11) <= VN627_data_out(0);
    CN50_sign_in(11) <= VN627_sign_out(0);
    CN50_data_in(12) <= VN702_data_out(0);
    CN50_sign_in(12) <= VN702_sign_out(0);
    CN50_data_in(13) <= VN773_data_out(0);
    CN50_sign_in(13) <= VN773_sign_out(0);
    CN50_data_in(14) <= VN808_data_out(0);
    CN50_sign_in(14) <= VN808_sign_out(0);
    CN50_data_in(15) <= VN865_data_out(0);
    CN50_sign_in(15) <= VN865_sign_out(0);
    CN50_data_in(16) <= VN939_data_out(0);
    CN50_sign_in(16) <= VN939_sign_out(0);
    CN50_data_in(17) <= VN1002_data_out(0);
    CN50_sign_in(17) <= VN1002_sign_out(0);
    CN50_data_in(18) <= VN1034_data_out(0);
    CN50_sign_in(18) <= VN1034_sign_out(0);
    CN50_data_in(19) <= VN1151_data_out(0);
    CN50_sign_in(19) <= VN1151_sign_out(0);
    CN50_data_in(20) <= VN1213_data_out(0);
    CN50_sign_in(20) <= VN1213_sign_out(0);
    CN50_data_in(21) <= VN1219_data_out(0);
    CN50_sign_in(21) <= VN1219_sign_out(0);
    CN50_data_in(22) <= VN1235_data_out(0);
    CN50_sign_in(22) <= VN1235_sign_out(0);
    CN50_data_in(23) <= VN1302_data_out(0);
    CN50_sign_in(23) <= VN1302_sign_out(0);
    CN50_data_in(24) <= VN1343_data_out(0);
    CN50_sign_in(24) <= VN1343_sign_out(0);
    CN50_data_in(25) <= VN1399_data_out(0);
    CN50_sign_in(25) <= VN1399_sign_out(0);
    CN50_data_in(26) <= VN1560_data_out(0);
    CN50_sign_in(26) <= VN1560_sign_out(0);
    CN50_data_in(27) <= VN1593_data_out(0);
    CN50_sign_in(27) <= VN1593_sign_out(0);
    CN50_data_in(28) <= VN1610_data_out(0);
    CN50_sign_in(28) <= VN1610_sign_out(0);
    CN50_data_in(29) <= VN1712_data_out(0);
    CN50_sign_in(29) <= VN1712_sign_out(0);
    CN50_data_in(30) <= VN1777_data_out(0);
    CN50_sign_in(30) <= VN1777_sign_out(0);
    CN50_data_in(31) <= VN1818_data_out(0);
    CN50_sign_in(31) <= VN1818_sign_out(0);
    CN51_data_in(0) <= VN4_data_out(0);
    CN51_sign_in(0) <= VN4_sign_out(0);
    CN51_data_in(1) <= VN103_data_out(0);
    CN51_sign_in(1) <= VN103_sign_out(0);
    CN51_data_in(2) <= VN182_data_out(0);
    CN51_sign_in(2) <= VN182_sign_out(0);
    CN51_data_in(3) <= VN250_data_out(0);
    CN51_sign_in(3) <= VN250_sign_out(0);
    CN51_data_in(4) <= VN319_data_out(0);
    CN51_sign_in(4) <= VN319_sign_out(0);
    CN51_data_in(5) <= VN369_data_out(0);
    CN51_sign_in(5) <= VN369_sign_out(0);
    CN51_data_in(6) <= VN420_data_out(0);
    CN51_sign_in(6) <= VN420_sign_out(0);
    CN51_data_in(7) <= VN485_data_out(0);
    CN51_sign_in(7) <= VN485_sign_out(0);
    CN51_data_in(8) <= VN525_data_out(0);
    CN51_sign_in(8) <= VN525_sign_out(0);
    CN51_data_in(9) <= VN610_data_out(0);
    CN51_sign_in(9) <= VN610_sign_out(0);
    CN51_data_in(10) <= VN626_data_out(0);
    CN51_sign_in(10) <= VN626_sign_out(0);
    CN51_data_in(11) <= VN701_data_out(0);
    CN51_sign_in(11) <= VN701_sign_out(0);
    CN51_data_in(12) <= VN807_data_out(0);
    CN51_sign_in(12) <= VN807_sign_out(0);
    CN51_data_in(13) <= VN938_data_out(0);
    CN51_sign_in(13) <= VN938_sign_out(0);
    CN51_data_in(14) <= VN1001_data_out(0);
    CN51_sign_in(14) <= VN1001_sign_out(0);
    CN51_data_in(15) <= VN1087_data_out(0);
    CN51_sign_in(15) <= VN1087_sign_out(0);
    CN51_data_in(16) <= VN1150_data_out(0);
    CN51_sign_in(16) <= VN1150_sign_out(0);
    CN51_data_in(17) <= VN1218_data_out(0);
    CN51_sign_in(17) <= VN1218_sign_out(0);
    CN51_data_in(18) <= VN1342_data_out(0);
    CN51_sign_in(18) <= VN1342_sign_out(0);
    CN51_data_in(19) <= VN1398_data_out(0);
    CN51_sign_in(19) <= VN1398_sign_out(0);
    CN51_data_in(20) <= VN1457_data_out(0);
    CN51_sign_in(20) <= VN1457_sign_out(0);
    CN51_data_in(21) <= VN1592_data_out(0);
    CN51_sign_in(21) <= VN1592_sign_out(0);
    CN51_data_in(22) <= VN1609_data_out(0);
    CN51_sign_in(22) <= VN1609_sign_out(0);
    CN51_data_in(23) <= VN1834_data_out(0);
    CN51_sign_in(23) <= VN1834_sign_out(0);
    CN51_data_in(24) <= VN1835_data_out(0);
    CN51_sign_in(24) <= VN1835_sign_out(0);
    CN51_data_in(25) <= VN1864_data_out(0);
    CN51_sign_in(25) <= VN1864_sign_out(0);
    CN51_data_in(26) <= VN1866_data_out(0);
    CN51_sign_in(26) <= VN1866_sign_out(0);
    CN51_data_in(27) <= VN1868_data_out(0);
    CN51_sign_in(27) <= VN1868_sign_out(0);
    CN51_data_in(28) <= VN1926_data_out(0);
    CN51_sign_in(28) <= VN1926_sign_out(0);
    CN51_data_in(29) <= VN1939_data_out(0);
    CN51_sign_in(29) <= VN1939_sign_out(0);
    CN51_data_in(30) <= VN1998_data_out(0);
    CN51_sign_in(30) <= VN1998_sign_out(0);
    CN51_data_in(31) <= VN2000_data_out(0);
    CN51_sign_in(31) <= VN2000_sign_out(0);
    CN52_data_in(0) <= VN102_data_out(0);
    CN52_sign_in(0) <= VN102_sign_out(0);
    CN52_data_in(1) <= VN151_data_out(0);
    CN52_sign_in(1) <= VN151_sign_out(0);
    CN52_data_in(2) <= VN181_data_out(0);
    CN52_sign_in(2) <= VN181_sign_out(0);
    CN52_data_in(3) <= VN318_data_out(0);
    CN52_sign_in(3) <= VN318_sign_out(0);
    CN52_data_in(4) <= VN368_data_out(0);
    CN52_sign_in(4) <= VN368_sign_out(0);
    CN52_data_in(5) <= VN419_data_out(0);
    CN52_sign_in(5) <= VN419_sign_out(0);
    CN52_data_in(6) <= VN524_data_out(0);
    CN52_sign_in(6) <= VN524_sign_out(0);
    CN52_data_in(7) <= VN609_data_out(0);
    CN52_sign_in(7) <= VN609_sign_out(0);
    CN52_data_in(8) <= VN625_data_out(0);
    CN52_sign_in(8) <= VN625_sign_out(0);
    CN52_data_in(9) <= VN700_data_out(0);
    CN52_sign_in(9) <= VN700_sign_out(0);
    CN52_data_in(10) <= VN772_data_out(0);
    CN52_sign_in(10) <= VN772_sign_out(0);
    CN52_data_in(11) <= VN806_data_out(0);
    CN52_sign_in(11) <= VN806_sign_out(0);
    CN52_data_in(12) <= VN864_data_out(0);
    CN52_sign_in(12) <= VN864_sign_out(0);
    CN52_data_in(13) <= VN937_data_out(0);
    CN52_sign_in(13) <= VN937_sign_out(0);
    CN52_data_in(14) <= VN1000_data_out(0);
    CN52_sign_in(14) <= VN1000_sign_out(0);
    CN52_data_in(15) <= VN1033_data_out(0);
    CN52_sign_in(15) <= VN1033_sign_out(0);
    CN52_data_in(16) <= VN1086_data_out(0);
    CN52_sign_in(16) <= VN1086_sign_out(0);
    CN52_data_in(17) <= VN1149_data_out(0);
    CN52_sign_in(17) <= VN1149_sign_out(0);
    CN52_data_in(18) <= VN1169_data_out(0);
    CN52_sign_in(18) <= VN1169_sign_out(0);
    CN52_data_in(19) <= VN1212_data_out(0);
    CN52_sign_in(19) <= VN1212_sign_out(0);
    CN52_data_in(20) <= VN1234_data_out(0);
    CN52_sign_in(20) <= VN1234_sign_out(0);
    CN52_data_in(21) <= VN1301_data_out(0);
    CN52_sign_in(21) <= VN1301_sign_out(0);
    CN52_data_in(22) <= VN1341_data_out(0);
    CN52_sign_in(22) <= VN1341_sign_out(0);
    CN52_data_in(23) <= VN1397_data_out(0);
    CN52_sign_in(23) <= VN1397_sign_out(0);
    CN52_data_in(24) <= VN1559_data_out(0);
    CN52_sign_in(24) <= VN1559_sign_out(0);
    CN52_data_in(25) <= VN1711_data_out(0);
    CN52_sign_in(25) <= VN1711_sign_out(0);
    CN52_data_in(26) <= VN1872_data_out(0);
    CN52_sign_in(26) <= VN1872_sign_out(0);
    CN52_data_in(27) <= VN1908_data_out(0);
    CN52_sign_in(27) <= VN1908_sign_out(0);
    CN52_data_in(28) <= VN1916_data_out(0);
    CN52_sign_in(28) <= VN1916_sign_out(0);
    CN52_data_in(29) <= VN1945_data_out(0);
    CN52_sign_in(29) <= VN1945_sign_out(0);
    CN52_data_in(30) <= VN2024_data_out(0);
    CN52_sign_in(30) <= VN2024_sign_out(0);
    CN52_data_in(31) <= VN2026_data_out(0);
    CN52_sign_in(31) <= VN2026_sign_out(0);
    CN53_data_in(0) <= VN3_data_out(0);
    CN53_sign_in(0) <= VN3_sign_out(0);
    CN53_data_in(1) <= VN150_data_out(0);
    CN53_sign_in(1) <= VN150_sign_out(0);
    CN53_data_in(2) <= VN180_data_out(0);
    CN53_sign_in(2) <= VN180_sign_out(0);
    CN53_data_in(3) <= VN249_data_out(0);
    CN53_sign_in(3) <= VN249_sign_out(0);
    CN53_data_in(4) <= VN317_data_out(0);
    CN53_sign_in(4) <= VN317_sign_out(0);
    CN53_data_in(5) <= VN367_data_out(0);
    CN53_sign_in(5) <= VN367_sign_out(0);
    CN53_data_in(6) <= VN418_data_out(0);
    CN53_sign_in(6) <= VN418_sign_out(0);
    CN53_data_in(7) <= VN484_data_out(0);
    CN53_sign_in(7) <= VN484_sign_out(0);
    CN53_data_in(8) <= VN608_data_out(0);
    CN53_sign_in(8) <= VN608_sign_out(0);
    CN53_data_in(9) <= VN699_data_out(0);
    CN53_sign_in(9) <= VN699_sign_out(0);
    CN53_data_in(10) <= VN771_data_out(0);
    CN53_sign_in(10) <= VN771_sign_out(0);
    CN53_data_in(11) <= VN863_data_out(0);
    CN53_sign_in(11) <= VN863_sign_out(0);
    CN53_data_in(12) <= VN936_data_out(0);
    CN53_sign_in(12) <= VN936_sign_out(0);
    CN53_data_in(13) <= VN1032_data_out(0);
    CN53_sign_in(13) <= VN1032_sign_out(0);
    CN53_data_in(14) <= VN1085_data_out(0);
    CN53_sign_in(14) <= VN1085_sign_out(0);
    CN53_data_in(15) <= VN1148_data_out(0);
    CN53_sign_in(15) <= VN1148_sign_out(0);
    CN53_data_in(16) <= VN1168_data_out(0);
    CN53_sign_in(16) <= VN1168_sign_out(0);
    CN53_data_in(17) <= VN1211_data_out(0);
    CN53_sign_in(17) <= VN1211_sign_out(0);
    CN53_data_in(18) <= VN1233_data_out(0);
    CN53_sign_in(18) <= VN1233_sign_out(0);
    CN53_data_in(19) <= VN1340_data_out(0);
    CN53_sign_in(19) <= VN1340_sign_out(0);
    CN53_data_in(20) <= VN1396_data_out(0);
    CN53_sign_in(20) <= VN1396_sign_out(0);
    CN53_data_in(21) <= VN1456_data_out(0);
    CN53_sign_in(21) <= VN1456_sign_out(0);
    CN53_data_in(22) <= VN1650_data_out(0);
    CN53_sign_in(22) <= VN1650_sign_out(0);
    CN53_data_in(23) <= VN1776_data_out(0);
    CN53_sign_in(23) <= VN1776_sign_out(0);
    CN53_data_in(24) <= VN1836_data_out(0);
    CN53_sign_in(24) <= VN1836_sign_out(0);
    CN53_data_in(25) <= VN1905_data_out(0);
    CN53_sign_in(25) <= VN1905_sign_out(0);
    CN53_data_in(26) <= VN1917_data_out(0);
    CN53_sign_in(26) <= VN1917_sign_out(0);
    CN53_data_in(27) <= VN1930_data_out(0);
    CN53_sign_in(27) <= VN1930_sign_out(0);
    CN53_data_in(28) <= VN2025_data_out(0);
    CN53_sign_in(28) <= VN2025_sign_out(0);
    CN53_data_in(29) <= VN2031_data_out(0);
    CN53_sign_in(29) <= VN2031_sign_out(0);
    CN53_data_in(30) <= VN2046_data_out(0);
    CN53_sign_in(30) <= VN2046_sign_out(0);
    CN53_data_in(31) <= VN2047_data_out(0);
    CN53_sign_in(31) <= VN2047_sign_out(0);
    CN54_data_in(0) <= VN2_data_out(0);
    CN54_sign_in(0) <= VN2_sign_out(0);
    CN54_data_in(1) <= VN101_data_out(0);
    CN54_sign_in(1) <= VN101_sign_out(0);
    CN54_data_in(2) <= VN149_data_out(0);
    CN54_sign_in(2) <= VN149_sign_out(0);
    CN54_data_in(3) <= VN179_data_out(0);
    CN54_sign_in(3) <= VN179_sign_out(0);
    CN54_data_in(4) <= VN316_data_out(0);
    CN54_sign_in(4) <= VN316_sign_out(0);
    CN54_data_in(5) <= VN366_data_out(0);
    CN54_sign_in(5) <= VN366_sign_out(0);
    CN54_data_in(6) <= VN417_data_out(0);
    CN54_sign_in(6) <= VN417_sign_out(0);
    CN54_data_in(7) <= VN523_data_out(0);
    CN54_sign_in(7) <= VN523_sign_out(0);
    CN54_data_in(8) <= VN698_data_out(0);
    CN54_sign_in(8) <= VN698_sign_out(0);
    CN54_data_in(9) <= VN770_data_out(0);
    CN54_sign_in(9) <= VN770_sign_out(0);
    CN54_data_in(10) <= VN805_data_out(0);
    CN54_sign_in(10) <= VN805_sign_out(0);
    CN54_data_in(11) <= VN862_data_out(0);
    CN54_sign_in(11) <= VN862_sign_out(0);
    CN54_data_in(12) <= VN935_data_out(0);
    CN54_sign_in(12) <= VN935_sign_out(0);
    CN54_data_in(13) <= VN999_data_out(0);
    CN54_sign_in(13) <= VN999_sign_out(0);
    CN54_data_in(14) <= VN1031_data_out(0);
    CN54_sign_in(14) <= VN1031_sign_out(0);
    CN54_data_in(15) <= VN1084_data_out(0);
    CN54_sign_in(15) <= VN1084_sign_out(0);
    CN54_data_in(16) <= VN1147_data_out(0);
    CN54_sign_in(16) <= VN1147_sign_out(0);
    CN54_data_in(17) <= VN1210_data_out(0);
    CN54_sign_in(17) <= VN1210_sign_out(0);
    CN54_data_in(18) <= VN1232_data_out(0);
    CN54_sign_in(18) <= VN1232_sign_out(0);
    CN54_data_in(19) <= VN1300_data_out(0);
    CN54_sign_in(19) <= VN1300_sign_out(0);
    CN54_data_in(20) <= VN1339_data_out(0);
    CN54_sign_in(20) <= VN1339_sign_out(0);
    CN54_data_in(21) <= VN1475_data_out(0);
    CN54_sign_in(21) <= VN1475_sign_out(0);
    CN54_data_in(22) <= VN1608_data_out(0);
    CN54_sign_in(22) <= VN1608_sign_out(0);
    CN54_data_in(23) <= VN1649_data_out(0);
    CN54_sign_in(23) <= VN1649_sign_out(0);
    CN54_data_in(24) <= VN1752_data_out(0);
    CN54_sign_in(24) <= VN1752_sign_out(0);
    CN54_data_in(25) <= VN1785_data_out(0);
    CN54_sign_in(25) <= VN1785_sign_out(0);
    CN54_data_in(26) <= VN1797_data_out(0);
    CN54_sign_in(26) <= VN1797_sign_out(0);
    CN54_data_in(27) <= VN1840_data_out(0);
    CN54_sign_in(27) <= VN1840_sign_out(0);
    CN54_data_in(28) <= VN1847_data_out(0);
    CN54_sign_in(28) <= VN1847_sign_out(0);
    CN54_data_in(29) <= VN1890_data_out(0);
    CN54_sign_in(29) <= VN1890_sign_out(0);
    CN54_data_in(30) <= VN1931_data_out(0);
    CN54_sign_in(30) <= VN1931_sign_out(0);
    CN54_data_in(31) <= VN1936_data_out(0);
    CN54_sign_in(31) <= VN1936_sign_out(0);
    CN55_data_in(0) <= VN1_data_out(0);
    CN55_sign_in(0) <= VN1_sign_out(0);
    CN55_data_in(1) <= VN100_data_out(0);
    CN55_sign_in(1) <= VN100_sign_out(0);
    CN55_data_in(2) <= VN148_data_out(0);
    CN55_sign_in(2) <= VN148_sign_out(0);
    CN55_data_in(3) <= VN178_data_out(0);
    CN55_sign_in(3) <= VN178_sign_out(0);
    CN55_data_in(4) <= VN248_data_out(0);
    CN55_sign_in(4) <= VN248_sign_out(0);
    CN55_data_in(5) <= VN315_data_out(0);
    CN55_sign_in(5) <= VN315_sign_out(0);
    CN55_data_in(6) <= VN365_data_out(0);
    CN55_sign_in(6) <= VN365_sign_out(0);
    CN55_data_in(7) <= VN416_data_out(0);
    CN55_sign_in(7) <= VN416_sign_out(0);
    CN55_data_in(8) <= VN483_data_out(0);
    CN55_sign_in(8) <= VN483_sign_out(0);
    CN55_data_in(9) <= VN522_data_out(0);
    CN55_sign_in(9) <= VN522_sign_out(0);
    CN55_data_in(10) <= VN607_data_out(0);
    CN55_sign_in(10) <= VN607_sign_out(0);
    CN55_data_in(11) <= VN624_data_out(0);
    CN55_sign_in(11) <= VN624_sign_out(0);
    CN55_data_in(12) <= VN697_data_out(0);
    CN55_sign_in(12) <= VN697_sign_out(0);
    CN55_data_in(13) <= VN769_data_out(0);
    CN55_sign_in(13) <= VN769_sign_out(0);
    CN55_data_in(14) <= VN804_data_out(0);
    CN55_sign_in(14) <= VN804_sign_out(0);
    CN55_data_in(15) <= VN861_data_out(0);
    CN55_sign_in(15) <= VN861_sign_out(0);
    CN55_data_in(16) <= VN934_data_out(0);
    CN55_sign_in(16) <= VN934_sign_out(0);
    CN55_data_in(17) <= VN998_data_out(0);
    CN55_sign_in(17) <= VN998_sign_out(0);
    CN55_data_in(18) <= VN1030_data_out(0);
    CN55_sign_in(18) <= VN1030_sign_out(0);
    CN55_data_in(19) <= VN1083_data_out(0);
    CN55_sign_in(19) <= VN1083_sign_out(0);
    CN55_data_in(20) <= VN1146_data_out(0);
    CN55_sign_in(20) <= VN1146_sign_out(0);
    CN55_data_in(21) <= VN1167_data_out(0);
    CN55_sign_in(21) <= VN1167_sign_out(0);
    CN55_data_in(22) <= VN1209_data_out(0);
    CN55_sign_in(22) <= VN1209_sign_out(0);
    CN55_data_in(23) <= VN1231_data_out(0);
    CN55_sign_in(23) <= VN1231_sign_out(0);
    CN55_data_in(24) <= VN1299_data_out(0);
    CN55_sign_in(24) <= VN1299_sign_out(0);
    CN55_data_in(25) <= VN1338_data_out(0);
    CN55_sign_in(25) <= VN1338_sign_out(0);
    CN55_data_in(26) <= VN1395_data_out(0);
    CN55_sign_in(26) <= VN1395_sign_out(0);
    CN55_data_in(27) <= VN1474_data_out(0);
    CN55_sign_in(27) <= VN1474_sign_out(0);
    CN55_data_in(28) <= VN1494_data_out(0);
    CN55_sign_in(28) <= VN1494_sign_out(0);
    CN55_data_in(29) <= VN1591_data_out(0);
    CN55_sign_in(29) <= VN1591_sign_out(0);
    CN55_data_in(30) <= VN1710_data_out(0);
    CN55_sign_in(30) <= VN1710_sign_out(0);
    CN55_data_in(31) <= VN1740_data_out(0);
    CN55_sign_in(31) <= VN1740_sign_out(0);
    CN56_data_in(0) <= VN0_data_out(0);
    CN56_sign_in(0) <= VN0_sign_out(0);
    CN56_data_in(1) <= VN99_data_out(0);
    CN56_sign_in(1) <= VN99_sign_out(0);
    CN56_data_in(2) <= VN147_data_out(0);
    CN56_sign_in(2) <= VN147_sign_out(0);
    CN56_data_in(3) <= VN177_data_out(0);
    CN56_sign_in(3) <= VN177_sign_out(0);
    CN56_data_in(4) <= VN247_data_out(0);
    CN56_sign_in(4) <= VN247_sign_out(0);
    CN56_data_in(5) <= VN314_data_out(0);
    CN56_sign_in(5) <= VN314_sign_out(0);
    CN56_data_in(6) <= VN364_data_out(0);
    CN56_sign_in(6) <= VN364_sign_out(0);
    CN56_data_in(7) <= VN415_data_out(0);
    CN56_sign_in(7) <= VN415_sign_out(0);
    CN56_data_in(8) <= VN482_data_out(0);
    CN56_sign_in(8) <= VN482_sign_out(0);
    CN56_data_in(9) <= VN521_data_out(0);
    CN56_sign_in(9) <= VN521_sign_out(0);
    CN56_data_in(10) <= VN606_data_out(0);
    CN56_sign_in(10) <= VN606_sign_out(0);
    CN56_data_in(11) <= VN623_data_out(0);
    CN56_sign_in(11) <= VN623_sign_out(0);
    CN56_data_in(12) <= VN696_data_out(0);
    CN56_sign_in(12) <= VN696_sign_out(0);
    CN56_data_in(13) <= VN803_data_out(0);
    CN56_sign_in(13) <= VN803_sign_out(0);
    CN56_data_in(14) <= VN860_data_out(0);
    CN56_sign_in(14) <= VN860_sign_out(0);
    CN56_data_in(15) <= VN933_data_out(0);
    CN56_sign_in(15) <= VN933_sign_out(0);
    CN56_data_in(16) <= VN997_data_out(0);
    CN56_sign_in(16) <= VN997_sign_out(0);
    CN56_data_in(17) <= VN1029_data_out(0);
    CN56_sign_in(17) <= VN1029_sign_out(0);
    CN56_data_in(18) <= VN1082_data_out(0);
    CN56_sign_in(18) <= VN1082_sign_out(0);
    CN56_data_in(19) <= VN1145_data_out(0);
    CN56_sign_in(19) <= VN1145_sign_out(0);
    CN56_data_in(20) <= VN1166_data_out(0);
    CN56_sign_in(20) <= VN1166_sign_out(0);
    CN56_data_in(21) <= VN1208_data_out(0);
    CN56_sign_in(21) <= VN1208_sign_out(0);
    CN56_data_in(22) <= VN1230_data_out(0);
    CN56_sign_in(22) <= VN1230_sign_out(0);
    CN56_data_in(23) <= VN1298_data_out(0);
    CN56_sign_in(23) <= VN1298_sign_out(0);
    CN56_data_in(24) <= VN1394_data_out(0);
    CN56_sign_in(24) <= VN1394_sign_out(0);
    CN56_data_in(25) <= VN1473_data_out(0);
    CN56_sign_in(25) <= VN1473_sign_out(0);
    CN56_data_in(26) <= VN1493_data_out(0);
    CN56_sign_in(26) <= VN1493_sign_out(0);
    CN56_data_in(27) <= VN1495_data_out(0);
    CN56_sign_in(27) <= VN1495_sign_out(0);
    CN56_data_in(28) <= VN1709_data_out(0);
    CN56_sign_in(28) <= VN1709_sign_out(0);
    CN56_data_in(29) <= VN1745_data_out(0);
    CN56_sign_in(29) <= VN1745_sign_out(0);
    CN56_data_in(30) <= VN1789_data_out(0);
    CN56_sign_in(30) <= VN1789_sign_out(0);
    CN56_data_in(31) <= VN1819_data_out(0);
    CN56_sign_in(31) <= VN1819_sign_out(0);
    CN57_data_in(0) <= VN98_data_out(0);
    CN57_sign_in(0) <= VN98_sign_out(0);
    CN57_data_in(1) <= VN146_data_out(0);
    CN57_sign_in(1) <= VN146_sign_out(0);
    CN57_data_in(2) <= VN176_data_out(0);
    CN57_sign_in(2) <= VN176_sign_out(0);
    CN57_data_in(3) <= VN246_data_out(0);
    CN57_sign_in(3) <= VN246_sign_out(0);
    CN57_data_in(4) <= VN313_data_out(0);
    CN57_sign_in(4) <= VN313_sign_out(0);
    CN57_data_in(5) <= VN363_data_out(0);
    CN57_sign_in(5) <= VN363_sign_out(0);
    CN57_data_in(6) <= VN414_data_out(0);
    CN57_sign_in(6) <= VN414_sign_out(0);
    CN57_data_in(7) <= VN481_data_out(0);
    CN57_sign_in(7) <= VN481_sign_out(0);
    CN57_data_in(8) <= VN520_data_out(0);
    CN57_sign_in(8) <= VN520_sign_out(0);
    CN57_data_in(9) <= VN605_data_out(0);
    CN57_sign_in(9) <= VN605_sign_out(0);
    CN57_data_in(10) <= VN622_data_out(0);
    CN57_sign_in(10) <= VN622_sign_out(0);
    CN57_data_in(11) <= VN695_data_out(0);
    CN57_sign_in(11) <= VN695_sign_out(0);
    CN57_data_in(12) <= VN768_data_out(0);
    CN57_sign_in(12) <= VN768_sign_out(0);
    CN57_data_in(13) <= VN802_data_out(0);
    CN57_sign_in(13) <= VN802_sign_out(0);
    CN57_data_in(14) <= VN859_data_out(0);
    CN57_sign_in(14) <= VN859_sign_out(0);
    CN57_data_in(15) <= VN932_data_out(0);
    CN57_sign_in(15) <= VN932_sign_out(0);
    CN57_data_in(16) <= VN996_data_out(0);
    CN57_sign_in(16) <= VN996_sign_out(0);
    CN57_data_in(17) <= VN1081_data_out(0);
    CN57_sign_in(17) <= VN1081_sign_out(0);
    CN57_data_in(18) <= VN1144_data_out(0);
    CN57_sign_in(18) <= VN1144_sign_out(0);
    CN57_data_in(19) <= VN1165_data_out(0);
    CN57_sign_in(19) <= VN1165_sign_out(0);
    CN57_data_in(20) <= VN1207_data_out(0);
    CN57_sign_in(20) <= VN1207_sign_out(0);
    CN57_data_in(21) <= VN1229_data_out(0);
    CN57_sign_in(21) <= VN1229_sign_out(0);
    CN57_data_in(22) <= VN1297_data_out(0);
    CN57_sign_in(22) <= VN1297_sign_out(0);
    CN57_data_in(23) <= VN1337_data_out(0);
    CN57_sign_in(23) <= VN1337_sign_out(0);
    CN57_data_in(24) <= VN1472_data_out(0);
    CN57_sign_in(24) <= VN1472_sign_out(0);
    CN57_data_in(25) <= VN1485_data_out(0);
    CN57_sign_in(25) <= VN1485_sign_out(0);
    CN57_data_in(26) <= VN1590_data_out(0);
    CN57_sign_in(26) <= VN1590_sign_out(0);
    CN57_data_in(27) <= VN1686_data_out(0);
    CN57_sign_in(27) <= VN1686_sign_out(0);
    CN57_data_in(28) <= VN1723_data_out(0);
    CN57_sign_in(28) <= VN1723_sign_out(0);
    CN57_data_in(29) <= VN1798_data_out(0);
    CN57_sign_in(29) <= VN1798_sign_out(0);
    CN57_data_in(30) <= VN1804_data_out(0);
    CN57_sign_in(30) <= VN1804_sign_out(0);
    CN57_data_in(31) <= VN1820_data_out(0);
    CN57_sign_in(31) <= VN1820_sign_out(0);
    CN58_data_in(0) <= VN97_data_out(0);
    CN58_sign_in(0) <= VN97_sign_out(0);
    CN58_data_in(1) <= VN145_data_out(0);
    CN58_sign_in(1) <= VN145_sign_out(0);
    CN58_data_in(2) <= VN175_data_out(0);
    CN58_sign_in(2) <= VN175_sign_out(0);
    CN58_data_in(3) <= VN312_data_out(0);
    CN58_sign_in(3) <= VN312_sign_out(0);
    CN58_data_in(4) <= VN362_data_out(0);
    CN58_sign_in(4) <= VN362_sign_out(0);
    CN58_data_in(5) <= VN413_data_out(0);
    CN58_sign_in(5) <= VN413_sign_out(0);
    CN58_data_in(6) <= VN480_data_out(0);
    CN58_sign_in(6) <= VN480_sign_out(0);
    CN58_data_in(7) <= VN519_data_out(0);
    CN58_sign_in(7) <= VN519_sign_out(0);
    CN58_data_in(8) <= VN604_data_out(0);
    CN58_sign_in(8) <= VN604_sign_out(0);
    CN58_data_in(9) <= VN621_data_out(0);
    CN58_sign_in(9) <= VN621_sign_out(0);
    CN58_data_in(10) <= VN694_data_out(0);
    CN58_sign_in(10) <= VN694_sign_out(0);
    CN58_data_in(11) <= VN767_data_out(0);
    CN58_sign_in(11) <= VN767_sign_out(0);
    CN58_data_in(12) <= VN801_data_out(0);
    CN58_sign_in(12) <= VN801_sign_out(0);
    CN58_data_in(13) <= VN858_data_out(0);
    CN58_sign_in(13) <= VN858_sign_out(0);
    CN58_data_in(14) <= VN931_data_out(0);
    CN58_sign_in(14) <= VN931_sign_out(0);
    CN58_data_in(15) <= VN995_data_out(0);
    CN58_sign_in(15) <= VN995_sign_out(0);
    CN58_data_in(16) <= VN1028_data_out(0);
    CN58_sign_in(16) <= VN1028_sign_out(0);
    CN58_data_in(17) <= VN1080_data_out(0);
    CN58_sign_in(17) <= VN1080_sign_out(0);
    CN58_data_in(18) <= VN1143_data_out(0);
    CN58_sign_in(18) <= VN1143_sign_out(0);
    CN58_data_in(19) <= VN1164_data_out(0);
    CN58_sign_in(19) <= VN1164_sign_out(0);
    CN58_data_in(20) <= VN1206_data_out(0);
    CN58_sign_in(20) <= VN1206_sign_out(0);
    CN58_data_in(21) <= VN1228_data_out(0);
    CN58_sign_in(21) <= VN1228_sign_out(0);
    CN58_data_in(22) <= VN1336_data_out(0);
    CN58_sign_in(22) <= VN1336_sign_out(0);
    CN58_data_in(23) <= VN1393_data_out(0);
    CN58_sign_in(23) <= VN1393_sign_out(0);
    CN58_data_in(24) <= VN1471_data_out(0);
    CN58_sign_in(24) <= VN1471_sign_out(0);
    CN58_data_in(25) <= VN1589_data_out(0);
    CN58_sign_in(25) <= VN1589_sign_out(0);
    CN58_data_in(26) <= VN1685_data_out(0);
    CN58_sign_in(26) <= VN1685_sign_out(0);
    CN58_data_in(27) <= VN1838_data_out(0);
    CN58_sign_in(27) <= VN1838_sign_out(0);
    CN58_data_in(28) <= VN1851_data_out(0);
    CN58_sign_in(28) <= VN1851_sign_out(0);
    CN58_data_in(29) <= VN1870_data_out(0);
    CN58_sign_in(29) <= VN1870_sign_out(0);
    CN58_data_in(30) <= VN1928_data_out(0);
    CN58_sign_in(30) <= VN1928_sign_out(0);
    CN58_data_in(31) <= VN1929_data_out(0);
    CN58_sign_in(31) <= VN1929_sign_out(0);
    CN59_data_in(0) <= VN144_data_out(0);
    CN59_sign_in(0) <= VN144_sign_out(0);
    CN59_data_in(1) <= VN174_data_out(0);
    CN59_sign_in(1) <= VN174_sign_out(0);
    CN59_data_in(2) <= VN245_data_out(0);
    CN59_sign_in(2) <= VN245_sign_out(0);
    CN59_data_in(3) <= VN311_data_out(0);
    CN59_sign_in(3) <= VN311_sign_out(0);
    CN59_data_in(4) <= VN361_data_out(0);
    CN59_sign_in(4) <= VN361_sign_out(0);
    CN59_data_in(5) <= VN412_data_out(0);
    CN59_sign_in(5) <= VN412_sign_out(0);
    CN59_data_in(6) <= VN479_data_out(0);
    CN59_sign_in(6) <= VN479_sign_out(0);
    CN59_data_in(7) <= VN603_data_out(0);
    CN59_sign_in(7) <= VN603_sign_out(0);
    CN59_data_in(8) <= VN693_data_out(0);
    CN59_sign_in(8) <= VN693_sign_out(0);
    CN59_data_in(9) <= VN766_data_out(0);
    CN59_sign_in(9) <= VN766_sign_out(0);
    CN59_data_in(10) <= VN857_data_out(0);
    CN59_sign_in(10) <= VN857_sign_out(0);
    CN59_data_in(11) <= VN994_data_out(0);
    CN59_sign_in(11) <= VN994_sign_out(0);
    CN59_data_in(12) <= VN1027_data_out(0);
    CN59_sign_in(12) <= VN1027_sign_out(0);
    CN59_data_in(13) <= VN1113_data_out(0);
    CN59_sign_in(13) <= VN1113_sign_out(0);
    CN59_data_in(14) <= VN1142_data_out(0);
    CN59_sign_in(14) <= VN1142_sign_out(0);
    CN59_data_in(15) <= VN1205_data_out(0);
    CN59_sign_in(15) <= VN1205_sign_out(0);
    CN59_data_in(16) <= VN1227_data_out(0);
    CN59_sign_in(16) <= VN1227_sign_out(0);
    CN59_data_in(17) <= VN1296_data_out(0);
    CN59_sign_in(17) <= VN1296_sign_out(0);
    CN59_data_in(18) <= VN1470_data_out(0);
    CN59_sign_in(18) <= VN1470_sign_out(0);
    CN59_data_in(19) <= VN1484_data_out(0);
    CN59_sign_in(19) <= VN1484_sign_out(0);
    CN59_data_in(20) <= VN1722_data_out(0);
    CN59_sign_in(20) <= VN1722_sign_out(0);
    CN59_data_in(21) <= VN1751_data_out(0);
    CN59_sign_in(21) <= VN1751_sign_out(0);
    CN59_data_in(22) <= VN1757_data_out(0);
    CN59_sign_in(22) <= VN1757_sign_out(0);
    CN59_data_in(23) <= VN1774_data_out(0);
    CN59_sign_in(23) <= VN1774_sign_out(0);
    CN59_data_in(24) <= VN1794_data_out(0);
    CN59_sign_in(24) <= VN1794_sign_out(0);
    CN59_data_in(25) <= VN1874_data_out(0);
    CN59_sign_in(25) <= VN1874_sign_out(0);
    CN59_data_in(26) <= VN1920_data_out(0);
    CN59_sign_in(26) <= VN1920_sign_out(0);
    CN59_data_in(27) <= VN1927_data_out(0);
    CN59_sign_in(27) <= VN1927_sign_out(0);
    CN59_data_in(28) <= VN1983_data_out(0);
    CN59_sign_in(28) <= VN1983_sign_out(0);
    CN59_data_in(29) <= VN2012_data_out(0);
    CN59_sign_in(29) <= VN2012_sign_out(0);
    CN59_data_in(30) <= VN2015_data_out(0);
    CN59_sign_in(30) <= VN2015_sign_out(0);
    CN59_data_in(31) <= VN2017_data_out(0);
    CN59_sign_in(31) <= VN2017_sign_out(0);
    CN60_data_in(0) <= VN96_data_out(0);
    CN60_sign_in(0) <= VN96_sign_out(0);
    CN60_data_in(1) <= VN143_data_out(0);
    CN60_sign_in(1) <= VN143_sign_out(0);
    CN60_data_in(2) <= VN173_data_out(0);
    CN60_sign_in(2) <= VN173_sign_out(0);
    CN60_data_in(3) <= VN244_data_out(0);
    CN60_sign_in(3) <= VN244_sign_out(0);
    CN60_data_in(4) <= VN310_data_out(0);
    CN60_sign_in(4) <= VN310_sign_out(0);
    CN60_data_in(5) <= VN360_data_out(0);
    CN60_sign_in(5) <= VN360_sign_out(0);
    CN60_data_in(6) <= VN411_data_out(0);
    CN60_sign_in(6) <= VN411_sign_out(0);
    CN60_data_in(7) <= VN478_data_out(0);
    CN60_sign_in(7) <= VN478_sign_out(0);
    CN60_data_in(8) <= VN518_data_out(0);
    CN60_sign_in(8) <= VN518_sign_out(0);
    CN60_data_in(9) <= VN692_data_out(0);
    CN60_sign_in(9) <= VN692_sign_out(0);
    CN60_data_in(10) <= VN765_data_out(0);
    CN60_sign_in(10) <= VN765_sign_out(0);
    CN60_data_in(11) <= VN800_data_out(0);
    CN60_sign_in(11) <= VN800_sign_out(0);
    CN60_data_in(12) <= VN993_data_out(0);
    CN60_sign_in(12) <= VN993_sign_out(0);
    CN60_data_in(13) <= VN1026_data_out(0);
    CN60_sign_in(13) <= VN1026_sign_out(0);
    CN60_data_in(14) <= VN1112_data_out(0);
    CN60_sign_in(14) <= VN1112_sign_out(0);
    CN60_data_in(15) <= VN1141_data_out(0);
    CN60_sign_in(15) <= VN1141_sign_out(0);
    CN60_data_in(16) <= VN1204_data_out(0);
    CN60_sign_in(16) <= VN1204_sign_out(0);
    CN60_data_in(17) <= VN1226_data_out(0);
    CN60_sign_in(17) <= VN1226_sign_out(0);
    CN60_data_in(18) <= VN1295_data_out(0);
    CN60_sign_in(18) <= VN1295_sign_out(0);
    CN60_data_in(19) <= VN1469_data_out(0);
    CN60_sign_in(19) <= VN1469_sign_out(0);
    CN60_data_in(20) <= VN1492_data_out(0);
    CN60_sign_in(20) <= VN1492_sign_out(0);
    CN60_data_in(21) <= VN1588_data_out(0);
    CN60_sign_in(21) <= VN1588_sign_out(0);
    CN60_data_in(22) <= VN1684_data_out(0);
    CN60_sign_in(22) <= VN1684_sign_out(0);
    CN60_data_in(23) <= VN1721_data_out(0);
    CN60_sign_in(23) <= VN1721_sign_out(0);
    CN60_data_in(24) <= VN1744_data_out(0);
    CN60_sign_in(24) <= VN1744_sign_out(0);
    CN60_data_in(25) <= VN1768_data_out(0);
    CN60_sign_in(25) <= VN1768_sign_out(0);
    CN60_data_in(26) <= VN1846_data_out(0);
    CN60_sign_in(26) <= VN1846_sign_out(0);
    CN60_data_in(27) <= VN1853_data_out(0);
    CN60_sign_in(27) <= VN1853_sign_out(0);
    CN60_data_in(28) <= VN1871_data_out(0);
    CN60_sign_in(28) <= VN1871_sign_out(0);
    CN60_data_in(29) <= VN1883_data_out(0);
    CN60_sign_in(29) <= VN1883_sign_out(0);
    CN60_data_in(30) <= VN1966_data_out(0);
    CN60_sign_in(30) <= VN1966_sign_out(0);
    CN60_data_in(31) <= VN1972_data_out(0);
    CN60_sign_in(31) <= VN1972_sign_out(0);
    CN61_data_in(0) <= VN95_data_out(0);
    CN61_sign_in(0) <= VN95_sign_out(0);
    CN61_data_in(1) <= VN142_data_out(0);
    CN61_sign_in(1) <= VN142_sign_out(0);
    CN61_data_in(2) <= VN172_data_out(0);
    CN61_sign_in(2) <= VN172_sign_out(0);
    CN61_data_in(3) <= VN243_data_out(0);
    CN61_sign_in(3) <= VN243_sign_out(0);
    CN61_data_in(4) <= VN309_data_out(0);
    CN61_sign_in(4) <= VN309_sign_out(0);
    CN61_data_in(5) <= VN359_data_out(0);
    CN61_sign_in(5) <= VN359_sign_out(0);
    CN61_data_in(6) <= VN410_data_out(0);
    CN61_sign_in(6) <= VN410_sign_out(0);
    CN61_data_in(7) <= VN477_data_out(0);
    CN61_sign_in(7) <= VN477_sign_out(0);
    CN61_data_in(8) <= VN517_data_out(0);
    CN61_sign_in(8) <= VN517_sign_out(0);
    CN61_data_in(9) <= VN602_data_out(0);
    CN61_sign_in(9) <= VN602_sign_out(0);
    CN61_data_in(10) <= VN620_data_out(0);
    CN61_sign_in(10) <= VN620_sign_out(0);
    CN61_data_in(11) <= VN691_data_out(0);
    CN61_sign_in(11) <= VN691_sign_out(0);
    CN61_data_in(12) <= VN764_data_out(0);
    CN61_sign_in(12) <= VN764_sign_out(0);
    CN61_data_in(13) <= VN856_data_out(0);
    CN61_sign_in(13) <= VN856_sign_out(0);
    CN61_data_in(14) <= VN930_data_out(0);
    CN61_sign_in(14) <= VN930_sign_out(0);
    CN61_data_in(15) <= VN992_data_out(0);
    CN61_sign_in(15) <= VN992_sign_out(0);
    CN61_data_in(16) <= VN1025_data_out(0);
    CN61_sign_in(16) <= VN1025_sign_out(0);
    CN61_data_in(17) <= VN1079_data_out(0);
    CN61_sign_in(17) <= VN1079_sign_out(0);
    CN61_data_in(18) <= VN1110_data_out(0);
    CN61_sign_in(18) <= VN1110_sign_out(0);
    CN61_data_in(19) <= VN1140_data_out(0);
    CN61_sign_in(19) <= VN1140_sign_out(0);
    CN61_data_in(20) <= VN1203_data_out(0);
    CN61_sign_in(20) <= VN1203_sign_out(0);
    CN61_data_in(21) <= VN1225_data_out(0);
    CN61_sign_in(21) <= VN1225_sign_out(0);
    CN61_data_in(22) <= VN1294_data_out(0);
    CN61_sign_in(22) <= VN1294_sign_out(0);
    CN61_data_in(23) <= VN1335_data_out(0);
    CN61_sign_in(23) <= VN1335_sign_out(0);
    CN61_data_in(24) <= VN1392_data_out(0);
    CN61_sign_in(24) <= VN1392_sign_out(0);
    CN61_data_in(25) <= VN1468_data_out(0);
    CN61_sign_in(25) <= VN1468_sign_out(0);
    CN61_data_in(26) <= VN1491_data_out(0);
    CN61_sign_in(26) <= VN1491_sign_out(0);
    CN61_data_in(27) <= VN1683_data_out(0);
    CN61_sign_in(27) <= VN1683_sign_out(0);
    CN61_data_in(28) <= VN1719_data_out(0);
    CN61_sign_in(28) <= VN1719_sign_out(0);
    CN61_data_in(29) <= VN1799_data_out(0);
    CN61_sign_in(29) <= VN1799_sign_out(0);
    CN61_data_in(30) <= VN1805_data_out(0);
    CN61_sign_in(30) <= VN1805_sign_out(0);
    CN61_data_in(31) <= VN1821_data_out(0);
    CN61_sign_in(31) <= VN1821_sign_out(0);
    CN62_data_in(0) <= VN94_data_out(0);
    CN62_sign_in(0) <= VN94_sign_out(0);
    CN62_data_in(1) <= VN141_data_out(0);
    CN62_sign_in(1) <= VN141_sign_out(0);
    CN62_data_in(2) <= VN171_data_out(0);
    CN62_sign_in(2) <= VN171_sign_out(0);
    CN62_data_in(3) <= VN242_data_out(0);
    CN62_sign_in(3) <= VN242_sign_out(0);
    CN62_data_in(4) <= VN308_data_out(0);
    CN62_sign_in(4) <= VN308_sign_out(0);
    CN62_data_in(5) <= VN358_data_out(0);
    CN62_sign_in(5) <= VN358_sign_out(0);
    CN62_data_in(6) <= VN409_data_out(0);
    CN62_sign_in(6) <= VN409_sign_out(0);
    CN62_data_in(7) <= VN619_data_out(0);
    CN62_sign_in(7) <= VN619_sign_out(0);
    CN62_data_in(8) <= VN690_data_out(0);
    CN62_sign_in(8) <= VN690_sign_out(0);
    CN62_data_in(9) <= VN799_data_out(0);
    CN62_sign_in(9) <= VN799_sign_out(0);
    CN62_data_in(10) <= VN855_data_out(0);
    CN62_sign_in(10) <= VN855_sign_out(0);
    CN62_data_in(11) <= VN929_data_out(0);
    CN62_sign_in(11) <= VN929_sign_out(0);
    CN62_data_in(12) <= VN1078_data_out(0);
    CN62_sign_in(12) <= VN1078_sign_out(0);
    CN62_data_in(13) <= VN1108_data_out(0);
    CN62_sign_in(13) <= VN1108_sign_out(0);
    CN62_data_in(14) <= VN1139_data_out(0);
    CN62_sign_in(14) <= VN1139_sign_out(0);
    CN62_data_in(15) <= VN1202_data_out(0);
    CN62_sign_in(15) <= VN1202_sign_out(0);
    CN62_data_in(16) <= VN1293_data_out(0);
    CN62_sign_in(16) <= VN1293_sign_out(0);
    CN62_data_in(17) <= VN1391_data_out(0);
    CN62_sign_in(17) <= VN1391_sign_out(0);
    CN62_data_in(18) <= VN1467_data_out(0);
    CN62_sign_in(18) <= VN1467_sign_out(0);
    CN62_data_in(19) <= VN1490_data_out(0);
    CN62_sign_in(19) <= VN1490_sign_out(0);
    CN62_data_in(20) <= VN1524_data_out(0);
    CN62_sign_in(20) <= VN1524_sign_out(0);
    CN62_data_in(21) <= VN1587_data_out(0);
    CN62_sign_in(21) <= VN1587_sign_out(0);
    CN62_data_in(22) <= VN1682_data_out(0);
    CN62_sign_in(22) <= VN1682_sign_out(0);
    CN62_data_in(23) <= VN1720_data_out(0);
    CN62_sign_in(23) <= VN1720_sign_out(0);
    CN62_data_in(24) <= VN1775_data_out(0);
    CN62_sign_in(24) <= VN1775_sign_out(0);
    CN62_data_in(25) <= VN1779_data_out(0);
    CN62_sign_in(25) <= VN1779_sign_out(0);
    CN62_data_in(26) <= VN1827_data_out(0);
    CN62_sign_in(26) <= VN1827_sign_out(0);
    CN62_data_in(27) <= VN1863_data_out(0);
    CN62_sign_in(27) <= VN1863_sign_out(0);
    CN62_data_in(28) <= VN1880_data_out(0);
    CN62_sign_in(28) <= VN1880_sign_out(0);
    CN62_data_in(29) <= VN2010_data_out(0);
    CN62_sign_in(29) <= VN2010_sign_out(0);
    CN62_data_in(30) <= VN2016_data_out(0);
    CN62_sign_in(30) <= VN2016_sign_out(0);
    CN62_data_in(31) <= VN2018_data_out(0);
    CN62_sign_in(31) <= VN2018_sign_out(0);
    CN63_data_in(0) <= VN52_data_out(0);
    CN63_sign_in(0) <= VN52_sign_out(0);
    CN63_data_in(1) <= VN93_data_out(0);
    CN63_sign_in(1) <= VN93_sign_out(0);
    CN63_data_in(2) <= VN140_data_out(0);
    CN63_sign_in(2) <= VN140_sign_out(0);
    CN63_data_in(3) <= VN357_data_out(0);
    CN63_sign_in(3) <= VN357_sign_out(0);
    CN63_data_in(4) <= VN516_data_out(0);
    CN63_sign_in(4) <= VN516_sign_out(0);
    CN63_data_in(5) <= VN601_data_out(0);
    CN63_sign_in(5) <= VN601_sign_out(0);
    CN63_data_in(6) <= VN618_data_out(0);
    CN63_sign_in(6) <= VN618_sign_out(0);
    CN63_data_in(7) <= VN763_data_out(0);
    CN63_sign_in(7) <= VN763_sign_out(0);
    CN63_data_in(8) <= VN798_data_out(0);
    CN63_sign_in(8) <= VN798_sign_out(0);
    CN63_data_in(9) <= VN928_data_out(0);
    CN63_sign_in(9) <= VN928_sign_out(0);
    CN63_data_in(10) <= VN991_data_out(0);
    CN63_sign_in(10) <= VN991_sign_out(0);
    CN63_data_in(11) <= VN1024_data_out(0);
    CN63_sign_in(11) <= VN1024_sign_out(0);
    CN63_data_in(12) <= VN1060_data_out(0);
    CN63_sign_in(12) <= VN1060_sign_out(0);
    CN63_data_in(13) <= VN1201_data_out(0);
    CN63_sign_in(13) <= VN1201_sign_out(0);
    CN63_data_in(14) <= VN1489_data_out(0);
    CN63_sign_in(14) <= VN1489_sign_out(0);
    CN63_data_in(15) <= VN1523_data_out(0);
    CN63_sign_in(15) <= VN1523_sign_out(0);
    CN63_data_in(16) <= VN1551_data_out(0);
    CN63_sign_in(16) <= VN1551_sign_out(0);
    CN63_data_in(17) <= VN1586_data_out(0);
    CN63_sign_in(17) <= VN1586_sign_out(0);
    CN63_data_in(18) <= VN1708_data_out(0);
    CN63_sign_in(18) <= VN1708_sign_out(0);
    CN63_data_in(19) <= VN1761_data_out(0);
    CN63_sign_in(19) <= VN1761_sign_out(0);
    CN63_data_in(20) <= VN1783_data_out(0);
    CN63_sign_in(20) <= VN1783_sign_out(0);
    CN63_data_in(21) <= VN1855_data_out(0);
    CN63_sign_in(21) <= VN1855_sign_out(0);
    CN63_data_in(22) <= VN1865_data_out(0);
    CN63_sign_in(22) <= VN1865_sign_out(0);
    CN63_data_in(23) <= VN1949_data_out(0);
    CN63_sign_in(23) <= VN1949_sign_out(0);
    CN63_data_in(24) <= VN1963_data_out(0);
    CN63_sign_in(24) <= VN1963_sign_out(0);
    CN63_data_in(25) <= VN1967_data_out(0);
    CN63_sign_in(25) <= VN1967_sign_out(0);
    CN63_data_in(26) <= VN1970_data_out(0);
    CN63_sign_in(26) <= VN1970_sign_out(0);
    CN63_data_in(27) <= VN1975_data_out(0);
    CN63_sign_in(27) <= VN1975_sign_out(0);
    CN63_data_in(28) <= VN2011_data_out(0);
    CN63_sign_in(28) <= VN2011_sign_out(0);
    CN63_data_in(29) <= VN2039_data_out(0);
    CN63_sign_in(29) <= VN2039_sign_out(0);
    CN63_data_in(30) <= VN2040_data_out(0);
    CN63_sign_in(30) <= VN2040_sign_out(0);
    CN63_data_in(31) <= VN2043_data_out(0);
    CN63_sign_in(31) <= VN2043_sign_out(0);
    CN64_data_in(0) <= VN53_data_out(1);
    CN64_sign_in(0) <= VN53_sign_out(1);
    CN64_data_in(1) <= VN109_data_out(1);
    CN64_sign_in(1) <= VN109_sign_out(1);
    CN64_data_in(2) <= VN130_data_out(1);
    CN64_sign_in(2) <= VN130_sign_out(1);
    CN64_data_in(3) <= VN245_data_out(1);
    CN64_sign_in(3) <= VN245_sign_out(1);
    CN64_data_in(4) <= VN299_data_out(1);
    CN64_sign_in(4) <= VN299_sign_out(1);
    CN64_data_in(5) <= VN342_data_out(1);
    CN64_sign_in(5) <= VN342_sign_out(1);
    CN64_data_in(6) <= VN442_data_out(1);
    CN64_sign_in(6) <= VN442_sign_out(1);
    CN64_data_in(7) <= VN458_data_out(1);
    CN64_sign_in(7) <= VN458_sign_out(1);
    CN64_data_in(8) <= VN535_data_out(1);
    CN64_sign_in(8) <= VN535_sign_out(1);
    CN64_data_in(9) <= VN580_data_out(1);
    CN64_sign_in(9) <= VN580_sign_out(1);
    CN64_data_in(10) <= VN641_data_out(1);
    CN64_sign_in(10) <= VN641_sign_out(1);
    CN64_data_in(11) <= VN763_data_out(1);
    CN64_sign_in(11) <= VN763_sign_out(1);
    CN64_data_in(12) <= VN796_data_out(1);
    CN64_sign_in(12) <= VN796_sign_out(1);
    CN64_data_in(13) <= VN859_data_out(1);
    CN64_sign_in(13) <= VN859_sign_out(1);
    CN64_data_in(14) <= VN894_data_out(1);
    CN64_sign_in(14) <= VN894_sign_out(1);
    CN64_data_in(15) <= VN944_data_out(1);
    CN64_sign_in(15) <= VN944_sign_out(1);
    CN64_data_in(16) <= VN1038_data_out(1);
    CN64_sign_in(16) <= VN1038_sign_out(1);
    CN64_data_in(17) <= VN1074_data_out(1);
    CN64_sign_in(17) <= VN1074_sign_out(1);
    CN64_data_in(18) <= VN1158_data_out(1);
    CN64_sign_in(18) <= VN1158_sign_out(1);
    CN64_data_in(19) <= VN1171_data_out(1);
    CN64_sign_in(19) <= VN1171_sign_out(1);
    CN64_data_in(20) <= VN1245_data_out(1);
    CN64_sign_in(20) <= VN1245_sign_out(1);
    CN64_data_in(21) <= VN1287_data_out(1);
    CN64_sign_in(21) <= VN1287_sign_out(1);
    CN64_data_in(22) <= VN1346_data_out(1);
    CN64_sign_in(22) <= VN1346_sign_out(1);
    CN64_data_in(23) <= VN1416_data_out(1);
    CN64_sign_in(23) <= VN1416_sign_out(1);
    CN64_data_in(24) <= VN1574_data_out(1);
    CN64_sign_in(24) <= VN1574_sign_out(1);
    CN64_data_in(25) <= VN1582_data_out(1);
    CN64_sign_in(25) <= VN1582_sign_out(1);
    CN64_data_in(26) <= VN1664_data_out(1);
    CN64_sign_in(26) <= VN1664_sign_out(1);
    CN64_data_in(27) <= VN1740_data_out(1);
    CN64_sign_in(27) <= VN1740_sign_out(1);
    CN64_data_in(28) <= VN1902_data_out(1);
    CN64_sign_in(28) <= VN1902_sign_out(1);
    CN64_data_in(29) <= VN1960_data_out(1);
    CN64_sign_in(29) <= VN1960_sign_out(1);
    CN64_data_in(30) <= VN1992_data_out(1);
    CN64_sign_in(30) <= VN1992_sign_out(1);
    CN64_data_in(31) <= VN1994_data_out(1);
    CN64_sign_in(31) <= VN1994_sign_out(1);
    CN65_data_in(0) <= VN51_data_out(1);
    CN65_sign_in(0) <= VN51_sign_out(1);
    CN65_data_in(1) <= VN74_data_out(1);
    CN65_sign_in(1) <= VN74_sign_out(1);
    CN65_data_in(2) <= VN141_data_out(1);
    CN65_sign_in(2) <= VN141_sign_out(1);
    CN65_data_in(3) <= VN189_data_out(1);
    CN65_sign_in(3) <= VN189_sign_out(1);
    CN65_data_in(4) <= VN286_data_out(1);
    CN65_sign_in(4) <= VN286_sign_out(1);
    CN65_data_in(5) <= VN386_data_out(1);
    CN65_sign_in(5) <= VN386_sign_out(1);
    CN65_data_in(6) <= VN399_data_out(1);
    CN65_sign_in(6) <= VN399_sign_out(1);
    CN65_data_in(7) <= VN478_data_out(1);
    CN65_sign_in(7) <= VN478_sign_out(1);
    CN65_data_in(8) <= VN521_data_out(1);
    CN65_sign_in(8) <= VN521_sign_out(1);
    CN65_data_in(9) <= VN587_data_out(1);
    CN65_sign_in(9) <= VN587_sign_out(1);
    CN65_data_in(10) <= VN655_data_out(1);
    CN65_sign_in(10) <= VN655_sign_out(1);
    CN65_data_in(11) <= VN707_data_out(1);
    CN65_sign_in(11) <= VN707_sign_out(1);
    CN65_data_in(12) <= VN757_data_out(1);
    CN65_sign_in(12) <= VN757_sign_out(1);
    CN65_data_in(13) <= VN787_data_out(1);
    CN65_sign_in(13) <= VN787_sign_out(1);
    CN65_data_in(14) <= VN943_data_out(1);
    CN65_sign_in(14) <= VN943_sign_out(1);
    CN65_data_in(15) <= VN982_data_out(1);
    CN65_sign_in(15) <= VN982_sign_out(1);
    CN65_data_in(16) <= VN1015_data_out(1);
    CN65_sign_in(16) <= VN1015_sign_out(1);
    CN65_data_in(17) <= VN1100_data_out(1);
    CN65_sign_in(17) <= VN1100_sign_out(1);
    CN65_data_in(18) <= VN1190_data_out(1);
    CN65_sign_in(18) <= VN1190_sign_out(1);
    CN65_data_in(19) <= VN1231_data_out(1);
    CN65_sign_in(19) <= VN1231_sign_out(1);
    CN65_data_in(20) <= VN1360_data_out(1);
    CN65_sign_in(20) <= VN1360_sign_out(1);
    CN65_data_in(21) <= VN1402_data_out(1);
    CN65_sign_in(21) <= VN1402_sign_out(1);
    CN65_data_in(22) <= VN1466_data_out(1);
    CN65_sign_in(22) <= VN1466_sign_out(1);
    CN65_data_in(23) <= VN1557_data_out(1);
    CN65_sign_in(23) <= VN1557_sign_out(1);
    CN65_data_in(24) <= VN1621_data_out(1);
    CN65_sign_in(24) <= VN1621_sign_out(1);
    CN65_data_in(25) <= VN1669_data_out(1);
    CN65_sign_in(25) <= VN1669_sign_out(1);
    CN65_data_in(26) <= VN1718_data_out(1);
    CN65_sign_in(26) <= VN1718_sign_out(1);
    CN65_data_in(27) <= VN1787_data_out(1);
    CN65_sign_in(27) <= VN1787_sign_out(1);
    CN65_data_in(28) <= VN1851_data_out(1);
    CN65_sign_in(28) <= VN1851_sign_out(1);
    CN65_data_in(29) <= VN1855_data_out(1);
    CN65_sign_in(29) <= VN1855_sign_out(1);
    CN65_data_in(30) <= VN1978_data_out(1);
    CN65_sign_in(30) <= VN1978_sign_out(1);
    CN65_data_in(31) <= VN1980_data_out(1);
    CN65_sign_in(31) <= VN1980_sign_out(1);
    CN66_data_in(0) <= VN50_data_out(1);
    CN66_sign_in(0) <= VN50_sign_out(1);
    CN66_data_in(1) <= VN66_data_out(1);
    CN66_sign_in(1) <= VN66_sign_out(1);
    CN66_data_in(2) <= VN155_data_out(1);
    CN66_sign_in(2) <= VN155_sign_out(1);
    CN66_data_in(3) <= VN244_data_out(1);
    CN66_sign_in(3) <= VN244_sign_out(1);
    CN66_data_in(4) <= VN404_data_out(1);
    CN66_sign_in(4) <= VN404_sign_out(1);
    CN66_data_in(5) <= VN480_data_out(1);
    CN66_sign_in(5) <= VN480_sign_out(1);
    CN66_data_in(6) <= VN531_data_out(1);
    CN66_sign_in(6) <= VN531_sign_out(1);
    CN66_data_in(7) <= VN609_data_out(1);
    CN66_sign_in(7) <= VN609_sign_out(1);
    CN66_data_in(8) <= VN666_data_out(1);
    CN66_sign_in(8) <= VN666_sign_out(1);
    CN66_data_in(9) <= VN701_data_out(1);
    CN66_sign_in(9) <= VN701_sign_out(1);
    CN66_data_in(10) <= VN751_data_out(1);
    CN66_sign_in(10) <= VN751_sign_out(1);
    CN66_data_in(11) <= VN871_data_out(1);
    CN66_sign_in(11) <= VN871_sign_out(1);
    CN66_data_in(12) <= VN933_data_out(1);
    CN66_sign_in(12) <= VN933_sign_out(1);
    CN66_data_in(13) <= VN973_data_out(1);
    CN66_sign_in(13) <= VN973_sign_out(1);
    CN66_data_in(14) <= VN1045_data_out(1);
    CN66_sign_in(14) <= VN1045_sign_out(1);
    CN66_data_in(15) <= VN1065_data_out(1);
    CN66_sign_in(15) <= VN1065_sign_out(1);
    CN66_data_in(16) <= VN1144_data_out(1);
    CN66_sign_in(16) <= VN1144_sign_out(1);
    CN66_data_in(17) <= VN1174_data_out(1);
    CN66_sign_in(17) <= VN1174_sign_out(1);
    CN66_data_in(18) <= VN1265_data_out(1);
    CN66_sign_in(18) <= VN1265_sign_out(1);
    CN66_data_in(19) <= VN1322_data_out(1);
    CN66_sign_in(19) <= VN1322_sign_out(1);
    CN66_data_in(20) <= VN1391_data_out(1);
    CN66_sign_in(20) <= VN1391_sign_out(1);
    CN66_data_in(21) <= VN1606_data_out(1);
    CN66_sign_in(21) <= VN1606_sign_out(1);
    CN66_data_in(22) <= VN1675_data_out(1);
    CN66_sign_in(22) <= VN1675_sign_out(1);
    CN66_data_in(23) <= VN1705_data_out(1);
    CN66_sign_in(23) <= VN1705_sign_out(1);
    CN66_data_in(24) <= VN1854_data_out(1);
    CN66_sign_in(24) <= VN1854_sign_out(1);
    CN66_data_in(25) <= VN1860_data_out(1);
    CN66_sign_in(25) <= VN1860_sign_out(1);
    CN66_data_in(26) <= VN1875_data_out(1);
    CN66_sign_in(26) <= VN1875_sign_out(1);
    CN66_data_in(27) <= VN1930_data_out(1);
    CN66_sign_in(27) <= VN1930_sign_out(1);
    CN66_data_in(28) <= VN1940_data_out(1);
    CN66_sign_in(28) <= VN1940_sign_out(1);
    CN66_data_in(29) <= VN1995_data_out(1);
    CN66_sign_in(29) <= VN1995_sign_out(1);
    CN66_data_in(30) <= VN2011_data_out(1);
    CN66_sign_in(30) <= VN2011_sign_out(1);
    CN66_data_in(31) <= VN2019_data_out(1);
    CN66_sign_in(31) <= VN2019_sign_out(1);
    CN67_data_in(0) <= VN97_data_out(1);
    CN67_sign_in(0) <= VN97_sign_out(1);
    CN67_data_in(1) <= VN275_data_out(1);
    CN67_sign_in(1) <= VN275_sign_out(1);
    CN67_data_in(2) <= VN322_data_out(1);
    CN67_sign_in(2) <= VN322_sign_out(1);
    CN67_data_in(3) <= VN365_data_out(1);
    CN67_sign_in(3) <= VN365_sign_out(1);
    CN67_data_in(4) <= VN393_data_out(1);
    CN67_sign_in(4) <= VN393_sign_out(1);
    CN67_data_in(5) <= VN449_data_out(1);
    CN67_sign_in(5) <= VN449_sign_out(1);
    CN67_data_in(6) <= VN524_data_out(1);
    CN67_sign_in(6) <= VN524_sign_out(1);
    CN67_data_in(7) <= VN561_data_out(1);
    CN67_sign_in(7) <= VN561_sign_out(1);
    CN67_data_in(8) <= VN638_data_out(1);
    CN67_sign_in(8) <= VN638_sign_out(1);
    CN67_data_in(9) <= VN734_data_out(1);
    CN67_sign_in(9) <= VN734_sign_out(1);
    CN67_data_in(10) <= VN874_data_out(1);
    CN67_sign_in(10) <= VN874_sign_out(1);
    CN67_data_in(11) <= VN960_data_out(1);
    CN67_sign_in(11) <= VN960_sign_out(1);
    CN67_data_in(12) <= VN1003_data_out(1);
    CN67_sign_in(12) <= VN1003_sign_out(1);
    CN67_data_in(13) <= VN1042_data_out(1);
    CN67_sign_in(13) <= VN1042_sign_out(1);
    CN67_data_in(14) <= VN1069_data_out(1);
    CN67_sign_in(14) <= VN1069_sign_out(1);
    CN67_data_in(15) <= VN1154_data_out(1);
    CN67_sign_in(15) <= VN1154_sign_out(1);
    CN67_data_in(16) <= VN1248_data_out(1);
    CN67_sign_in(16) <= VN1248_sign_out(1);
    CN67_data_in(17) <= VN1313_data_out(1);
    CN67_sign_in(17) <= VN1313_sign_out(1);
    CN67_data_in(18) <= VN1353_data_out(1);
    CN67_sign_in(18) <= VN1353_sign_out(1);
    CN67_data_in(19) <= VN1405_data_out(1);
    CN67_sign_in(19) <= VN1405_sign_out(1);
    CN67_data_in(20) <= VN1483_data_out(1);
    CN67_sign_in(20) <= VN1483_sign_out(1);
    CN67_data_in(21) <= VN1500_data_out(1);
    CN67_sign_in(21) <= VN1500_sign_out(1);
    CN67_data_in(22) <= VN1561_data_out(1);
    CN67_sign_in(22) <= VN1561_sign_out(1);
    CN67_data_in(23) <= VN1702_data_out(1);
    CN67_sign_in(23) <= VN1702_sign_out(1);
    CN67_data_in(24) <= VN1811_data_out(1);
    CN67_sign_in(24) <= VN1811_sign_out(1);
    CN67_data_in(25) <= VN1812_data_out(1);
    CN67_sign_in(25) <= VN1812_sign_out(1);
    CN67_data_in(26) <= VN1833_data_out(1);
    CN67_sign_in(26) <= VN1833_sign_out(1);
    CN67_data_in(27) <= VN1849_data_out(1);
    CN67_sign_in(27) <= VN1849_sign_out(1);
    CN67_data_in(28) <= VN1900_data_out(1);
    CN67_sign_in(28) <= VN1900_sign_out(1);
    CN67_data_in(29) <= VN1926_data_out(1);
    CN67_sign_in(29) <= VN1926_sign_out(1);
    CN67_data_in(30) <= VN2014_data_out(1);
    CN67_sign_in(30) <= VN2014_sign_out(1);
    CN67_data_in(31) <= VN2020_data_out(1);
    CN67_sign_in(31) <= VN2020_sign_out(1);
    CN68_data_in(0) <= VN49_data_out(1);
    CN68_sign_in(0) <= VN49_sign_out(1);
    CN68_data_in(1) <= VN112_data_out(1);
    CN68_sign_in(1) <= VN112_sign_out(1);
    CN68_data_in(2) <= VN210_data_out(1);
    CN68_sign_in(2) <= VN210_sign_out(1);
    CN68_data_in(3) <= VN256_data_out(1);
    CN68_sign_in(3) <= VN256_sign_out(1);
    CN68_data_in(4) <= VN318_data_out(1);
    CN68_sign_in(4) <= VN318_sign_out(1);
    CN68_data_in(5) <= VN381_data_out(1);
    CN68_sign_in(5) <= VN381_sign_out(1);
    CN68_data_in(6) <= VN417_data_out(1);
    CN68_sign_in(6) <= VN417_sign_out(1);
    CN68_data_in(7) <= VN485_data_out(1);
    CN68_sign_in(7) <= VN485_sign_out(1);
    CN68_data_in(8) <= VN528_data_out(1);
    CN68_sign_in(8) <= VN528_sign_out(1);
    CN68_data_in(9) <= VN601_data_out(1);
    CN68_sign_in(9) <= VN601_sign_out(1);
    CN68_data_in(10) <= VN627_data_out(1);
    CN68_sign_in(10) <= VN627_sign_out(1);
    CN68_data_in(11) <= VN694_data_out(1);
    CN68_sign_in(11) <= VN694_sign_out(1);
    CN68_data_in(12) <= VN741_data_out(1);
    CN68_sign_in(12) <= VN741_sign_out(1);
    CN68_data_in(13) <= VN791_data_out(1);
    CN68_sign_in(13) <= VN791_sign_out(1);
    CN68_data_in(14) <= VN861_data_out(1);
    CN68_sign_in(14) <= VN861_sign_out(1);
    CN68_data_in(15) <= VN897_data_out(1);
    CN68_sign_in(15) <= VN897_sign_out(1);
    CN68_data_in(16) <= VN979_data_out(1);
    CN68_sign_in(16) <= VN979_sign_out(1);
    CN68_data_in(17) <= VN1148_data_out(1);
    CN68_sign_in(17) <= VN1148_sign_out(1);
    CN68_data_in(18) <= VN1195_data_out(1);
    CN68_sign_in(18) <= VN1195_sign_out(1);
    CN68_data_in(19) <= VN1260_data_out(1);
    CN68_sign_in(19) <= VN1260_sign_out(1);
    CN68_data_in(20) <= VN1350_data_out(1);
    CN68_sign_in(20) <= VN1350_sign_out(1);
    CN68_data_in(21) <= VN1424_data_out(1);
    CN68_sign_in(21) <= VN1424_sign_out(1);
    CN68_data_in(22) <= VN1442_data_out(1);
    CN68_sign_in(22) <= VN1442_sign_out(1);
    CN68_data_in(23) <= VN1485_data_out(1);
    CN68_sign_in(23) <= VN1485_sign_out(1);
    CN68_data_in(24) <= VN1504_data_out(1);
    CN68_sign_in(24) <= VN1504_sign_out(1);
    CN68_data_in(25) <= VN1509_data_out(1);
    CN68_sign_in(25) <= VN1509_sign_out(1);
    CN68_data_in(26) <= VN1529_data_out(1);
    CN68_sign_in(26) <= VN1529_sign_out(1);
    CN68_data_in(27) <= VN1556_data_out(1);
    CN68_sign_in(27) <= VN1556_sign_out(1);
    CN68_data_in(28) <= VN1578_data_out(1);
    CN68_sign_in(28) <= VN1578_sign_out(1);
    CN68_data_in(29) <= VN1676_data_out(1);
    CN68_sign_in(29) <= VN1676_sign_out(1);
    CN68_data_in(30) <= VN1690_data_out(1);
    CN68_sign_in(30) <= VN1690_sign_out(1);
    CN68_data_in(31) <= VN1741_data_out(1);
    CN68_sign_in(31) <= VN1741_sign_out(1);
    CN69_data_in(0) <= VN48_data_out(1);
    CN69_sign_in(0) <= VN48_sign_out(1);
    CN69_data_in(1) <= VN101_data_out(1);
    CN69_sign_in(1) <= VN101_sign_out(1);
    CN69_data_in(2) <= VN135_data_out(1);
    CN69_sign_in(2) <= VN135_sign_out(1);
    CN69_data_in(3) <= VN215_data_out(1);
    CN69_sign_in(3) <= VN215_sign_out(1);
    CN69_data_in(4) <= VN259_data_out(1);
    CN69_sign_in(4) <= VN259_sign_out(1);
    CN69_data_in(5) <= VN283_data_out(1);
    CN69_sign_in(5) <= VN283_sign_out(1);
    CN69_data_in(6) <= VN351_data_out(1);
    CN69_sign_in(6) <= VN351_sign_out(1);
    CN69_data_in(7) <= VN498_data_out(1);
    CN69_sign_in(7) <= VN498_sign_out(1);
    CN69_data_in(8) <= VN602_data_out(1);
    CN69_sign_in(8) <= VN602_sign_out(1);
    CN69_data_in(9) <= VN674_data_out(1);
    CN69_sign_in(9) <= VN674_sign_out(1);
    CN69_data_in(10) <= VN785_data_out(1);
    CN69_sign_in(10) <= VN785_sign_out(1);
    CN69_data_in(11) <= VN836_data_out(1);
    CN69_sign_in(11) <= VN836_sign_out(1);
    CN69_data_in(12) <= VN910_data_out(1);
    CN69_sign_in(12) <= VN910_sign_out(1);
    CN69_data_in(13) <= VN951_data_out(1);
    CN69_sign_in(13) <= VN951_sign_out(1);
    CN69_data_in(14) <= VN1051_data_out(1);
    CN69_sign_in(14) <= VN1051_sign_out(1);
    CN69_data_in(15) <= VN1152_data_out(1);
    CN69_sign_in(15) <= VN1152_sign_out(1);
    CN69_data_in(16) <= VN1272_data_out(1);
    CN69_sign_in(16) <= VN1272_sign_out(1);
    CN69_data_in(17) <= VN1282_data_out(1);
    CN69_sign_in(17) <= VN1282_sign_out(1);
    CN69_data_in(18) <= VN1364_data_out(1);
    CN69_sign_in(18) <= VN1364_sign_out(1);
    CN69_data_in(19) <= VN1517_data_out(1);
    CN69_sign_in(19) <= VN1517_sign_out(1);
    CN69_data_in(20) <= VN1540_data_out(1);
    CN69_sign_in(20) <= VN1540_sign_out(1);
    CN69_data_in(21) <= VN1563_data_out(1);
    CN69_sign_in(21) <= VN1563_sign_out(1);
    CN69_data_in(22) <= VN1607_data_out(1);
    CN69_sign_in(22) <= VN1607_sign_out(1);
    CN69_data_in(23) <= VN1759_data_out(1);
    CN69_sign_in(23) <= VN1759_sign_out(1);
    CN69_data_in(24) <= VN1773_data_out(1);
    CN69_sign_in(24) <= VN1773_sign_out(1);
    CN69_data_in(25) <= VN1779_data_out(1);
    CN69_sign_in(25) <= VN1779_sign_out(1);
    CN69_data_in(26) <= VN1839_data_out(1);
    CN69_sign_in(26) <= VN1839_sign_out(1);
    CN69_data_in(27) <= VN1948_data_out(1);
    CN69_sign_in(27) <= VN1948_sign_out(1);
    CN69_data_in(28) <= VN1951_data_out(1);
    CN69_sign_in(28) <= VN1951_sign_out(1);
    CN69_data_in(29) <= VN1982_data_out(1);
    CN69_sign_in(29) <= VN1982_sign_out(1);
    CN69_data_in(30) <= VN2015_data_out(1);
    CN69_sign_in(30) <= VN2015_sign_out(1);
    CN69_data_in(31) <= VN2021_data_out(1);
    CN69_sign_in(31) <= VN2021_sign_out(1);
    CN70_data_in(0) <= VN47_data_out(1);
    CN70_sign_in(0) <= VN47_sign_out(1);
    CN70_data_in(1) <= VN104_data_out(1);
    CN70_sign_in(1) <= VN104_sign_out(1);
    CN70_data_in(2) <= VN136_data_out(1);
    CN70_sign_in(2) <= VN136_sign_out(1);
    CN70_data_in(3) <= VN206_data_out(1);
    CN70_sign_in(3) <= VN206_sign_out(1);
    CN70_data_in(4) <= VN246_data_out(1);
    CN70_sign_in(4) <= VN246_sign_out(1);
    CN70_data_in(5) <= VN301_data_out(1);
    CN70_sign_in(5) <= VN301_sign_out(1);
    CN70_data_in(6) <= VN389_data_out(1);
    CN70_sign_in(6) <= VN389_sign_out(1);
    CN70_data_in(7) <= VN407_data_out(1);
    CN70_sign_in(7) <= VN407_sign_out(1);
    CN70_data_in(8) <= VN450_data_out(1);
    CN70_sign_in(8) <= VN450_sign_out(1);
    CN70_data_in(9) <= VN556_data_out(1);
    CN70_sign_in(9) <= VN556_sign_out(1);
    CN70_data_in(10) <= VN572_data_out(1);
    CN70_sign_in(10) <= VN572_sign_out(1);
    CN70_data_in(11) <= VN629_data_out(1);
    CN70_sign_in(11) <= VN629_sign_out(1);
    CN70_data_in(12) <= VN713_data_out(1);
    CN70_sign_in(12) <= VN713_sign_out(1);
    CN70_data_in(13) <= VN762_data_out(1);
    CN70_sign_in(13) <= VN762_sign_out(1);
    CN70_data_in(14) <= VN822_data_out(1);
    CN70_sign_in(14) <= VN822_sign_out(1);
    CN70_data_in(15) <= VN857_data_out(1);
    CN70_sign_in(15) <= VN857_sign_out(1);
    CN70_data_in(16) <= VN921_data_out(1);
    CN70_sign_in(16) <= VN921_sign_out(1);
    CN70_data_in(17) <= VN948_data_out(1);
    CN70_sign_in(17) <= VN948_sign_out(1);
    CN70_data_in(18) <= VN1025_data_out(1);
    CN70_sign_in(18) <= VN1025_sign_out(1);
    CN70_data_in(19) <= VN1063_data_out(1);
    CN70_sign_in(19) <= VN1063_sign_out(1);
    CN70_data_in(20) <= VN1141_data_out(1);
    CN70_sign_in(20) <= VN1141_sign_out(1);
    CN70_data_in(21) <= VN1212_data_out(1);
    CN70_sign_in(21) <= VN1212_sign_out(1);
    CN70_data_in(22) <= VN1242_data_out(1);
    CN70_sign_in(22) <= VN1242_sign_out(1);
    CN70_data_in(23) <= VN1388_data_out(1);
    CN70_sign_in(23) <= VN1388_sign_out(1);
    CN70_data_in(24) <= VN1448_data_out(1);
    CN70_sign_in(24) <= VN1448_sign_out(1);
    CN70_data_in(25) <= VN1495_data_out(1);
    CN70_sign_in(25) <= VN1495_sign_out(1);
    CN70_data_in(26) <= VN1532_data_out(1);
    CN70_sign_in(26) <= VN1532_sign_out(1);
    CN70_data_in(27) <= VN1577_data_out(1);
    CN70_sign_in(27) <= VN1577_sign_out(1);
    CN70_data_in(28) <= VN1614_data_out(1);
    CN70_sign_in(28) <= VN1614_sign_out(1);
    CN70_data_in(29) <= VN1708_data_out(1);
    CN70_sign_in(29) <= VN1708_sign_out(1);
    CN70_data_in(30) <= VN1786_data_out(1);
    CN70_sign_in(30) <= VN1786_sign_out(1);
    CN70_data_in(31) <= VN1822_data_out(1);
    CN70_sign_in(31) <= VN1822_sign_out(1);
    CN71_data_in(0) <= VN46_data_out(1);
    CN71_sign_in(0) <= VN46_sign_out(1);
    CN71_data_in(1) <= VN95_data_out(1);
    CN71_sign_in(1) <= VN95_sign_out(1);
    CN71_data_in(2) <= VN176_data_out(1);
    CN71_sign_in(2) <= VN176_sign_out(1);
    CN71_data_in(3) <= VN276_data_out(1);
    CN71_sign_in(3) <= VN276_sign_out(1);
    CN71_data_in(4) <= VN302_data_out(1);
    CN71_sign_in(4) <= VN302_sign_out(1);
    CN71_data_in(5) <= VN353_data_out(1);
    CN71_sign_in(5) <= VN353_sign_out(1);
    CN71_data_in(6) <= VN479_data_out(1);
    CN71_sign_in(6) <= VN479_sign_out(1);
    CN71_data_in(7) <= VN538_data_out(1);
    CN71_sign_in(7) <= VN538_sign_out(1);
    CN71_data_in(8) <= VN650_data_out(1);
    CN71_sign_in(8) <= VN650_sign_out(1);
    CN71_data_in(9) <= VN739_data_out(1);
    CN71_sign_in(9) <= VN739_sign_out(1);
    CN71_data_in(10) <= VN828_data_out(1);
    CN71_sign_in(10) <= VN828_sign_out(1);
    CN71_data_in(11) <= VN883_data_out(1);
    CN71_sign_in(11) <= VN883_sign_out(1);
    CN71_data_in(12) <= VN891_data_out(1);
    CN71_sign_in(12) <= VN891_sign_out(1);
    CN71_data_in(13) <= VN964_data_out(1);
    CN71_sign_in(13) <= VN964_sign_out(1);
    CN71_data_in(14) <= VN1034_data_out(1);
    CN71_sign_in(14) <= VN1034_sign_out(1);
    CN71_data_in(15) <= VN1121_data_out(1);
    CN71_sign_in(15) <= VN1121_sign_out(1);
    CN71_data_in(16) <= VN1198_data_out(1);
    CN71_sign_in(16) <= VN1198_sign_out(1);
    CN71_data_in(17) <= VN1233_data_out(1);
    CN71_sign_in(17) <= VN1233_sign_out(1);
    CN71_data_in(18) <= VN1284_data_out(1);
    CN71_sign_in(18) <= VN1284_sign_out(1);
    CN71_data_in(19) <= VN1431_data_out(1);
    CN71_sign_in(19) <= VN1431_sign_out(1);
    CN71_data_in(20) <= VN1452_data_out(1);
    CN71_sign_in(20) <= VN1452_sign_out(1);
    CN71_data_in(21) <= VN1481_data_out(1);
    CN71_sign_in(21) <= VN1481_sign_out(1);
    CN71_data_in(22) <= VN1541_data_out(1);
    CN71_sign_in(22) <= VN1541_sign_out(1);
    CN71_data_in(23) <= VN1651_data_out(1);
    CN71_sign_in(23) <= VN1651_sign_out(1);
    CN71_data_in(24) <= VN1707_data_out(1);
    CN71_sign_in(24) <= VN1707_sign_out(1);
    CN71_data_in(25) <= VN1813_data_out(1);
    CN71_sign_in(25) <= VN1813_sign_out(1);
    CN71_data_in(26) <= VN1847_data_out(1);
    CN71_sign_in(26) <= VN1847_sign_out(1);
    CN71_data_in(27) <= VN1937_data_out(1);
    CN71_sign_in(27) <= VN1937_sign_out(1);
    CN71_data_in(28) <= VN1952_data_out(1);
    CN71_sign_in(28) <= VN1952_sign_out(1);
    CN71_data_in(29) <= VN2018_data_out(1);
    CN71_sign_in(29) <= VN2018_sign_out(1);
    CN71_data_in(30) <= VN2030_data_out(1);
    CN71_sign_in(30) <= VN2030_sign_out(1);
    CN71_data_in(31) <= VN2039_data_out(1);
    CN71_sign_in(31) <= VN2039_sign_out(1);
    CN72_data_in(0) <= VN45_data_out(1);
    CN72_sign_in(0) <= VN45_sign_out(1);
    CN72_data_in(1) <= VN75_data_out(1);
    CN72_sign_in(1) <= VN75_sign_out(1);
    CN72_data_in(2) <= VN162_data_out(1);
    CN72_sign_in(2) <= VN162_sign_out(1);
    CN72_data_in(3) <= VN183_data_out(1);
    CN72_sign_in(3) <= VN183_sign_out(1);
    CN72_data_in(4) <= VN243_data_out(1);
    CN72_sign_in(4) <= VN243_sign_out(1);
    CN72_data_in(5) <= VN367_data_out(1);
    CN72_sign_in(5) <= VN367_sign_out(1);
    CN72_data_in(6) <= VN435_data_out(1);
    CN72_sign_in(6) <= VN435_sign_out(1);
    CN72_data_in(7) <= VN493_data_out(1);
    CN72_sign_in(7) <= VN493_sign_out(1);
    CN72_data_in(8) <= VN552_data_out(1);
    CN72_sign_in(8) <= VN552_sign_out(1);
    CN72_data_in(9) <= VN565_data_out(1);
    CN72_sign_in(9) <= VN565_sign_out(1);
    CN72_data_in(10) <= VN657_data_out(1);
    CN72_sign_in(10) <= VN657_sign_out(1);
    CN72_data_in(11) <= VN680_data_out(1);
    CN72_sign_in(11) <= VN680_sign_out(1);
    CN72_data_in(12) <= VN775_data_out(1);
    CN72_sign_in(12) <= VN775_sign_out(1);
    CN72_data_in(13) <= VN867_data_out(1);
    CN72_sign_in(13) <= VN867_sign_out(1);
    CN72_data_in(14) <= VN935_data_out(1);
    CN72_sign_in(14) <= VN935_sign_out(1);
    CN72_data_in(15) <= VN957_data_out(1);
    CN72_sign_in(15) <= VN957_sign_out(1);
    CN72_data_in(16) <= VN1104_data_out(1);
    CN72_sign_in(16) <= VN1104_sign_out(1);
    CN72_data_in(17) <= VN1161_data_out(1);
    CN72_sign_in(17) <= VN1161_sign_out(1);
    CN72_data_in(18) <= VN1214_data_out(1);
    CN72_sign_in(18) <= VN1214_sign_out(1);
    CN72_data_in(19) <= VN1275_data_out(1);
    CN72_sign_in(19) <= VN1275_sign_out(1);
    CN72_data_in(20) <= VN1342_data_out(1);
    CN72_sign_in(20) <= VN1342_sign_out(1);
    CN72_data_in(21) <= VN1423_data_out(1);
    CN72_sign_in(21) <= VN1423_sign_out(1);
    CN72_data_in(22) <= VN1527_data_out(1);
    CN72_sign_in(22) <= VN1527_sign_out(1);
    CN72_data_in(23) <= VN1603_data_out(1);
    CN72_sign_in(23) <= VN1603_sign_out(1);
    CN72_data_in(24) <= VN1629_data_out(1);
    CN72_sign_in(24) <= VN1629_sign_out(1);
    CN72_data_in(25) <= VN1679_data_out(1);
    CN72_sign_in(25) <= VN1679_sign_out(1);
    CN72_data_in(26) <= VN1724_data_out(1);
    CN72_sign_in(26) <= VN1724_sign_out(1);
    CN72_data_in(27) <= VN1820_data_out(1);
    CN72_sign_in(27) <= VN1820_sign_out(1);
    CN72_data_in(28) <= VN1848_data_out(1);
    CN72_sign_in(28) <= VN1848_sign_out(1);
    CN72_data_in(29) <= VN1986_data_out(1);
    CN72_sign_in(29) <= VN1986_sign_out(1);
    CN72_data_in(30) <= VN2003_data_out(1);
    CN72_sign_in(30) <= VN2003_sign_out(1);
    CN72_data_in(31) <= VN2008_data_out(1);
    CN72_sign_in(31) <= VN2008_sign_out(1);
    CN73_data_in(0) <= VN44_data_out(1);
    CN73_sign_in(0) <= VN44_sign_out(1);
    CN73_data_in(1) <= VN56_data_out(1);
    CN73_sign_in(1) <= VN56_sign_out(1);
    CN73_data_in(2) <= VN121_data_out(1);
    CN73_sign_in(2) <= VN121_sign_out(1);
    CN73_data_in(3) <= VN219_data_out(1);
    CN73_sign_in(3) <= VN219_sign_out(1);
    CN73_data_in(4) <= VN328_data_out(1);
    CN73_sign_in(4) <= VN328_sign_out(1);
    CN73_data_in(5) <= VN363_data_out(1);
    CN73_sign_in(5) <= VN363_sign_out(1);
    CN73_data_in(6) <= VN415_data_out(1);
    CN73_sign_in(6) <= VN415_sign_out(1);
    CN73_data_in(7) <= VN507_data_out(1);
    CN73_sign_in(7) <= VN507_sign_out(1);
    CN73_data_in(8) <= VN573_data_out(1);
    CN73_sign_in(8) <= VN573_sign_out(1);
    CN73_data_in(9) <= VN708_data_out(1);
    CN73_sign_in(9) <= VN708_sign_out(1);
    CN73_data_in(10) <= VN723_data_out(1);
    CN73_sign_in(10) <= VN723_sign_out(1);
    CN73_data_in(11) <= VN795_data_out(1);
    CN73_sign_in(11) <= VN795_sign_out(1);
    CN73_data_in(12) <= VN838_data_out(1);
    CN73_sign_in(12) <= VN838_sign_out(1);
    CN73_data_in(13) <= VN923_data_out(1);
    CN73_sign_in(13) <= VN923_sign_out(1);
    CN73_data_in(14) <= VN990_data_out(1);
    CN73_sign_in(14) <= VN990_sign_out(1);
    CN73_data_in(15) <= VN1032_data_out(1);
    CN73_sign_in(15) <= VN1032_sign_out(1);
    CN73_data_in(16) <= VN1075_data_out(1);
    CN73_sign_in(16) <= VN1075_sign_out(1);
    CN73_data_in(17) <= VN1116_data_out(1);
    CN73_sign_in(17) <= VN1116_sign_out(1);
    CN73_data_in(18) <= VN1178_data_out(1);
    CN73_sign_in(18) <= VN1178_sign_out(1);
    CN73_data_in(19) <= VN1235_data_out(1);
    CN73_sign_in(19) <= VN1235_sign_out(1);
    CN73_data_in(20) <= VN1311_data_out(1);
    CN73_sign_in(20) <= VN1311_sign_out(1);
    CN73_data_in(21) <= VN1336_data_out(1);
    CN73_sign_in(21) <= VN1336_sign_out(1);
    CN73_data_in(22) <= VN1432_data_out(1);
    CN73_sign_in(22) <= VN1432_sign_out(1);
    CN73_data_in(23) <= VN1451_data_out(1);
    CN73_sign_in(23) <= VN1451_sign_out(1);
    CN73_data_in(24) <= VN1462_data_out(1);
    CN73_sign_in(24) <= VN1462_sign_out(1);
    CN73_data_in(25) <= VN1619_data_out(1);
    CN73_sign_in(25) <= VN1619_sign_out(1);
    CN73_data_in(26) <= VN1739_data_out(1);
    CN73_sign_in(26) <= VN1739_sign_out(1);
    CN73_data_in(27) <= VN1837_data_out(1);
    CN73_sign_in(27) <= VN1837_sign_out(1);
    CN73_data_in(28) <= VN1857_data_out(1);
    CN73_sign_in(28) <= VN1857_sign_out(1);
    CN73_data_in(29) <= VN1914_data_out(1);
    CN73_sign_in(29) <= VN1914_sign_out(1);
    CN73_data_in(30) <= VN1920_data_out(1);
    CN73_sign_in(30) <= VN1920_sign_out(1);
    CN73_data_in(31) <= VN1921_data_out(1);
    CN73_sign_in(31) <= VN1921_sign_out(1);
    CN74_data_in(0) <= VN43_data_out(1);
    CN74_sign_in(0) <= VN43_sign_out(1);
    CN74_data_in(1) <= VN70_data_out(1);
    CN74_sign_in(1) <= VN70_sign_out(1);
    CN74_data_in(2) <= VN125_data_out(1);
    CN74_sign_in(2) <= VN125_sign_out(1);
    CN74_data_in(3) <= VN221_data_out(1);
    CN74_sign_in(3) <= VN221_sign_out(1);
    CN74_data_in(4) <= VN290_data_out(1);
    CN74_sign_in(4) <= VN290_sign_out(1);
    CN74_data_in(5) <= VN384_data_out(1);
    CN74_sign_in(5) <= VN384_sign_out(1);
    CN74_data_in(6) <= VN427_data_out(1);
    CN74_sign_in(6) <= VN427_sign_out(1);
    CN74_data_in(7) <= VN501_data_out(1);
    CN74_sign_in(7) <= VN501_sign_out(1);
    CN74_data_in(8) <= VN532_data_out(1);
    CN74_sign_in(8) <= VN532_sign_out(1);
    CN74_data_in(9) <= VN658_data_out(1);
    CN74_sign_in(9) <= VN658_sign_out(1);
    CN74_data_in(10) <= VN696_data_out(1);
    CN74_sign_in(10) <= VN696_sign_out(1);
    CN74_data_in(11) <= VN764_data_out(1);
    CN74_sign_in(11) <= VN764_sign_out(1);
    CN74_data_in(12) <= VN885_data_out(1);
    CN74_sign_in(12) <= VN885_sign_out(1);
    CN74_data_in(13) <= VN938_data_out(1);
    CN74_sign_in(13) <= VN938_sign_out(1);
    CN74_data_in(14) <= VN1023_data_out(1);
    CN74_sign_in(14) <= VN1023_sign_out(1);
    CN74_data_in(15) <= VN1073_data_out(1);
    CN74_sign_in(15) <= VN1073_sign_out(1);
    CN74_data_in(16) <= VN1127_data_out(1);
    CN74_sign_in(16) <= VN1127_sign_out(1);
    CN74_data_in(17) <= VN1187_data_out(1);
    CN74_sign_in(17) <= VN1187_sign_out(1);
    CN74_data_in(18) <= VN1254_data_out(1);
    CN74_sign_in(18) <= VN1254_sign_out(1);
    CN74_data_in(19) <= VN1318_data_out(1);
    CN74_sign_in(19) <= VN1318_sign_out(1);
    CN74_data_in(20) <= VN1339_data_out(1);
    CN74_sign_in(20) <= VN1339_sign_out(1);
    CN74_data_in(21) <= VN1387_data_out(1);
    CN74_sign_in(21) <= VN1387_sign_out(1);
    CN74_data_in(22) <= VN1397_data_out(1);
    CN74_sign_in(22) <= VN1397_sign_out(1);
    CN74_data_in(23) <= VN1446_data_out(1);
    CN74_sign_in(23) <= VN1446_sign_out(1);
    CN74_data_in(24) <= VN1583_data_out(1);
    CN74_sign_in(24) <= VN1583_sign_out(1);
    CN74_data_in(25) <= VN1634_data_out(1);
    CN74_sign_in(25) <= VN1634_sign_out(1);
    CN74_data_in(26) <= VN1658_data_out(1);
    CN74_sign_in(26) <= VN1658_sign_out(1);
    CN74_data_in(27) <= VN1758_data_out(1);
    CN74_sign_in(27) <= VN1758_sign_out(1);
    CN74_data_in(28) <= VN1791_data_out(1);
    CN74_sign_in(28) <= VN1791_sign_out(1);
    CN74_data_in(29) <= VN1796_data_out(1);
    CN74_sign_in(29) <= VN1796_sign_out(1);
    CN74_data_in(30) <= VN1836_data_out(1);
    CN74_sign_in(30) <= VN1836_sign_out(1);
    CN74_data_in(31) <= VN1880_data_out(1);
    CN74_sign_in(31) <= VN1880_sign_out(1);
    CN75_data_in(0) <= VN42_data_out(1);
    CN75_sign_in(0) <= VN42_sign_out(1);
    CN75_data_in(1) <= VN81_data_out(1);
    CN75_sign_in(1) <= VN81_sign_out(1);
    CN75_data_in(2) <= VN170_data_out(1);
    CN75_sign_in(2) <= VN170_sign_out(1);
    CN75_data_in(3) <= VN192_data_out(1);
    CN75_sign_in(3) <= VN192_sign_out(1);
    CN75_data_in(4) <= VN278_data_out(1);
    CN75_sign_in(4) <= VN278_sign_out(1);
    CN75_data_in(5) <= VN294_data_out(1);
    CN75_sign_in(5) <= VN294_sign_out(1);
    CN75_data_in(6) <= VN347_data_out(1);
    CN75_sign_in(6) <= VN347_sign_out(1);
    CN75_data_in(7) <= VN436_data_out(1);
    CN75_sign_in(7) <= VN436_sign_out(1);
    CN75_data_in(8) <= VN468_data_out(1);
    CN75_sign_in(8) <= VN468_sign_out(1);
    CN75_data_in(9) <= VN520_data_out(1);
    CN75_sign_in(9) <= VN520_sign_out(1);
    CN75_data_in(10) <= VN615_data_out(1);
    CN75_sign_in(10) <= VN615_sign_out(1);
    CN75_data_in(11) <= VN649_data_out(1);
    CN75_sign_in(11) <= VN649_sign_out(1);
    CN75_data_in(12) <= VN682_data_out(1);
    CN75_sign_in(12) <= VN682_sign_out(1);
    CN75_data_in(13) <= VN740_data_out(1);
    CN75_sign_in(13) <= VN740_sign_out(1);
    CN75_data_in(14) <= VN807_data_out(1);
    CN75_sign_in(14) <= VN807_sign_out(1);
    CN75_data_in(15) <= VN872_data_out(1);
    CN75_sign_in(15) <= VN872_sign_out(1);
    CN75_data_in(16) <= VN903_data_out(1);
    CN75_sign_in(16) <= VN903_sign_out(1);
    CN75_data_in(17) <= VN993_data_out(1);
    CN75_sign_in(17) <= VN993_sign_out(1);
    CN75_data_in(18) <= VN1004_data_out(1);
    CN75_sign_in(18) <= VN1004_sign_out(1);
    CN75_data_in(19) <= VN1102_data_out(1);
    CN75_sign_in(19) <= VN1102_sign_out(1);
    CN75_data_in(20) <= VN1155_data_out(1);
    CN75_sign_in(20) <= VN1155_sign_out(1);
    CN75_data_in(21) <= VN1183_data_out(1);
    CN75_sign_in(21) <= VN1183_sign_out(1);
    CN75_data_in(22) <= VN1262_data_out(1);
    CN75_sign_in(22) <= VN1262_sign_out(1);
    CN75_data_in(23) <= VN1279_data_out(1);
    CN75_sign_in(23) <= VN1279_sign_out(1);
    CN75_data_in(24) <= VN1288_data_out(1);
    CN75_sign_in(24) <= VN1288_sign_out(1);
    CN75_data_in(25) <= VN1468_data_out(1);
    CN75_sign_in(25) <= VN1468_sign_out(1);
    CN75_data_in(26) <= VN1534_data_out(1);
    CN75_sign_in(26) <= VN1534_sign_out(1);
    CN75_data_in(27) <= VN1545_data_out(1);
    CN75_sign_in(27) <= VN1545_sign_out(1);
    CN75_data_in(28) <= VN1581_data_out(1);
    CN75_sign_in(28) <= VN1581_sign_out(1);
    CN75_data_in(29) <= VN1685_data_out(1);
    CN75_sign_in(29) <= VN1685_sign_out(1);
    CN75_data_in(30) <= VN1775_data_out(1);
    CN75_sign_in(30) <= VN1775_sign_out(1);
    CN75_data_in(31) <= VN1823_data_out(1);
    CN75_sign_in(31) <= VN1823_sign_out(1);
    CN76_data_in(0) <= VN41_data_out(1);
    CN76_sign_in(0) <= VN41_sign_out(1);
    CN76_data_in(1) <= VN106_data_out(1);
    CN76_sign_in(1) <= VN106_sign_out(1);
    CN76_data_in(2) <= VN124_data_out(1);
    CN76_sign_in(2) <= VN124_sign_out(1);
    CN76_data_in(3) <= VN174_data_out(1);
    CN76_sign_in(3) <= VN174_sign_out(1);
    CN76_data_in(4) <= VN270_data_out(1);
    CN76_sign_in(4) <= VN270_sign_out(1);
    CN76_data_in(5) <= VN332_data_out(1);
    CN76_sign_in(5) <= VN332_sign_out(1);
    CN76_data_in(6) <= VN348_data_out(1);
    CN76_sign_in(6) <= VN348_sign_out(1);
    CN76_data_in(7) <= VN408_data_out(1);
    CN76_sign_in(7) <= VN408_sign_out(1);
    CN76_data_in(8) <= VN481_data_out(1);
    CN76_sign_in(8) <= VN481_sign_out(1);
    CN76_data_in(9) <= VN509_data_out(1);
    CN76_sign_in(9) <= VN509_sign_out(1);
    CN76_data_in(10) <= VN588_data_out(1);
    CN76_sign_in(10) <= VN588_sign_out(1);
    CN76_data_in(11) <= VN619_data_out(1);
    CN76_sign_in(11) <= VN619_sign_out(1);
    CN76_data_in(12) <= VN699_data_out(1);
    CN76_sign_in(12) <= VN699_sign_out(1);
    CN76_data_in(13) <= VN761_data_out(1);
    CN76_sign_in(13) <= VN761_sign_out(1);
    CN76_data_in(14) <= VN810_data_out(1);
    CN76_sign_in(14) <= VN810_sign_out(1);
    CN76_data_in(15) <= VN835_data_out(1);
    CN76_sign_in(15) <= VN835_sign_out(1);
    CN76_data_in(16) <= VN912_data_out(1);
    CN76_sign_in(16) <= VN912_sign_out(1);
    CN76_data_in(17) <= VN997_data_out(1);
    CN76_sign_in(17) <= VN997_sign_out(1);
    CN76_data_in(18) <= VN1041_data_out(1);
    CN76_sign_in(18) <= VN1041_sign_out(1);
    CN76_data_in(19) <= VN1086_data_out(1);
    CN76_sign_in(19) <= VN1086_sign_out(1);
    CN76_data_in(20) <= VN1143_data_out(1);
    CN76_sign_in(20) <= VN1143_sign_out(1);
    CN76_data_in(21) <= VN1188_data_out(1);
    CN76_sign_in(21) <= VN1188_sign_out(1);
    CN76_data_in(22) <= VN1257_data_out(1);
    CN76_sign_in(22) <= VN1257_sign_out(1);
    CN76_data_in(23) <= VN1286_data_out(1);
    CN76_sign_in(23) <= VN1286_sign_out(1);
    CN76_data_in(24) <= VN1365_data_out(1);
    CN76_sign_in(24) <= VN1365_sign_out(1);
    CN76_data_in(25) <= VN1460_data_out(1);
    CN76_sign_in(25) <= VN1460_sign_out(1);
    CN76_data_in(26) <= VN1475_data_out(1);
    CN76_sign_in(26) <= VN1475_sign_out(1);
    CN76_data_in(27) <= VN1547_data_out(1);
    CN76_sign_in(27) <= VN1547_sign_out(1);
    CN76_data_in(28) <= VN1609_data_out(1);
    CN76_sign_in(28) <= VN1609_sign_out(1);
    CN76_data_in(29) <= VN1653_data_out(1);
    CN76_sign_in(29) <= VN1653_sign_out(1);
    CN76_data_in(30) <= VN1694_data_out(1);
    CN76_sign_in(30) <= VN1694_sign_out(1);
    CN76_data_in(31) <= VN1742_data_out(1);
    CN76_sign_in(31) <= VN1742_sign_out(1);
    CN77_data_in(0) <= VN119_data_out(1);
    CN77_sign_in(0) <= VN119_sign_out(1);
    CN77_data_in(1) <= VN185_data_out(1);
    CN77_sign_in(1) <= VN185_sign_out(1);
    CN77_data_in(2) <= VN257_data_out(1);
    CN77_sign_in(2) <= VN257_sign_out(1);
    CN77_data_in(3) <= VN293_data_out(1);
    CN77_sign_in(3) <= VN293_sign_out(1);
    CN77_data_in(4) <= VN383_data_out(1);
    CN77_sign_in(4) <= VN383_sign_out(1);
    CN77_data_in(5) <= VN423_data_out(1);
    CN77_sign_in(5) <= VN423_sign_out(1);
    CN77_data_in(6) <= VN477_data_out(1);
    CN77_sign_in(6) <= VN477_sign_out(1);
    CN77_data_in(7) <= VN523_data_out(1);
    CN77_sign_in(7) <= VN523_sign_out(1);
    CN77_data_in(8) <= VN568_data_out(1);
    CN77_sign_in(8) <= VN568_sign_out(1);
    CN77_data_in(9) <= VN624_data_out(1);
    CN77_sign_in(9) <= VN624_sign_out(1);
    CN77_data_in(10) <= VN717_data_out(1);
    CN77_sign_in(10) <= VN717_sign_out(1);
    CN77_data_in(11) <= VN722_data_out(1);
    CN77_sign_in(11) <= VN722_sign_out(1);
    CN77_data_in(12) <= VN731_data_out(1);
    CN77_sign_in(12) <= VN731_sign_out(1);
    CN77_data_in(13) <= VN797_data_out(1);
    CN77_sign_in(13) <= VN797_sign_out(1);
    CN77_data_in(14) <= VN865_data_out(1);
    CN77_sign_in(14) <= VN865_sign_out(1);
    CN77_data_in(15) <= VN908_data_out(1);
    CN77_sign_in(15) <= VN908_sign_out(1);
    CN77_data_in(16) <= VN987_data_out(1);
    CN77_sign_in(16) <= VN987_sign_out(1);
    CN77_data_in(17) <= VN1055_data_out(1);
    CN77_sign_in(17) <= VN1055_sign_out(1);
    CN77_data_in(18) <= VN1088_data_out(1);
    CN77_sign_in(18) <= VN1088_sign_out(1);
    CN77_data_in(19) <= VN1177_data_out(1);
    CN77_sign_in(19) <= VN1177_sign_out(1);
    CN77_data_in(20) <= VN1263_data_out(1);
    CN77_sign_in(20) <= VN1263_sign_out(1);
    CN77_data_in(21) <= VN1316_data_out(1);
    CN77_sign_in(21) <= VN1316_sign_out(1);
    CN77_data_in(22) <= VN1349_data_out(1);
    CN77_sign_in(22) <= VN1349_sign_out(1);
    CN77_data_in(23) <= VN1409_data_out(1);
    CN77_sign_in(23) <= VN1409_sign_out(1);
    CN77_data_in(24) <= VN1435_data_out(1);
    CN77_sign_in(24) <= VN1435_sign_out(1);
    CN77_data_in(25) <= VN1624_data_out(1);
    CN77_sign_in(25) <= VN1624_sign_out(1);
    CN77_data_in(26) <= VN1659_data_out(1);
    CN77_sign_in(26) <= VN1659_sign_out(1);
    CN77_data_in(27) <= VN1810_data_out(1);
    CN77_sign_in(27) <= VN1810_sign_out(1);
    CN77_data_in(28) <= VN1845_data_out(1);
    CN77_sign_in(28) <= VN1845_sign_out(1);
    CN77_data_in(29) <= VN2013_data_out(1);
    CN77_sign_in(29) <= VN2013_sign_out(1);
    CN77_data_in(30) <= VN2017_data_out(1);
    CN77_sign_in(30) <= VN2017_sign_out(1);
    CN77_data_in(31) <= VN2031_data_out(1);
    CN77_sign_in(31) <= VN2031_sign_out(1);
    CN78_data_in(0) <= VN40_data_out(1);
    CN78_sign_in(0) <= VN40_sign_out(1);
    CN78_data_in(1) <= VN84_data_out(1);
    CN78_sign_in(1) <= VN84_sign_out(1);
    CN78_data_in(2) <= VN159_data_out(1);
    CN78_sign_in(2) <= VN159_sign_out(1);
    CN78_data_in(3) <= VN193_data_out(1);
    CN78_sign_in(3) <= VN193_sign_out(1);
    CN78_data_in(4) <= VN274_data_out(1);
    CN78_sign_in(4) <= VN274_sign_out(1);
    CN78_data_in(5) <= VN288_data_out(1);
    CN78_sign_in(5) <= VN288_sign_out(1);
    CN78_data_in(6) <= VN374_data_out(1);
    CN78_sign_in(6) <= VN374_sign_out(1);
    CN78_data_in(7) <= VN391_data_out(1);
    CN78_sign_in(7) <= VN391_sign_out(1);
    CN78_data_in(8) <= VN395_data_out(1);
    CN78_sign_in(8) <= VN395_sign_out(1);
    CN78_data_in(9) <= VN496_data_out(1);
    CN78_sign_in(9) <= VN496_sign_out(1);
    CN78_data_in(10) <= VN544_data_out(1);
    CN78_sign_in(10) <= VN544_sign_out(1);
    CN78_data_in(11) <= VN590_data_out(1);
    CN78_sign_in(11) <= VN590_sign_out(1);
    CN78_data_in(12) <= VN662_data_out(1);
    CN78_sign_in(12) <= VN662_sign_out(1);
    CN78_data_in(13) <= VN672_data_out(1);
    CN78_sign_in(13) <= VN672_sign_out(1);
    CN78_data_in(14) <= VN772_data_out(1);
    CN78_sign_in(14) <= VN772_sign_out(1);
    CN78_data_in(15) <= VN827_data_out(1);
    CN78_sign_in(15) <= VN827_sign_out(1);
    CN78_data_in(16) <= VN863_data_out(1);
    CN78_sign_in(16) <= VN863_sign_out(1);
    CN78_data_in(17) <= VN913_data_out(1);
    CN78_sign_in(17) <= VN913_sign_out(1);
    CN78_data_in(18) <= VN965_data_out(1);
    CN78_sign_in(18) <= VN965_sign_out(1);
    CN78_data_in(19) <= VN1009_data_out(1);
    CN78_sign_in(19) <= VN1009_sign_out(1);
    CN78_data_in(20) <= VN1076_data_out(1);
    CN78_sign_in(20) <= VN1076_sign_out(1);
    CN78_data_in(21) <= VN1146_data_out(1);
    CN78_sign_in(21) <= VN1146_sign_out(1);
    CN78_data_in(22) <= VN1200_data_out(1);
    CN78_sign_in(22) <= VN1200_sign_out(1);
    CN78_data_in(23) <= VN1253_data_out(1);
    CN78_sign_in(23) <= VN1253_sign_out(1);
    CN78_data_in(24) <= VN1300_data_out(1);
    CN78_sign_in(24) <= VN1300_sign_out(1);
    CN78_data_in(25) <= VN1361_data_out(1);
    CN78_sign_in(25) <= VN1361_sign_out(1);
    CN78_data_in(26) <= VN1392_data_out(1);
    CN78_sign_in(26) <= VN1392_sign_out(1);
    CN78_data_in(27) <= VN1437_data_out(1);
    CN78_sign_in(27) <= VN1437_sign_out(1);
    CN78_data_in(28) <= VN1593_data_out(1);
    CN78_sign_in(28) <= VN1593_sign_out(1);
    CN78_data_in(29) <= VN1616_data_out(1);
    CN78_sign_in(29) <= VN1616_sign_out(1);
    CN78_data_in(30) <= VN1680_data_out(1);
    CN78_sign_in(30) <= VN1680_sign_out(1);
    CN78_data_in(31) <= VN1743_data_out(1);
    CN78_sign_in(31) <= VN1743_sign_out(1);
    CN79_data_in(0) <= VN39_data_out(1);
    CN79_sign_in(0) <= VN39_sign_out(1);
    CN79_data_in(1) <= VN99_data_out(1);
    CN79_sign_in(1) <= VN99_sign_out(1);
    CN79_data_in(2) <= VN167_data_out(1);
    CN79_sign_in(2) <= VN167_sign_out(1);
    CN79_data_in(3) <= VN220_data_out(1);
    CN79_sign_in(3) <= VN220_sign_out(1);
    CN79_data_in(4) <= VN325_data_out(1);
    CN79_sign_in(4) <= VN325_sign_out(1);
    CN79_data_in(5) <= VN430_data_out(1);
    CN79_sign_in(5) <= VN430_sign_out(1);
    CN79_data_in(6) <= VN463_data_out(1);
    CN79_sign_in(6) <= VN463_sign_out(1);
    CN79_data_in(7) <= VN721_data_out(1);
    CN79_sign_in(7) <= VN721_sign_out(1);
    CN79_data_in(8) <= VN742_data_out(1);
    CN79_sign_in(8) <= VN742_sign_out(1);
    CN79_data_in(9) <= VN794_data_out(1);
    CN79_sign_in(9) <= VN794_sign_out(1);
    CN79_data_in(10) <= VN902_data_out(1);
    CN79_sign_in(10) <= VN902_sign_out(1);
    CN79_data_in(11) <= VN947_data_out(1);
    CN79_sign_in(11) <= VN947_sign_out(1);
    CN79_data_in(12) <= VN1035_data_out(1);
    CN79_sign_in(12) <= VN1035_sign_out(1);
    CN79_data_in(13) <= VN1103_data_out(1);
    CN79_sign_in(13) <= VN1103_sign_out(1);
    CN79_data_in(14) <= VN1207_data_out(1);
    CN79_sign_in(14) <= VN1207_sign_out(1);
    CN79_data_in(15) <= VN1331_data_out(1);
    CN79_sign_in(15) <= VN1331_sign_out(1);
    CN79_data_in(16) <= VN1371_data_out(1);
    CN79_sign_in(16) <= VN1371_sign_out(1);
    CN79_data_in(17) <= VN1401_data_out(1);
    CN79_sign_in(17) <= VN1401_sign_out(1);
    CN79_data_in(18) <= VN1512_data_out(1);
    CN79_sign_in(18) <= VN1512_sign_out(1);
    CN79_data_in(19) <= VN1521_data_out(1);
    CN79_sign_in(19) <= VN1521_sign_out(1);
    CN79_data_in(20) <= VN1567_data_out(1);
    CN79_sign_in(20) <= VN1567_sign_out(1);
    CN79_data_in(21) <= VN1727_data_out(1);
    CN79_sign_in(21) <= VN1727_sign_out(1);
    CN79_data_in(22) <= VN1769_data_out(1);
    CN79_sign_in(22) <= VN1769_sign_out(1);
    CN79_data_in(23) <= VN1776_data_out(1);
    CN79_sign_in(23) <= VN1776_sign_out(1);
    CN79_data_in(24) <= VN1777_data_out(1);
    CN79_sign_in(24) <= VN1777_sign_out(1);
    CN79_data_in(25) <= VN1801_data_out(1);
    CN79_sign_in(25) <= VN1801_sign_out(1);
    CN79_data_in(26) <= VN1866_data_out(1);
    CN79_sign_in(26) <= VN1866_sign_out(1);
    CN79_data_in(27) <= VN1883_data_out(1);
    CN79_sign_in(27) <= VN1883_sign_out(1);
    CN79_data_in(28) <= VN1891_data_out(1);
    CN79_sign_in(28) <= VN1891_sign_out(1);
    CN79_data_in(29) <= VN1950_data_out(1);
    CN79_sign_in(29) <= VN1950_sign_out(1);
    CN79_data_in(30) <= VN2026_data_out(1);
    CN79_sign_in(30) <= VN2026_sign_out(1);
    CN79_data_in(31) <= VN2032_data_out(1);
    CN79_sign_in(31) <= VN2032_sign_out(1);
    CN80_data_in(0) <= VN38_data_out(1);
    CN80_sign_in(0) <= VN38_sign_out(1);
    CN80_data_in(1) <= VN62_data_out(1);
    CN80_sign_in(1) <= VN62_sign_out(1);
    CN80_data_in(2) <= VN131_data_out(1);
    CN80_sign_in(2) <= VN131_sign_out(1);
    CN80_data_in(3) <= VN182_data_out(1);
    CN80_sign_in(3) <= VN182_sign_out(1);
    CN80_data_in(4) <= VN248_data_out(1);
    CN80_sign_in(4) <= VN248_sign_out(1);
    CN80_data_in(5) <= VN337_data_out(1);
    CN80_sign_in(5) <= VN337_sign_out(1);
    CN80_data_in(6) <= VN397_data_out(1);
    CN80_sign_in(6) <= VN397_sign_out(1);
    CN80_data_in(7) <= VN549_data_out(1);
    CN80_sign_in(7) <= VN549_sign_out(1);
    CN80_data_in(8) <= VN600_data_out(1);
    CN80_sign_in(8) <= VN600_sign_out(1);
    CN80_data_in(9) <= VN632_data_out(1);
    CN80_sign_in(9) <= VN632_sign_out(1);
    CN80_data_in(10) <= VN673_data_out(1);
    CN80_sign_in(10) <= VN673_sign_out(1);
    CN80_data_in(11) <= VN733_data_out(1);
    CN80_sign_in(11) <= VN733_sign_out(1);
    CN80_data_in(12) <= VN869_data_out(1);
    CN80_sign_in(12) <= VN869_sign_out(1);
    CN80_data_in(13) <= VN926_data_out(1);
    CN80_sign_in(13) <= VN926_sign_out(1);
    CN80_data_in(14) <= VN961_data_out(1);
    CN80_sign_in(14) <= VN961_sign_out(1);
    CN80_data_in(15) <= VN1072_data_out(1);
    CN80_sign_in(15) <= VN1072_sign_out(1);
    CN80_data_in(16) <= VN1118_data_out(1);
    CN80_sign_in(16) <= VN1118_sign_out(1);
    CN80_data_in(17) <= VN1166_data_out(1);
    CN80_sign_in(17) <= VN1166_sign_out(1);
    CN80_data_in(18) <= VN1192_data_out(1);
    CN80_sign_in(18) <= VN1192_sign_out(1);
    CN80_data_in(19) <= VN1228_data_out(1);
    CN80_sign_in(19) <= VN1228_sign_out(1);
    CN80_data_in(20) <= VN1289_data_out(1);
    CN80_sign_in(20) <= VN1289_sign_out(1);
    CN80_data_in(21) <= VN1343_data_out(1);
    CN80_sign_in(21) <= VN1343_sign_out(1);
    CN80_data_in(22) <= VN1410_data_out(1);
    CN80_sign_in(22) <= VN1410_sign_out(1);
    CN80_data_in(23) <= VN1461_data_out(1);
    CN80_sign_in(23) <= VN1461_sign_out(1);
    CN80_data_in(24) <= VN1484_data_out(1);
    CN80_sign_in(24) <= VN1484_sign_out(1);
    CN80_data_in(25) <= VN1695_data_out(1);
    CN80_sign_in(25) <= VN1695_sign_out(1);
    CN80_data_in(26) <= VN1730_data_out(1);
    CN80_sign_in(26) <= VN1730_sign_out(1);
    CN80_data_in(27) <= VN1915_data_out(1);
    CN80_sign_in(27) <= VN1915_sign_out(1);
    CN80_data_in(28) <= VN1961_data_out(1);
    CN80_sign_in(28) <= VN1961_sign_out(1);
    CN80_data_in(29) <= VN1967_data_out(1);
    CN80_sign_in(29) <= VN1967_sign_out(1);
    CN80_data_in(30) <= VN2010_data_out(1);
    CN80_sign_in(30) <= VN2010_sign_out(1);
    CN80_data_in(31) <= VN2022_data_out(1);
    CN80_sign_in(31) <= VN2022_sign_out(1);
    CN81_data_in(0) <= VN37_data_out(1);
    CN81_sign_in(0) <= VN37_sign_out(1);
    CN81_data_in(1) <= VN72_data_out(1);
    CN81_sign_in(1) <= VN72_sign_out(1);
    CN81_data_in(2) <= VN129_data_out(1);
    CN81_sign_in(2) <= VN129_sign_out(1);
    CN81_data_in(3) <= VN262_data_out(1);
    CN81_sign_in(3) <= VN262_sign_out(1);
    CN81_data_in(4) <= VN409_data_out(1);
    CN81_sign_in(4) <= VN409_sign_out(1);
    CN81_data_in(5) <= VN495_data_out(1);
    CN81_sign_in(5) <= VN495_sign_out(1);
    CN81_data_in(6) <= VN554_data_out(1);
    CN81_sign_in(6) <= VN554_sign_out(1);
    CN81_data_in(7) <= VN563_data_out(1);
    CN81_sign_in(7) <= VN563_sign_out(1);
    CN81_data_in(8) <= VN617_data_out(1);
    CN81_sign_in(8) <= VN617_sign_out(1);
    CN81_data_in(9) <= VN804_data_out(1);
    CN81_sign_in(9) <= VN804_sign_out(1);
    CN81_data_in(10) <= VN846_data_out(1);
    CN81_sign_in(10) <= VN846_sign_out(1);
    CN81_data_in(11) <= VN972_data_out(1);
    CN81_sign_in(11) <= VN972_sign_out(1);
    CN81_data_in(12) <= VN1012_data_out(1);
    CN81_sign_in(12) <= VN1012_sign_out(1);
    CN81_data_in(13) <= VN1095_data_out(1);
    CN81_sign_in(13) <= VN1095_sign_out(1);
    CN81_data_in(14) <= VN1114_data_out(1);
    CN81_sign_in(14) <= VN1114_sign_out(1);
    CN81_data_in(15) <= VN1168_data_out(1);
    CN81_sign_in(15) <= VN1168_sign_out(1);
    CN81_data_in(16) <= VN1267_data_out(1);
    CN81_sign_in(16) <= VN1267_sign_out(1);
    CN81_data_in(17) <= VN1317_data_out(1);
    CN81_sign_in(17) <= VN1317_sign_out(1);
    CN81_data_in(18) <= VN1496_data_out(1);
    CN81_sign_in(18) <= VN1496_sign_out(1);
    CN81_data_in(19) <= VN1546_data_out(1);
    CN81_sign_in(19) <= VN1546_sign_out(1);
    CN81_data_in(20) <= VN1560_data_out(1);
    CN81_sign_in(20) <= VN1560_sign_out(1);
    CN81_data_in(21) <= VN1580_data_out(1);
    CN81_sign_in(21) <= VN1580_sign_out(1);
    CN81_data_in(22) <= VN1647_data_out(1);
    CN81_sign_in(22) <= VN1647_sign_out(1);
    CN81_data_in(23) <= VN1655_data_out(1);
    CN81_sign_in(23) <= VN1655_sign_out(1);
    CN81_data_in(24) <= VN1867_data_out(1);
    CN81_sign_in(24) <= VN1867_sign_out(1);
    CN81_data_in(25) <= VN1874_data_out(1);
    CN81_sign_in(25) <= VN1874_sign_out(1);
    CN81_data_in(26) <= VN1878_data_out(1);
    CN81_sign_in(26) <= VN1878_sign_out(1);
    CN81_data_in(27) <= VN1949_data_out(1);
    CN81_sign_in(27) <= VN1949_sign_out(1);
    CN81_data_in(28) <= VN1956_data_out(1);
    CN81_sign_in(28) <= VN1956_sign_out(1);
    CN81_data_in(29) <= VN1957_data_out(1);
    CN81_sign_in(29) <= VN1957_sign_out(1);
    CN81_data_in(30) <= VN1971_data_out(1);
    CN81_sign_in(30) <= VN1971_sign_out(1);
    CN81_data_in(31) <= VN1973_data_out(1);
    CN81_sign_in(31) <= VN1973_sign_out(1);
    CN82_data_in(0) <= VN36_data_out(1);
    CN82_sign_in(0) <= VN36_sign_out(1);
    CN82_data_in(1) <= VN67_data_out(1);
    CN82_sign_in(1) <= VN67_sign_out(1);
    CN82_data_in(2) <= VN165_data_out(1);
    CN82_sign_in(2) <= VN165_sign_out(1);
    CN82_data_in(3) <= VN188_data_out(1);
    CN82_sign_in(3) <= VN188_sign_out(1);
    CN82_data_in(4) <= VN254_data_out(1);
    CN82_sign_in(4) <= VN254_sign_out(1);
    CN82_data_in(5) <= VN298_data_out(1);
    CN82_sign_in(5) <= VN298_sign_out(1);
    CN82_data_in(6) <= VN336_data_out(1);
    CN82_sign_in(6) <= VN336_sign_out(1);
    CN82_data_in(7) <= VN486_data_out(1);
    CN82_sign_in(7) <= VN486_sign_out(1);
    CN82_data_in(8) <= VN543_data_out(1);
    CN82_sign_in(8) <= VN543_sign_out(1);
    CN82_data_in(9) <= VN584_data_out(1);
    CN82_sign_in(9) <= VN584_sign_out(1);
    CN82_data_in(10) <= VN626_data_out(1);
    CN82_sign_in(10) <= VN626_sign_out(1);
    CN82_data_in(11) <= VN685_data_out(1);
    CN82_sign_in(11) <= VN685_sign_out(1);
    CN82_data_in(12) <= VN738_data_out(1);
    CN82_sign_in(12) <= VN738_sign_out(1);
    CN82_data_in(13) <= VN777_data_out(1);
    CN82_sign_in(13) <= VN777_sign_out(1);
    CN82_data_in(14) <= VN829_data_out(1);
    CN82_sign_in(14) <= VN829_sign_out(1);
    CN82_data_in(15) <= VN856_data_out(1);
    CN82_sign_in(15) <= VN856_sign_out(1);
    CN82_data_in(16) <= VN916_data_out(1);
    CN82_sign_in(16) <= VN916_sign_out(1);
    CN82_data_in(17) <= VN1000_data_out(1);
    CN82_sign_in(17) <= VN1000_sign_out(1);
    CN82_data_in(18) <= VN1027_data_out(1);
    CN82_sign_in(18) <= VN1027_sign_out(1);
    CN82_data_in(19) <= VN1082_data_out(1);
    CN82_sign_in(19) <= VN1082_sign_out(1);
    CN82_data_in(20) <= VN1119_data_out(1);
    CN82_sign_in(20) <= VN1119_sign_out(1);
    CN82_data_in(21) <= VN1216_data_out(1);
    CN82_sign_in(21) <= VN1216_sign_out(1);
    CN82_data_in(22) <= VN1269_data_out(1);
    CN82_sign_in(22) <= VN1269_sign_out(1);
    CN82_data_in(23) <= VN1374_data_out(1);
    CN82_sign_in(23) <= VN1374_sign_out(1);
    CN82_data_in(24) <= VN1396_data_out(1);
    CN82_sign_in(24) <= VN1396_sign_out(1);
    CN82_data_in(25) <= VN1490_data_out(1);
    CN82_sign_in(25) <= VN1490_sign_out(1);
    CN82_data_in(26) <= VN1568_data_out(1);
    CN82_sign_in(26) <= VN1568_sign_out(1);
    CN82_data_in(27) <= VN1601_data_out(1);
    CN82_sign_in(27) <= VN1601_sign_out(1);
    CN82_data_in(28) <= VN1670_data_out(1);
    CN82_sign_in(28) <= VN1670_sign_out(1);
    CN82_data_in(29) <= VN1763_data_out(1);
    CN82_sign_in(29) <= VN1763_sign_out(1);
    CN82_data_in(30) <= VN1788_data_out(1);
    CN82_sign_in(30) <= VN1788_sign_out(1);
    CN82_data_in(31) <= VN1824_data_out(1);
    CN82_sign_in(31) <= VN1824_sign_out(1);
    CN83_data_in(0) <= VN35_data_out(1);
    CN83_sign_in(0) <= VN35_sign_out(1);
    CN83_data_in(1) <= VN73_data_out(1);
    CN83_sign_in(1) <= VN73_sign_out(1);
    CN83_data_in(2) <= VN144_data_out(1);
    CN83_sign_in(2) <= VN144_sign_out(1);
    CN83_data_in(3) <= VN208_data_out(1);
    CN83_sign_in(3) <= VN208_sign_out(1);
    CN83_data_in(4) <= VN232_data_out(1);
    CN83_sign_in(4) <= VN232_sign_out(1);
    CN83_data_in(5) <= VN330_data_out(1);
    CN83_sign_in(5) <= VN330_sign_out(1);
    CN83_data_in(6) <= VN425_data_out(1);
    CN83_sign_in(6) <= VN425_sign_out(1);
    CN83_data_in(7) <= VN448_data_out(1);
    CN83_sign_in(7) <= VN448_sign_out(1);
    CN83_data_in(8) <= VN511_data_out(1);
    CN83_sign_in(8) <= VN511_sign_out(1);
    CN83_data_in(9) <= VN585_data_out(1);
    CN83_sign_in(9) <= VN585_sign_out(1);
    CN83_data_in(10) <= VN633_data_out(1);
    CN83_sign_in(10) <= VN633_sign_out(1);
    CN83_data_in(11) <= VN691_data_out(1);
    CN83_sign_in(11) <= VN691_sign_out(1);
    CN83_data_in(12) <= VN821_data_out(1);
    CN83_sign_in(12) <= VN821_sign_out(1);
    CN83_data_in(13) <= VN850_data_out(1);
    CN83_sign_in(13) <= VN850_sign_out(1);
    CN83_data_in(14) <= VN918_data_out(1);
    CN83_sign_in(14) <= VN918_sign_out(1);
    CN83_data_in(15) <= VN989_data_out(1);
    CN83_sign_in(15) <= VN989_sign_out(1);
    CN83_data_in(16) <= VN1047_data_out(1);
    CN83_sign_in(16) <= VN1047_sign_out(1);
    CN83_data_in(17) <= VN1105_data_out(1);
    CN83_sign_in(17) <= VN1105_sign_out(1);
    CN83_data_in(18) <= VN1239_data_out(1);
    CN83_sign_in(18) <= VN1239_sign_out(1);
    CN83_data_in(19) <= VN1309_data_out(1);
    CN83_sign_in(19) <= VN1309_sign_out(1);
    CN83_data_in(20) <= VN1332_data_out(1);
    CN83_sign_in(20) <= VN1332_sign_out(1);
    CN83_data_in(21) <= VN1425_data_out(1);
    CN83_sign_in(21) <= VN1425_sign_out(1);
    CN83_data_in(22) <= VN1436_data_out(1);
    CN83_sign_in(22) <= VN1436_sign_out(1);
    CN83_data_in(23) <= VN1511_data_out(1);
    CN83_sign_in(23) <= VN1511_sign_out(1);
    CN83_data_in(24) <= VN1590_data_out(1);
    CN83_sign_in(24) <= VN1590_sign_out(1);
    CN83_data_in(25) <= VN1641_data_out(1);
    CN83_sign_in(25) <= VN1641_sign_out(1);
    CN83_data_in(26) <= VN1681_data_out(1);
    CN83_sign_in(26) <= VN1681_sign_out(1);
    CN83_data_in(27) <= VN1693_data_out(1);
    CN83_sign_in(27) <= VN1693_sign_out(1);
    CN83_data_in(28) <= VN1819_data_out(1);
    CN83_sign_in(28) <= VN1819_sign_out(1);
    CN83_data_in(29) <= VN1871_data_out(1);
    CN83_sign_in(29) <= VN1871_sign_out(1);
    CN83_data_in(30) <= VN1919_data_out(1);
    CN83_sign_in(30) <= VN1919_sign_out(1);
    CN83_data_in(31) <= VN1922_data_out(1);
    CN83_sign_in(31) <= VN1922_sign_out(1);
    CN84_data_in(0) <= VN34_data_out(1);
    CN84_sign_in(0) <= VN34_sign_out(1);
    CN84_data_in(1) <= VN61_data_out(1);
    CN84_sign_in(1) <= VN61_sign_out(1);
    CN84_data_in(2) <= VN147_data_out(1);
    CN84_sign_in(2) <= VN147_sign_out(1);
    CN84_data_in(3) <= VN222_data_out(1);
    CN84_sign_in(3) <= VN222_sign_out(1);
    CN84_data_in(4) <= VN310_data_out(1);
    CN84_sign_in(4) <= VN310_sign_out(1);
    CN84_data_in(5) <= VN371_data_out(1);
    CN84_sign_in(5) <= VN371_sign_out(1);
    CN84_data_in(6) <= VN392_data_out(1);
    CN84_sign_in(6) <= VN392_sign_out(1);
    CN84_data_in(7) <= VN453_data_out(1);
    CN84_sign_in(7) <= VN453_sign_out(1);
    CN84_data_in(8) <= VN562_data_out(1);
    CN84_sign_in(8) <= VN562_sign_out(1);
    CN84_data_in(9) <= VN663_data_out(1);
    CN84_sign_in(9) <= VN663_sign_out(1);
    CN84_data_in(10) <= VN676_data_out(1);
    CN84_sign_in(10) <= VN676_sign_out(1);
    CN84_data_in(11) <= VN766_data_out(1);
    CN84_sign_in(11) <= VN766_sign_out(1);
    CN84_data_in(12) <= VN808_data_out(1);
    CN84_sign_in(12) <= VN808_sign_out(1);
    CN84_data_in(13) <= VN854_data_out(1);
    CN84_sign_in(13) <= VN854_sign_out(1);
    CN84_data_in(14) <= VN942_data_out(1);
    CN84_sign_in(14) <= VN942_sign_out(1);
    CN84_data_in(15) <= VN975_data_out(1);
    CN84_sign_in(15) <= VN975_sign_out(1);
    CN84_data_in(16) <= VN1057_data_out(1);
    CN84_sign_in(16) <= VN1057_sign_out(1);
    CN84_data_in(17) <= VN1097_data_out(1);
    CN84_sign_in(17) <= VN1097_sign_out(1);
    CN84_data_in(18) <= VN1132_data_out(1);
    CN84_sign_in(18) <= VN1132_sign_out(1);
    CN84_data_in(19) <= VN1211_data_out(1);
    CN84_sign_in(19) <= VN1211_sign_out(1);
    CN84_data_in(20) <= VN1404_data_out(1);
    CN84_sign_in(20) <= VN1404_sign_out(1);
    CN84_data_in(21) <= VN1455_data_out(1);
    CN84_sign_in(21) <= VN1455_sign_out(1);
    CN84_data_in(22) <= VN1463_data_out(1);
    CN84_sign_in(22) <= VN1463_sign_out(1);
    CN84_data_in(23) <= VN1474_data_out(1);
    CN84_sign_in(23) <= VN1474_sign_out(1);
    CN84_data_in(24) <= VN1625_data_out(1);
    CN84_sign_in(24) <= VN1625_sign_out(1);
    CN84_data_in(25) <= VN1678_data_out(1);
    CN84_sign_in(25) <= VN1678_sign_out(1);
    CN84_data_in(26) <= VN1761_data_out(1);
    CN84_sign_in(26) <= VN1761_sign_out(1);
    CN84_data_in(27) <= VN1804_data_out(1);
    CN84_sign_in(27) <= VN1804_sign_out(1);
    CN84_data_in(28) <= VN1863_data_out(1);
    CN84_sign_in(28) <= VN1863_sign_out(1);
    CN84_data_in(29) <= VN1870_data_out(1);
    CN84_sign_in(29) <= VN1870_sign_out(1);
    CN84_data_in(30) <= VN1897_data_out(1);
    CN84_sign_in(30) <= VN1897_sign_out(1);
    CN84_data_in(31) <= VN1907_data_out(1);
    CN84_sign_in(31) <= VN1907_sign_out(1);
    CN85_data_in(0) <= VN33_data_out(1);
    CN85_sign_in(0) <= VN33_sign_out(1);
    CN85_data_in(1) <= VN132_data_out(1);
    CN85_sign_in(1) <= VN132_sign_out(1);
    CN85_data_in(2) <= VN218_data_out(1);
    CN85_sign_in(2) <= VN218_sign_out(1);
    CN85_data_in(3) <= VN235_data_out(1);
    CN85_sign_in(3) <= VN235_sign_out(1);
    CN85_data_in(4) <= VN313_data_out(1);
    CN85_sign_in(4) <= VN313_sign_out(1);
    CN85_data_in(5) <= VN379_data_out(1);
    CN85_sign_in(5) <= VN379_sign_out(1);
    CN85_data_in(6) <= VN505_data_out(1);
    CN85_sign_in(6) <= VN505_sign_out(1);
    CN85_data_in(7) <= VN558_data_out(1);
    CN85_sign_in(7) <= VN558_sign_out(1);
    CN85_data_in(8) <= VN608_data_out(1);
    CN85_sign_in(8) <= VN608_sign_out(1);
    CN85_data_in(9) <= VN623_data_out(1);
    CN85_sign_in(9) <= VN623_sign_out(1);
    CN85_data_in(10) <= VN677_data_out(1);
    CN85_sign_in(10) <= VN677_sign_out(1);
    CN85_data_in(11) <= VN725_data_out(1);
    CN85_sign_in(11) <= VN725_sign_out(1);
    CN85_data_in(12) <= VN843_data_out(1);
    CN85_sign_in(12) <= VN843_sign_out(1);
    CN85_data_in(13) <= VN924_data_out(1);
    CN85_sign_in(13) <= VN924_sign_out(1);
    CN85_data_in(14) <= VN1052_data_out(1);
    CN85_sign_in(14) <= VN1052_sign_out(1);
    CN85_data_in(15) <= VN1087_data_out(1);
    CN85_sign_in(15) <= VN1087_sign_out(1);
    CN85_data_in(16) <= VN1217_data_out(1);
    CN85_sign_in(16) <= VN1217_sign_out(1);
    CN85_data_in(17) <= VN1232_data_out(1);
    CN85_sign_in(17) <= VN1232_sign_out(1);
    CN85_data_in(18) <= VN1277_data_out(1);
    CN85_sign_in(18) <= VN1277_sign_out(1);
    CN85_data_in(19) <= VN1319_data_out(1);
    CN85_sign_in(19) <= VN1319_sign_out(1);
    CN85_data_in(20) <= VN1363_data_out(1);
    CN85_sign_in(20) <= VN1363_sign_out(1);
    CN85_data_in(21) <= VN1389_data_out(1);
    CN85_sign_in(21) <= VN1389_sign_out(1);
    CN85_data_in(22) <= VN1652_data_out(1);
    CN85_sign_in(22) <= VN1652_sign_out(1);
    CN85_data_in(23) <= VN1768_data_out(1);
    CN85_sign_in(23) <= VN1768_sign_out(1);
    CN85_data_in(24) <= VN1770_data_out(1);
    CN85_sign_in(24) <= VN1770_sign_out(1);
    CN85_data_in(25) <= VN1772_data_out(1);
    CN85_sign_in(25) <= VN1772_sign_out(1);
    CN85_data_in(26) <= VN1815_data_out(1);
    CN85_sign_in(26) <= VN1815_sign_out(1);
    CN85_data_in(27) <= VN1872_data_out(1);
    CN85_sign_in(27) <= VN1872_sign_out(1);
    CN85_data_in(28) <= VN1909_data_out(1);
    CN85_sign_in(28) <= VN1909_sign_out(1);
    CN85_data_in(29) <= VN2016_data_out(1);
    CN85_sign_in(29) <= VN2016_sign_out(1);
    CN85_data_in(30) <= VN2038_data_out(1);
    CN85_sign_in(30) <= VN2038_sign_out(1);
    CN85_data_in(31) <= VN2043_data_out(1);
    CN85_sign_in(31) <= VN2043_sign_out(1);
    CN86_data_in(0) <= VN32_data_out(1);
    CN86_sign_in(0) <= VN32_sign_out(1);
    CN86_data_in(1) <= VN166_data_out(1);
    CN86_sign_in(1) <= VN166_sign_out(1);
    CN86_data_in(2) <= VN239_data_out(1);
    CN86_sign_in(2) <= VN239_sign_out(1);
    CN86_data_in(3) <= VN343_data_out(1);
    CN86_sign_in(3) <= VN343_sign_out(1);
    CN86_data_in(4) <= VN424_data_out(1);
    CN86_sign_in(4) <= VN424_sign_out(1);
    CN86_data_in(5) <= VN452_data_out(1);
    CN86_sign_in(5) <= VN452_sign_out(1);
    CN86_data_in(6) <= VN559_data_out(1);
    CN86_sign_in(6) <= VN559_sign_out(1);
    CN86_data_in(7) <= VN571_data_out(1);
    CN86_sign_in(7) <= VN571_sign_out(1);
    CN86_data_in(8) <= VN651_data_out(1);
    CN86_sign_in(8) <= VN651_sign_out(1);
    CN86_data_in(9) <= VN703_data_out(1);
    CN86_sign_in(9) <= VN703_sign_out(1);
    CN86_data_in(10) <= VN773_data_out(1);
    CN86_sign_in(10) <= VN773_sign_out(1);
    CN86_data_in(11) <= VN877_data_out(1);
    CN86_sign_in(11) <= VN877_sign_out(1);
    CN86_data_in(12) <= VN934_data_out(1);
    CN86_sign_in(12) <= VN934_sign_out(1);
    CN86_data_in(13) <= VN953_data_out(1);
    CN86_sign_in(13) <= VN953_sign_out(1);
    CN86_data_in(14) <= VN1058_data_out(1);
    CN86_sign_in(14) <= VN1058_sign_out(1);
    CN86_data_in(15) <= VN1101_data_out(1);
    CN86_sign_in(15) <= VN1101_sign_out(1);
    CN86_data_in(16) <= VN1112_data_out(1);
    CN86_sign_in(16) <= VN1112_sign_out(1);
    CN86_data_in(17) <= VN1122_data_out(1);
    CN86_sign_in(17) <= VN1122_sign_out(1);
    CN86_data_in(18) <= VN1310_data_out(1);
    CN86_sign_in(18) <= VN1310_sign_out(1);
    CN86_data_in(19) <= VN1358_data_out(1);
    CN86_sign_in(19) <= VN1358_sign_out(1);
    CN86_data_in(20) <= VN1620_data_out(1);
    CN86_sign_in(20) <= VN1620_sign_out(1);
    CN86_data_in(21) <= VN1756_data_out(1);
    CN86_sign_in(21) <= VN1756_sign_out(1);
    CN86_data_in(22) <= VN1762_data_out(1);
    CN86_sign_in(22) <= VN1762_sign_out(1);
    CN86_data_in(23) <= VN1802_data_out(1);
    CN86_sign_in(23) <= VN1802_sign_out(1);
    CN86_data_in(24) <= VN1916_data_out(1);
    CN86_sign_in(24) <= VN1916_sign_out(1);
    CN86_data_in(25) <= VN1944_data_out(1);
    CN86_sign_in(25) <= VN1944_sign_out(1);
    CN86_data_in(26) <= VN1946_data_out(1);
    CN86_sign_in(26) <= VN1946_sign_out(1);
    CN86_data_in(27) <= VN1954_data_out(1);
    CN86_sign_in(27) <= VN1954_sign_out(1);
    CN86_data_in(28) <= VN1983_data_out(1);
    CN86_sign_in(28) <= VN1983_sign_out(1);
    CN86_data_in(29) <= VN1993_data_out(1);
    CN86_sign_in(29) <= VN1993_sign_out(1);
    CN86_data_in(30) <= VN1996_data_out(1);
    CN86_sign_in(30) <= VN1996_sign_out(1);
    CN86_data_in(31) <= VN2001_data_out(1);
    CN86_sign_in(31) <= VN2001_sign_out(1);
    CN87_data_in(0) <= VN31_data_out(1);
    CN87_sign_in(0) <= VN31_sign_out(1);
    CN87_data_in(1) <= VN77_data_out(1);
    CN87_sign_in(1) <= VN77_sign_out(1);
    CN87_data_in(2) <= VN128_data_out(1);
    CN87_sign_in(2) <= VN128_sign_out(1);
    CN87_data_in(3) <= VN203_data_out(1);
    CN87_sign_in(3) <= VN203_sign_out(1);
    CN87_data_in(4) <= VN229_data_out(1);
    CN87_sign_in(4) <= VN229_sign_out(1);
    CN87_data_in(5) <= VN331_data_out(1);
    CN87_sign_in(5) <= VN331_sign_out(1);
    CN87_data_in(6) <= VN341_data_out(1);
    CN87_sign_in(6) <= VN341_sign_out(1);
    CN87_data_in(7) <= VN416_data_out(1);
    CN87_sign_in(7) <= VN416_sign_out(1);
    CN87_data_in(8) <= VN503_data_out(1);
    CN87_sign_in(8) <= VN503_sign_out(1);
    CN87_data_in(9) <= VN526_data_out(1);
    CN87_sign_in(9) <= VN526_sign_out(1);
    CN87_data_in(10) <= VN576_data_out(1);
    CN87_sign_in(10) <= VN576_sign_out(1);
    CN87_data_in(11) <= VN683_data_out(1);
    CN87_sign_in(11) <= VN683_sign_out(1);
    CN87_data_in(12) <= VN799_data_out(1);
    CN87_sign_in(12) <= VN799_sign_out(1);
    CN87_data_in(13) <= VN862_data_out(1);
    CN87_sign_in(13) <= VN862_sign_out(1);
    CN87_data_in(14) <= VN963_data_out(1);
    CN87_sign_in(14) <= VN963_sign_out(1);
    CN87_data_in(15) <= VN1046_data_out(1);
    CN87_sign_in(15) <= VN1046_sign_out(1);
    CN87_data_in(16) <= VN1124_data_out(1);
    CN87_sign_in(16) <= VN1124_sign_out(1);
    CN87_data_in(17) <= VN1206_data_out(1);
    CN87_sign_in(17) <= VN1206_sign_out(1);
    CN87_data_in(18) <= VN1268_data_out(1);
    CN87_sign_in(18) <= VN1268_sign_out(1);
    CN87_data_in(19) <= VN1426_data_out(1);
    CN87_sign_in(19) <= VN1426_sign_out(1);
    CN87_data_in(20) <= VN1459_data_out(1);
    CN87_sign_in(20) <= VN1459_sign_out(1);
    CN87_data_in(21) <= VN1544_data_out(1);
    CN87_sign_in(21) <= VN1544_sign_out(1);
    CN87_data_in(22) <= VN1554_data_out(1);
    CN87_sign_in(22) <= VN1554_sign_out(1);
    CN87_data_in(23) <= VN1731_data_out(1);
    CN87_sign_in(23) <= VN1731_sign_out(1);
    CN87_data_in(24) <= VN1765_data_out(1);
    CN87_sign_in(24) <= VN1765_sign_out(1);
    CN87_data_in(25) <= VN1832_data_out(1);
    CN87_sign_in(25) <= VN1832_sign_out(1);
    CN87_data_in(26) <= VN1842_data_out(1);
    CN87_sign_in(26) <= VN1842_sign_out(1);
    CN87_data_in(27) <= VN1853_data_out(1);
    CN87_sign_in(27) <= VN1853_sign_out(1);
    CN87_data_in(28) <= VN1869_data_out(1);
    CN87_sign_in(28) <= VN1869_sign_out(1);
    CN87_data_in(29) <= VN1917_data_out(1);
    CN87_sign_in(29) <= VN1917_sign_out(1);
    CN87_data_in(30) <= VN2000_data_out(1);
    CN87_sign_in(30) <= VN2000_sign_out(1);
    CN87_data_in(31) <= VN2005_data_out(1);
    CN87_sign_in(31) <= VN2005_sign_out(1);
    CN88_data_in(0) <= VN30_data_out(1);
    CN88_sign_in(0) <= VN30_sign_out(1);
    CN88_data_in(1) <= VN79_data_out(1);
    CN88_sign_in(1) <= VN79_sign_out(1);
    CN88_data_in(2) <= VN156_data_out(1);
    CN88_sign_in(2) <= VN156_sign_out(1);
    CN88_data_in(3) <= VN204_data_out(1);
    CN88_sign_in(3) <= VN204_sign_out(1);
    CN88_data_in(4) <= VN263_data_out(1);
    CN88_sign_in(4) <= VN263_sign_out(1);
    CN88_data_in(5) <= VN297_data_out(1);
    CN88_sign_in(5) <= VN297_sign_out(1);
    CN88_data_in(6) <= VN377_data_out(1);
    CN88_sign_in(6) <= VN377_sign_out(1);
    CN88_data_in(7) <= VN434_data_out(1);
    CN88_sign_in(7) <= VN434_sign_out(1);
    CN88_data_in(8) <= VN484_data_out(1);
    CN88_sign_in(8) <= VN484_sign_out(1);
    CN88_data_in(9) <= VN616_data_out(1);
    CN88_sign_in(9) <= VN616_sign_out(1);
    CN88_data_in(10) <= VN695_data_out(1);
    CN88_sign_in(10) <= VN695_sign_out(1);
    CN88_data_in(11) <= VN759_data_out(1);
    CN88_sign_in(11) <= VN759_sign_out(1);
    CN88_data_in(12) <= VN813_data_out(1);
    CN88_sign_in(12) <= VN813_sign_out(1);
    CN88_data_in(13) <= VN873_data_out(1);
    CN88_sign_in(13) <= VN873_sign_out(1);
    CN88_data_in(14) <= VN917_data_out(1);
    CN88_sign_in(14) <= VN917_sign_out(1);
    CN88_data_in(15) <= VN958_data_out(1);
    CN88_sign_in(15) <= VN958_sign_out(1);
    CN88_data_in(16) <= VN1014_data_out(1);
    CN88_sign_in(16) <= VN1014_sign_out(1);
    CN88_data_in(17) <= VN1150_data_out(1);
    CN88_sign_in(17) <= VN1150_sign_out(1);
    CN88_data_in(18) <= VN1179_data_out(1);
    CN88_sign_in(18) <= VN1179_sign_out(1);
    CN88_data_in(19) <= VN1227_data_out(1);
    CN88_sign_in(19) <= VN1227_sign_out(1);
    CN88_data_in(20) <= VN1278_data_out(1);
    CN88_sign_in(20) <= VN1278_sign_out(1);
    CN88_data_in(21) <= VN1315_data_out(1);
    CN88_sign_in(21) <= VN1315_sign_out(1);
    CN88_data_in(22) <= VN1354_data_out(1);
    CN88_sign_in(22) <= VN1354_sign_out(1);
    CN88_data_in(23) <= VN1399_data_out(1);
    CN88_sign_in(23) <= VN1399_sign_out(1);
    CN88_data_in(24) <= VN1438_data_out(1);
    CN88_sign_in(24) <= VN1438_sign_out(1);
    CN88_data_in(25) <= VN1700_data_out(1);
    CN88_sign_in(25) <= VN1700_sign_out(1);
    CN88_data_in(26) <= VN1799_data_out(1);
    CN88_sign_in(26) <= VN1799_sign_out(1);
    CN88_data_in(27) <= VN1903_data_out(1);
    CN88_sign_in(27) <= VN1903_sign_out(1);
    CN88_data_in(28) <= VN1911_data_out(1);
    CN88_sign_in(28) <= VN1911_sign_out(1);
    CN88_data_in(29) <= VN1929_data_out(1);
    CN88_sign_in(29) <= VN1929_sign_out(1);
    CN88_data_in(30) <= VN2037_data_out(1);
    CN88_sign_in(30) <= VN2037_sign_out(1);
    CN88_data_in(31) <= VN2040_data_out(1);
    CN88_sign_in(31) <= VN2040_sign_out(1);
    CN89_data_in(0) <= VN29_data_out(1);
    CN89_sign_in(0) <= VN29_sign_out(1);
    CN89_data_in(1) <= VN102_data_out(1);
    CN89_sign_in(1) <= VN102_sign_out(1);
    CN89_data_in(2) <= VN140_data_out(1);
    CN89_sign_in(2) <= VN140_sign_out(1);
    CN89_data_in(3) <= VN184_data_out(1);
    CN89_sign_in(3) <= VN184_sign_out(1);
    CN89_data_in(4) <= VN247_data_out(1);
    CN89_sign_in(4) <= VN247_sign_out(1);
    CN89_data_in(5) <= VN355_data_out(1);
    CN89_sign_in(5) <= VN355_sign_out(1);
    CN89_data_in(6) <= VN438_data_out(1);
    CN89_sign_in(6) <= VN438_sign_out(1);
    CN89_data_in(7) <= VN491_data_out(1);
    CN89_sign_in(7) <= VN491_sign_out(1);
    CN89_data_in(8) <= VN519_data_out(1);
    CN89_sign_in(8) <= VN519_sign_out(1);
    CN89_data_in(9) <= VN575_data_out(1);
    CN89_sign_in(9) <= VN575_sign_out(1);
    CN89_data_in(10) <= VN664_data_out(1);
    CN89_sign_in(10) <= VN664_sign_out(1);
    CN89_data_in(11) <= VN704_data_out(1);
    CN89_sign_in(11) <= VN704_sign_out(1);
    CN89_data_in(12) <= VN752_data_out(1);
    CN89_sign_in(12) <= VN752_sign_out(1);
    CN89_data_in(13) <= VN884_data_out(1);
    CN89_sign_in(13) <= VN884_sign_out(1);
    CN89_data_in(14) <= VN1130_data_out(1);
    CN89_sign_in(14) <= VN1130_sign_out(1);
    CN89_data_in(15) <= VN1167_data_out(1);
    CN89_sign_in(15) <= VN1167_sign_out(1);
    CN89_data_in(16) <= VN1213_data_out(1);
    CN89_sign_in(16) <= VN1213_sign_out(1);
    CN89_data_in(17) <= VN1293_data_out(1);
    CN89_sign_in(17) <= VN1293_sign_out(1);
    CN89_data_in(18) <= VN1377_data_out(1);
    CN89_sign_in(18) <= VN1377_sign_out(1);
    CN89_data_in(19) <= VN1421_data_out(1);
    CN89_sign_in(19) <= VN1421_sign_out(1);
    CN89_data_in(20) <= VN1585_data_out(1);
    CN89_sign_in(20) <= VN1585_sign_out(1);
    CN89_data_in(21) <= VN1643_data_out(1);
    CN89_sign_in(21) <= VN1643_sign_out(1);
    CN89_data_in(22) <= VN1686_data_out(1);
    CN89_sign_in(22) <= VN1686_sign_out(1);
    CN89_data_in(23) <= VN1725_data_out(1);
    CN89_sign_in(23) <= VN1725_sign_out(1);
    CN89_data_in(24) <= VN1861_data_out(1);
    CN89_sign_in(24) <= VN1861_sign_out(1);
    CN89_data_in(25) <= VN1892_data_out(1);
    CN89_sign_in(25) <= VN1892_sign_out(1);
    CN89_data_in(26) <= VN1894_data_out(1);
    CN89_sign_in(26) <= VN1894_sign_out(1);
    CN89_data_in(27) <= VN1918_data_out(1);
    CN89_sign_in(27) <= VN1918_sign_out(1);
    CN89_data_in(28) <= VN1935_data_out(1);
    CN89_sign_in(28) <= VN1935_sign_out(1);
    CN89_data_in(29) <= VN1972_data_out(1);
    CN89_sign_in(29) <= VN1972_sign_out(1);
    CN89_data_in(30) <= VN2025_data_out(1);
    CN89_sign_in(30) <= VN2025_sign_out(1);
    CN89_data_in(31) <= VN2033_data_out(1);
    CN89_sign_in(31) <= VN2033_sign_out(1);
    CN90_data_in(0) <= VN28_data_out(1);
    CN90_sign_in(0) <= VN28_sign_out(1);
    CN90_data_in(1) <= VN85_data_out(1);
    CN90_sign_in(1) <= VN85_sign_out(1);
    CN90_data_in(2) <= VN168_data_out(1);
    CN90_sign_in(2) <= VN168_sign_out(1);
    CN90_data_in(3) <= VN175_data_out(1);
    CN90_sign_in(3) <= VN175_sign_out(1);
    CN90_data_in(4) <= VN258_data_out(1);
    CN90_sign_in(4) <= VN258_sign_out(1);
    CN90_data_in(5) <= VN307_data_out(1);
    CN90_sign_in(5) <= VN307_sign_out(1);
    CN90_data_in(6) <= VN358_data_out(1);
    CN90_sign_in(6) <= VN358_sign_out(1);
    CN90_data_in(7) <= VN447_data_out(1);
    CN90_sign_in(7) <= VN447_sign_out(1);
    CN90_data_in(8) <= VN459_data_out(1);
    CN90_sign_in(8) <= VN459_sign_out(1);
    CN90_data_in(9) <= VN527_data_out(1);
    CN90_sign_in(9) <= VN527_sign_out(1);
    CN90_data_in(10) <= VN661_data_out(1);
    CN90_sign_in(10) <= VN661_sign_out(1);
    CN90_data_in(11) <= VN756_data_out(1);
    CN90_sign_in(11) <= VN756_sign_out(1);
    CN90_data_in(12) <= VN783_data_out(1);
    CN90_sign_in(12) <= VN783_sign_out(1);
    CN90_data_in(13) <= VN904_data_out(1);
    CN90_sign_in(13) <= VN904_sign_out(1);
    CN90_data_in(14) <= VN952_data_out(1);
    CN90_sign_in(14) <= VN952_sign_out(1);
    CN90_data_in(15) <= VN1084_data_out(1);
    CN90_sign_in(15) <= VN1084_sign_out(1);
    CN90_data_in(16) <= VN1142_data_out(1);
    CN90_sign_in(16) <= VN1142_sign_out(1);
    CN90_data_in(17) <= VN1181_data_out(1);
    CN90_sign_in(17) <= VN1181_sign_out(1);
    CN90_data_in(18) <= VN1291_data_out(1);
    CN90_sign_in(18) <= VN1291_sign_out(1);
    CN90_data_in(19) <= VN1330_data_out(1);
    CN90_sign_in(19) <= VN1330_sign_out(1);
    CN90_data_in(20) <= VN1383_data_out(1);
    CN90_sign_in(20) <= VN1383_sign_out(1);
    CN90_data_in(21) <= VN1559_data_out(1);
    CN90_sign_in(21) <= VN1559_sign_out(1);
    CN90_data_in(22) <= VN1630_data_out(1);
    CN90_sign_in(22) <= VN1630_sign_out(1);
    CN90_data_in(23) <= VN1703_data_out(1);
    CN90_sign_in(23) <= VN1703_sign_out(1);
    CN90_data_in(24) <= VN1834_data_out(1);
    CN90_sign_in(24) <= VN1834_sign_out(1);
    CN90_data_in(25) <= VN1841_data_out(1);
    CN90_sign_in(25) <= VN1841_sign_out(1);
    CN90_data_in(26) <= VN1846_data_out(1);
    CN90_sign_in(26) <= VN1846_sign_out(1);
    CN90_data_in(27) <= VN1881_data_out(1);
    CN90_sign_in(27) <= VN1881_sign_out(1);
    CN90_data_in(28) <= VN1882_data_out(1);
    CN90_sign_in(28) <= VN1882_sign_out(1);
    CN90_data_in(29) <= VN1888_data_out(1);
    CN90_sign_in(29) <= VN1888_sign_out(1);
    CN90_data_in(30) <= VN1923_data_out(1);
    CN90_sign_in(30) <= VN1923_sign_out(1);
    CN90_data_in(31) <= VN1925_data_out(1);
    CN90_sign_in(31) <= VN1925_sign_out(1);
    CN91_data_in(0) <= VN27_data_out(1);
    CN91_sign_in(0) <= VN27_sign_out(1);
    CN91_data_in(1) <= VN96_data_out(1);
    CN91_sign_in(1) <= VN96_sign_out(1);
    CN91_data_in(2) <= VN158_data_out(1);
    CN91_sign_in(2) <= VN158_sign_out(1);
    CN91_data_in(3) <= VN191_data_out(1);
    CN91_sign_in(3) <= VN191_sign_out(1);
    CN91_data_in(4) <= VN269_data_out(1);
    CN91_sign_in(4) <= VN269_sign_out(1);
    CN91_data_in(5) <= VN280_data_out(1);
    CN91_sign_in(5) <= VN280_sign_out(1);
    CN91_data_in(6) <= VN344_data_out(1);
    CN91_sign_in(6) <= VN344_sign_out(1);
    CN91_data_in(7) <= VN457_data_out(1);
    CN91_sign_in(7) <= VN457_sign_out(1);
    CN91_data_in(8) <= VN606_data_out(1);
    CN91_sign_in(8) <= VN606_sign_out(1);
    CN91_data_in(9) <= VN690_data_out(1);
    CN91_sign_in(9) <= VN690_sign_out(1);
    CN91_data_in(10) <= VN746_data_out(1);
    CN91_sign_in(10) <= VN746_sign_out(1);
    CN91_data_in(11) <= VN792_data_out(1);
    CN91_sign_in(11) <= VN792_sign_out(1);
    CN91_data_in(12) <= VN845_data_out(1);
    CN91_sign_in(12) <= VN845_sign_out(1);
    CN91_data_in(13) <= VN937_data_out(1);
    CN91_sign_in(13) <= VN937_sign_out(1);
    CN91_data_in(14) <= VN978_data_out(1);
    CN91_sign_in(14) <= VN978_sign_out(1);
    CN91_data_in(15) <= VN1007_data_out(1);
    CN91_sign_in(15) <= VN1007_sign_out(1);
    CN91_data_in(16) <= VN1059_data_out(1);
    CN91_sign_in(16) <= VN1059_sign_out(1);
    CN91_data_in(17) <= VN1151_data_out(1);
    CN91_sign_in(17) <= VN1151_sign_out(1);
    CN91_data_in(18) <= VN1193_data_out(1);
    CN91_sign_in(18) <= VN1193_sign_out(1);
    CN91_data_in(19) <= VN1256_data_out(1);
    CN91_sign_in(19) <= VN1256_sign_out(1);
    CN91_data_in(20) <= VN1367_data_out(1);
    CN91_sign_in(20) <= VN1367_sign_out(1);
    CN91_data_in(21) <= VN1384_data_out(1);
    CN91_sign_in(21) <= VN1384_sign_out(1);
    CN91_data_in(22) <= VN1398_data_out(1);
    CN91_sign_in(22) <= VN1398_sign_out(1);
    CN91_data_in(23) <= VN1591_data_out(1);
    CN91_sign_in(23) <= VN1591_sign_out(1);
    CN91_data_in(24) <= VN1645_data_out(1);
    CN91_sign_in(24) <= VN1645_sign_out(1);
    CN91_data_in(25) <= VN1733_data_out(1);
    CN91_sign_in(25) <= VN1733_sign_out(1);
    CN91_data_in(26) <= VN1792_data_out(1);
    CN91_sign_in(26) <= VN1792_sign_out(1);
    CN91_data_in(27) <= VN1905_data_out(1);
    CN91_sign_in(27) <= VN1905_sign_out(1);
    CN91_data_in(28) <= VN1979_data_out(1);
    CN91_sign_in(28) <= VN1979_sign_out(1);
    CN91_data_in(29) <= VN1999_data_out(1);
    CN91_sign_in(29) <= VN1999_sign_out(1);
    CN91_data_in(30) <= VN2028_data_out(1);
    CN91_sign_in(30) <= VN2028_sign_out(1);
    CN91_data_in(31) <= VN2034_data_out(1);
    CN91_sign_in(31) <= VN2034_sign_out(1);
    CN92_data_in(0) <= VN26_data_out(1);
    CN92_sign_in(0) <= VN26_sign_out(1);
    CN92_data_in(1) <= VN103_data_out(1);
    CN92_sign_in(1) <= VN103_sign_out(1);
    CN92_data_in(2) <= VN145_data_out(1);
    CN92_sign_in(2) <= VN145_sign_out(1);
    CN92_data_in(3) <= VN195_data_out(1);
    CN92_sign_in(3) <= VN195_sign_out(1);
    CN92_data_in(4) <= VN242_data_out(1);
    CN92_sign_in(4) <= VN242_sign_out(1);
    CN92_data_in(5) <= VN324_data_out(1);
    CN92_sign_in(5) <= VN324_sign_out(1);
    CN92_data_in(6) <= VN378_data_out(1);
    CN92_sign_in(6) <= VN378_sign_out(1);
    CN92_data_in(7) <= VN432_data_out(1);
    CN92_sign_in(7) <= VN432_sign_out(1);
    CN92_data_in(8) <= VN489_data_out(1);
    CN92_sign_in(8) <= VN489_sign_out(1);
    CN92_data_in(9) <= VN516_data_out(1);
    CN92_sign_in(9) <= VN516_sign_out(1);
    CN92_data_in(10) <= VN613_data_out(1);
    CN92_sign_in(10) <= VN613_sign_out(1);
    CN92_data_in(11) <= VN646_data_out(1);
    CN92_sign_in(11) <= VN646_sign_out(1);
    CN92_data_in(12) <= VN718_data_out(1);
    CN92_sign_in(12) <= VN718_sign_out(1);
    CN92_data_in(13) <= VN726_data_out(1);
    CN92_sign_in(13) <= VN726_sign_out(1);
    CN92_data_in(14) <= VN786_data_out(1);
    CN92_sign_in(14) <= VN786_sign_out(1);
    CN92_data_in(15) <= VN831_data_out(1);
    CN92_sign_in(15) <= VN831_sign_out(1);
    CN92_data_in(16) <= VN887_data_out(1);
    CN92_sign_in(16) <= VN887_sign_out(1);
    CN92_data_in(17) <= VN906_data_out(1);
    CN92_sign_in(17) <= VN906_sign_out(1);
    CN92_data_in(18) <= VN984_data_out(1);
    CN92_sign_in(18) <= VN984_sign_out(1);
    CN92_data_in(19) <= VN1030_data_out(1);
    CN92_sign_in(19) <= VN1030_sign_out(1);
    CN92_data_in(20) <= VN1070_data_out(1);
    CN92_sign_in(20) <= VN1070_sign_out(1);
    CN92_data_in(21) <= VN1123_data_out(1);
    CN92_sign_in(21) <= VN1123_sign_out(1);
    CN92_data_in(22) <= VN1191_data_out(1);
    CN92_sign_in(22) <= VN1191_sign_out(1);
    CN92_data_in(23) <= VN1270_data_out(1);
    CN92_sign_in(23) <= VN1270_sign_out(1);
    CN92_data_in(24) <= VN1298_data_out(1);
    CN92_sign_in(24) <= VN1298_sign_out(1);
    CN92_data_in(25) <= VN1369_data_out(1);
    CN92_sign_in(25) <= VN1369_sign_out(1);
    CN92_data_in(26) <= VN1385_data_out(1);
    CN92_sign_in(26) <= VN1385_sign_out(1);
    CN92_data_in(27) <= VN1478_data_out(1);
    CN92_sign_in(27) <= VN1478_sign_out(1);
    CN92_data_in(28) <= VN1613_data_out(1);
    CN92_sign_in(28) <= VN1613_sign_out(1);
    CN92_data_in(29) <= VN1687_data_out(1);
    CN92_sign_in(29) <= VN1687_sign_out(1);
    CN92_data_in(30) <= VN1697_data_out(1);
    CN92_sign_in(30) <= VN1697_sign_out(1);
    CN92_data_in(31) <= VN1744_data_out(1);
    CN92_sign_in(31) <= VN1744_sign_out(1);
    CN93_data_in(0) <= VN25_data_out(1);
    CN93_sign_in(0) <= VN25_sign_out(1);
    CN93_data_in(1) <= VN78_data_out(1);
    CN93_sign_in(1) <= VN78_sign_out(1);
    CN93_data_in(2) <= VN164_data_out(1);
    CN93_sign_in(2) <= VN164_sign_out(1);
    CN93_data_in(3) <= VN224_data_out(1);
    CN93_sign_in(3) <= VN224_sign_out(1);
    CN93_data_in(4) <= VN231_data_out(1);
    CN93_sign_in(4) <= VN231_sign_out(1);
    CN93_data_in(5) <= VN311_data_out(1);
    CN93_sign_in(5) <= VN311_sign_out(1);
    CN93_data_in(6) <= VN340_data_out(1);
    CN93_sign_in(6) <= VN340_sign_out(1);
    CN93_data_in(7) <= VN413_data_out(1);
    CN93_sign_in(7) <= VN413_sign_out(1);
    CN93_data_in(8) <= VN471_data_out(1);
    CN93_sign_in(8) <= VN471_sign_out(1);
    CN93_data_in(9) <= VN545_data_out(1);
    CN93_sign_in(9) <= VN545_sign_out(1);
    CN93_data_in(10) <= VN581_data_out(1);
    CN93_sign_in(10) <= VN581_sign_out(1);
    CN93_data_in(11) <= VN647_data_out(1);
    CN93_sign_in(11) <= VN647_sign_out(1);
    CN93_data_in(12) <= VN698_data_out(1);
    CN93_sign_in(12) <= VN698_sign_out(1);
    CN93_data_in(13) <= VN765_data_out(1);
    CN93_sign_in(13) <= VN765_sign_out(1);
    CN93_data_in(14) <= VN790_data_out(1);
    CN93_sign_in(14) <= VN790_sign_out(1);
    CN93_data_in(15) <= VN848_data_out(1);
    CN93_sign_in(15) <= VN848_sign_out(1);
    CN93_data_in(16) <= VN919_data_out(1);
    CN93_sign_in(16) <= VN919_sign_out(1);
    CN93_data_in(17) <= VN967_data_out(1);
    CN93_sign_in(17) <= VN967_sign_out(1);
    CN93_data_in(18) <= VN1013_data_out(1);
    CN93_sign_in(18) <= VN1013_sign_out(1);
    CN93_data_in(19) <= VN1064_data_out(1);
    CN93_sign_in(19) <= VN1064_sign_out(1);
    CN93_data_in(20) <= VN1138_data_out(1);
    CN93_sign_in(20) <= VN1138_sign_out(1);
    CN93_data_in(21) <= VN1209_data_out(1);
    CN93_sign_in(21) <= VN1209_sign_out(1);
    CN93_data_in(22) <= VN1219_data_out(1);
    CN93_sign_in(22) <= VN1219_sign_out(1);
    CN93_data_in(23) <= VN1266_data_out(1);
    CN93_sign_in(23) <= VN1266_sign_out(1);
    CN93_data_in(24) <= VN1327_data_out(1);
    CN93_sign_in(24) <= VN1327_sign_out(1);
    CN93_data_in(25) <= VN1408_data_out(1);
    CN93_sign_in(25) <= VN1408_sign_out(1);
    CN93_data_in(26) <= VN1456_data_out(1);
    CN93_sign_in(26) <= VN1456_sign_out(1);
    CN93_data_in(27) <= VN1579_data_out(1);
    CN93_sign_in(27) <= VN1579_sign_out(1);
    CN93_data_in(28) <= VN1622_data_out(1);
    CN93_sign_in(28) <= VN1622_sign_out(1);
    CN93_data_in(29) <= VN1661_data_out(1);
    CN93_sign_in(29) <= VN1661_sign_out(1);
    CN93_data_in(30) <= VN1715_data_out(1);
    CN93_sign_in(30) <= VN1715_sign_out(1);
    CN93_data_in(31) <= VN1745_data_out(1);
    CN93_sign_in(31) <= VN1745_sign_out(1);
    CN94_data_in(0) <= VN24_data_out(1);
    CN94_sign_in(0) <= VN24_sign_out(1);
    CN94_data_in(1) <= VN92_data_out(1);
    CN94_sign_in(1) <= VN92_sign_out(1);
    CN94_data_in(2) <= VN194_data_out(1);
    CN94_sign_in(2) <= VN194_sign_out(1);
    CN94_data_in(3) <= VN329_data_out(1);
    CN94_sign_in(3) <= VN329_sign_out(1);
    CN94_data_in(4) <= VN368_data_out(1);
    CN94_sign_in(4) <= VN368_sign_out(1);
    CN94_data_in(5) <= VN421_data_out(1);
    CN94_sign_in(5) <= VN421_sign_out(1);
    CN94_data_in(6) <= VN474_data_out(1);
    CN94_sign_in(6) <= VN474_sign_out(1);
    CN94_data_in(7) <= VN522_data_out(1);
    CN94_sign_in(7) <= VN522_sign_out(1);
    CN94_data_in(8) <= VN579_data_out(1);
    CN94_sign_in(8) <= VN579_sign_out(1);
    CN94_data_in(9) <= VN719_data_out(1);
    CN94_sign_in(9) <= VN719_sign_out(1);
    CN94_data_in(10) <= VN776_data_out(1);
    CN94_sign_in(10) <= VN776_sign_out(1);
    CN94_data_in(11) <= VN780_data_out(1);
    CN94_sign_in(11) <= VN780_sign_out(1);
    CN94_data_in(12) <= VN915_data_out(1);
    CN94_sign_in(12) <= VN915_sign_out(1);
    CN94_data_in(13) <= VN969_data_out(1);
    CN94_sign_in(13) <= VN969_sign_out(1);
    CN94_data_in(14) <= VN1024_data_out(1);
    CN94_sign_in(14) <= VN1024_sign_out(1);
    CN94_data_in(15) <= VN1068_data_out(1);
    CN94_sign_in(15) <= VN1068_sign_out(1);
    CN94_data_in(16) <= VN1164_data_out(1);
    CN94_sign_in(16) <= VN1164_sign_out(1);
    CN94_data_in(17) <= VN1175_data_out(1);
    CN94_sign_in(17) <= VN1175_sign_out(1);
    CN94_data_in(18) <= VN1230_data_out(1);
    CN94_sign_in(18) <= VN1230_sign_out(1);
    CN94_data_in(19) <= VN1375_data_out(1);
    CN94_sign_in(19) <= VN1375_sign_out(1);
    CN94_data_in(20) <= VN1412_data_out(1);
    CN94_sign_in(20) <= VN1412_sign_out(1);
    CN94_data_in(21) <= VN1467_data_out(1);
    CN94_sign_in(21) <= VN1467_sign_out(1);
    CN94_data_in(22) <= VN1482_data_out(1);
    CN94_sign_in(22) <= VN1482_sign_out(1);
    CN94_data_in(23) <= VN1617_data_out(1);
    CN94_sign_in(23) <= VN1617_sign_out(1);
    CN94_data_in(24) <= VN1656_data_out(1);
    CN94_sign_in(24) <= VN1656_sign_out(1);
    CN94_data_in(25) <= VN1805_data_out(1);
    CN94_sign_in(25) <= VN1805_sign_out(1);
    CN94_data_in(26) <= VN1887_data_out(1);
    CN94_sign_in(26) <= VN1887_sign_out(1);
    CN94_data_in(27) <= VN1895_data_out(1);
    CN94_sign_in(27) <= VN1895_sign_out(1);
    CN94_data_in(28) <= VN1901_data_out(1);
    CN94_sign_in(28) <= VN1901_sign_out(1);
    CN94_data_in(29) <= VN1933_data_out(1);
    CN94_sign_in(29) <= VN1933_sign_out(1);
    CN94_data_in(30) <= VN1936_data_out(1);
    CN94_sign_in(30) <= VN1936_sign_out(1);
    CN94_data_in(31) <= VN1943_data_out(1);
    CN94_sign_in(31) <= VN1943_sign_out(1);
    CN95_data_in(0) <= VN23_data_out(1);
    CN95_sign_in(0) <= VN23_sign_out(1);
    CN95_data_in(1) <= VN63_data_out(1);
    CN95_sign_in(1) <= VN63_sign_out(1);
    CN95_data_in(2) <= VN134_data_out(1);
    CN95_sign_in(2) <= VN134_sign_out(1);
    CN95_data_in(3) <= VN190_data_out(1);
    CN95_sign_in(3) <= VN190_sign_out(1);
    CN95_data_in(4) <= VN234_data_out(1);
    CN95_sign_in(4) <= VN234_sign_out(1);
    CN95_data_in(5) <= VN303_data_out(1);
    CN95_sign_in(5) <= VN303_sign_out(1);
    CN95_data_in(6) <= VN352_data_out(1);
    CN95_sign_in(6) <= VN352_sign_out(1);
    CN95_data_in(7) <= VN443_data_out(1);
    CN95_sign_in(7) <= VN443_sign_out(1);
    CN95_data_in(8) <= VN460_data_out(1);
    CN95_sign_in(8) <= VN460_sign_out(1);
    CN95_data_in(9) <= VN547_data_out(1);
    CN95_sign_in(9) <= VN547_sign_out(1);
    CN95_data_in(10) <= VN611_data_out(1);
    CN95_sign_in(10) <= VN611_sign_out(1);
    CN95_data_in(11) <= VN618_data_out(1);
    CN95_sign_in(11) <= VN618_sign_out(1);
    CN95_data_in(12) <= VN678_data_out(1);
    CN95_sign_in(12) <= VN678_sign_out(1);
    CN95_data_in(13) <= VN732_data_out(1);
    CN95_sign_in(13) <= VN732_sign_out(1);
    CN95_data_in(14) <= VN814_data_out(1);
    CN95_sign_in(14) <= VN814_sign_out(1);
    CN95_data_in(15) <= VN875_data_out(1);
    CN95_sign_in(15) <= VN875_sign_out(1);
    CN95_data_in(16) <= VN932_data_out(1);
    CN95_sign_in(16) <= VN932_sign_out(1);
    CN95_data_in(17) <= VN995_data_out(1);
    CN95_sign_in(17) <= VN995_sign_out(1);
    CN95_data_in(18) <= VN1031_data_out(1);
    CN95_sign_in(18) <= VN1031_sign_out(1);
    CN95_data_in(19) <= VN1145_data_out(1);
    CN95_sign_in(19) <= VN1145_sign_out(1);
    CN95_data_in(20) <= VN1176_data_out(1);
    CN95_sign_in(20) <= VN1176_sign_out(1);
    CN95_data_in(21) <= VN1250_data_out(1);
    CN95_sign_in(21) <= VN1250_sign_out(1);
    CN95_data_in(22) <= VN1444_data_out(1);
    CN95_sign_in(22) <= VN1444_sign_out(1);
    CN95_data_in(23) <= VN1487_data_out(1);
    CN95_sign_in(23) <= VN1487_sign_out(1);
    CN95_data_in(24) <= VN1507_data_out(1);
    CN95_sign_in(24) <= VN1507_sign_out(1);
    CN95_data_in(25) <= VN1528_data_out(1);
    CN95_sign_in(25) <= VN1528_sign_out(1);
    CN95_data_in(26) <= VN1535_data_out(1);
    CN95_sign_in(26) <= VN1535_sign_out(1);
    CN95_data_in(27) <= VN1552_data_out(1);
    CN95_sign_in(27) <= VN1552_sign_out(1);
    CN95_data_in(28) <= VN1566_data_out(1);
    CN95_sign_in(28) <= VN1566_sign_out(1);
    CN95_data_in(29) <= VN1623_data_out(1);
    CN95_sign_in(29) <= VN1623_sign_out(1);
    CN95_data_in(30) <= VN1684_data_out(1);
    CN95_sign_in(30) <= VN1684_sign_out(1);
    CN95_data_in(31) <= VN1746_data_out(1);
    CN95_sign_in(31) <= VN1746_sign_out(1);
    CN96_data_in(0) <= VN22_data_out(1);
    CN96_sign_in(0) <= VN22_sign_out(1);
    CN96_data_in(1) <= VN98_data_out(1);
    CN96_sign_in(1) <= VN98_sign_out(1);
    CN96_data_in(2) <= VN150_data_out(1);
    CN96_sign_in(2) <= VN150_sign_out(1);
    CN96_data_in(3) <= VN172_data_out(1);
    CN96_sign_in(3) <= VN172_sign_out(1);
    CN96_data_in(4) <= VN251_data_out(1);
    CN96_sign_in(4) <= VN251_sign_out(1);
    CN96_data_in(5) <= VN380_data_out(1);
    CN96_sign_in(5) <= VN380_sign_out(1);
    CN96_data_in(6) <= VN441_data_out(1);
    CN96_sign_in(6) <= VN441_sign_out(1);
    CN96_data_in(7) <= VN490_data_out(1);
    CN96_sign_in(7) <= VN490_sign_out(1);
    CN96_data_in(8) <= VN560_data_out(1);
    CN96_sign_in(8) <= VN560_sign_out(1);
    CN96_data_in(9) <= VN592_data_out(1);
    CN96_sign_in(9) <= VN592_sign_out(1);
    CN96_data_in(10) <= VN631_data_out(1);
    CN96_sign_in(10) <= VN631_sign_out(1);
    CN96_data_in(11) <= VN675_data_out(1);
    CN96_sign_in(11) <= VN675_sign_out(1);
    CN96_data_in(12) <= VN760_data_out(1);
    CN96_sign_in(12) <= VN760_sign_out(1);
    CN96_data_in(13) <= VN798_data_out(1);
    CN96_sign_in(13) <= VN798_sign_out(1);
    CN96_data_in(14) <= VN870_data_out(1);
    CN96_sign_in(14) <= VN870_sign_out(1);
    CN96_data_in(15) <= VN899_data_out(1);
    CN96_sign_in(15) <= VN899_sign_out(1);
    CN96_data_in(16) <= VN976_data_out(1);
    CN96_sign_in(16) <= VN976_sign_out(1);
    CN96_data_in(17) <= VN1006_data_out(1);
    CN96_sign_in(17) <= VN1006_sign_out(1);
    CN96_data_in(18) <= VN1090_data_out(1);
    CN96_sign_in(18) <= VN1090_sign_out(1);
    CN96_data_in(19) <= VN1208_data_out(1);
    CN96_sign_in(19) <= VN1208_sign_out(1);
    CN96_data_in(20) <= VN1251_data_out(1);
    CN96_sign_in(20) <= VN1251_sign_out(1);
    CN96_data_in(21) <= VN1283_data_out(1);
    CN96_sign_in(21) <= VN1283_sign_out(1);
    CN96_data_in(22) <= VN1338_data_out(1);
    CN96_sign_in(22) <= VN1338_sign_out(1);
    CN96_data_in(23) <= VN1453_data_out(1);
    CN96_sign_in(23) <= VN1453_sign_out(1);
    CN96_data_in(24) <= VN1476_data_out(1);
    CN96_sign_in(24) <= VN1476_sign_out(1);
    CN96_data_in(25) <= VN1513_data_out(1);
    CN96_sign_in(25) <= VN1513_sign_out(1);
    CN96_data_in(26) <= VN1571_data_out(1);
    CN96_sign_in(26) <= VN1571_sign_out(1);
    CN96_data_in(27) <= VN1612_data_out(1);
    CN96_sign_in(27) <= VN1612_sign_out(1);
    CN96_data_in(28) <= VN1689_data_out(1);
    CN96_sign_in(28) <= VN1689_sign_out(1);
    CN96_data_in(29) <= VN1735_data_out(1);
    CN96_sign_in(29) <= VN1735_sign_out(1);
    CN96_data_in(30) <= VN1886_data_out(1);
    CN96_sign_in(30) <= VN1886_sign_out(1);
    CN96_data_in(31) <= VN1908_data_out(1);
    CN96_sign_in(31) <= VN1908_sign_out(1);
    CN97_data_in(0) <= VN21_data_out(1);
    CN97_sign_in(0) <= VN21_sign_out(1);
    CN97_data_in(1) <= VN65_data_out(1);
    CN97_sign_in(1) <= VN65_sign_out(1);
    CN97_data_in(2) <= VN142_data_out(1);
    CN97_sign_in(2) <= VN142_sign_out(1);
    CN97_data_in(3) <= VN180_data_out(1);
    CN97_sign_in(3) <= VN180_sign_out(1);
    CN97_data_in(4) <= VN260_data_out(1);
    CN97_sign_in(4) <= VN260_sign_out(1);
    CN97_data_in(5) <= VN316_data_out(1);
    CN97_sign_in(5) <= VN316_sign_out(1);
    CN97_data_in(6) <= VN370_data_out(1);
    CN97_sign_in(6) <= VN370_sign_out(1);
    CN97_data_in(7) <= VN419_data_out(1);
    CN97_sign_in(7) <= VN419_sign_out(1);
    CN97_data_in(8) <= VN456_data_out(1);
    CN97_sign_in(8) <= VN456_sign_out(1);
    CN97_data_in(9) <= VN557_data_out(1);
    CN97_sign_in(9) <= VN557_sign_out(1);
    CN97_data_in(10) <= VN595_data_out(1);
    CN97_sign_in(10) <= VN595_sign_out(1);
    CN97_data_in(11) <= VN636_data_out(1);
    CN97_sign_in(11) <= VN636_sign_out(1);
    CN97_data_in(12) <= VN693_data_out(1);
    CN97_sign_in(12) <= VN693_sign_out(1);
    CN97_data_in(13) <= VN748_data_out(1);
    CN97_sign_in(13) <= VN748_sign_out(1);
    CN97_data_in(14) <= VN809_data_out(1);
    CN97_sign_in(14) <= VN809_sign_out(1);
    CN97_data_in(15) <= VN876_data_out(1);
    CN97_sign_in(15) <= VN876_sign_out(1);
    CN97_data_in(16) <= VN900_data_out(1);
    CN97_sign_in(16) <= VN900_sign_out(1);
    CN97_data_in(17) <= VN988_data_out(1);
    CN97_sign_in(17) <= VN988_sign_out(1);
    CN97_data_in(18) <= VN1020_data_out(1);
    CN97_sign_in(18) <= VN1020_sign_out(1);
    CN97_data_in(19) <= VN1077_data_out(1);
    CN97_sign_in(19) <= VN1077_sign_out(1);
    CN97_data_in(20) <= VN1125_data_out(1);
    CN97_sign_in(20) <= VN1125_sign_out(1);
    CN97_data_in(21) <= VN1199_data_out(1);
    CN97_sign_in(21) <= VN1199_sign_out(1);
    CN97_data_in(22) <= VN1229_data_out(1);
    CN97_sign_in(22) <= VN1229_sign_out(1);
    CN97_data_in(23) <= VN1324_data_out(1);
    CN97_sign_in(23) <= VN1324_sign_out(1);
    CN97_data_in(24) <= VN1368_data_out(1);
    CN97_sign_in(24) <= VN1368_sign_out(1);
    CN97_data_in(25) <= VN1406_data_out(1);
    CN97_sign_in(25) <= VN1406_sign_out(1);
    CN97_data_in(26) <= VN1447_data_out(1);
    CN97_sign_in(26) <= VN1447_sign_out(1);
    CN97_data_in(27) <= VN1575_data_out(1);
    CN97_sign_in(27) <= VN1575_sign_out(1);
    CN97_data_in(28) <= VN1596_data_out(1);
    CN97_sign_in(28) <= VN1596_sign_out(1);
    CN97_data_in(29) <= VN1633_data_out(1);
    CN97_sign_in(29) <= VN1633_sign_out(1);
    CN97_data_in(30) <= VN1665_data_out(1);
    CN97_sign_in(30) <= VN1665_sign_out(1);
    CN97_data_in(31) <= VN1747_data_out(1);
    CN97_sign_in(31) <= VN1747_sign_out(1);
    CN98_data_in(0) <= VN20_data_out(1);
    CN98_sign_in(0) <= VN20_sign_out(1);
    CN98_data_in(1) <= VN116_data_out(1);
    CN98_sign_in(1) <= VN116_sign_out(1);
    CN98_data_in(2) <= VN199_data_out(1);
    CN98_sign_in(2) <= VN199_sign_out(1);
    CN98_data_in(3) <= VN255_data_out(1);
    CN98_sign_in(3) <= VN255_sign_out(1);
    CN98_data_in(4) <= VN308_data_out(1);
    CN98_sign_in(4) <= VN308_sign_out(1);
    CN98_data_in(5) <= VN356_data_out(1);
    CN98_sign_in(5) <= VN356_sign_out(1);
    CN98_data_in(6) <= VN400_data_out(1);
    CN98_sign_in(6) <= VN400_sign_out(1);
    CN98_data_in(7) <= VN482_data_out(1);
    CN98_sign_in(7) <= VN482_sign_out(1);
    CN98_data_in(8) <= VN518_data_out(1);
    CN98_sign_in(8) <= VN518_sign_out(1);
    CN98_data_in(9) <= VN582_data_out(1);
    CN98_sign_in(9) <= VN582_sign_out(1);
    CN98_data_in(10) <= VN668_data_out(1);
    CN98_sign_in(10) <= VN668_sign_out(1);
    CN98_data_in(11) <= VN714_data_out(1);
    CN98_sign_in(11) <= VN714_sign_out(1);
    CN98_data_in(12) <= VN735_data_out(1);
    CN98_sign_in(12) <= VN735_sign_out(1);
    CN98_data_in(13) <= VN820_data_out(1);
    CN98_sign_in(13) <= VN820_sign_out(1);
    CN98_data_in(14) <= VN866_data_out(1);
    CN98_sign_in(14) <= VN866_sign_out(1);
    CN98_data_in(15) <= VN931_data_out(1);
    CN98_sign_in(15) <= VN931_sign_out(1);
    CN98_data_in(16) <= VN996_data_out(1);
    CN98_sign_in(16) <= VN996_sign_out(1);
    CN98_data_in(17) <= VN1048_data_out(1);
    CN98_sign_in(17) <= VN1048_sign_out(1);
    CN98_data_in(18) <= VN1215_data_out(1);
    CN98_sign_in(18) <= VN1215_sign_out(1);
    CN98_data_in(19) <= VN1382_data_out(1);
    CN98_sign_in(19) <= VN1382_sign_out(1);
    CN98_data_in(20) <= VN1450_data_out(1);
    CN98_sign_in(20) <= VN1450_sign_out(1);
    CN98_data_in(21) <= VN1520_data_out(1);
    CN98_sign_in(21) <= VN1520_sign_out(1);
    CN98_data_in(22) <= VN1551_data_out(1);
    CN98_sign_in(22) <= VN1551_sign_out(1);
    CN98_data_in(23) <= VN1570_data_out(1);
    CN98_sign_in(23) <= VN1570_sign_out(1);
    CN98_data_in(24) <= VN1584_data_out(1);
    CN98_sign_in(24) <= VN1584_sign_out(1);
    CN98_data_in(25) <= VN1638_data_out(1);
    CN98_sign_in(25) <= VN1638_sign_out(1);
    CN98_data_in(26) <= VN1699_data_out(1);
    CN98_sign_in(26) <= VN1699_sign_out(1);
    CN98_data_in(27) <= VN1781_data_out(1);
    CN98_sign_in(27) <= VN1781_sign_out(1);
    CN98_data_in(28) <= VN1818_data_out(1);
    CN98_sign_in(28) <= VN1818_sign_out(1);
    CN98_data_in(29) <= VN1968_data_out(1);
    CN98_sign_in(29) <= VN1968_sign_out(1);
    CN98_data_in(30) <= VN2036_data_out(1);
    CN98_sign_in(30) <= VN2036_sign_out(1);
    CN98_data_in(31) <= VN2041_data_out(1);
    CN98_sign_in(31) <= VN2041_sign_out(1);
    CN99_data_in(0) <= VN19_data_out(1);
    CN99_sign_in(0) <= VN19_sign_out(1);
    CN99_data_in(1) <= VN76_data_out(1);
    CN99_sign_in(1) <= VN76_sign_out(1);
    CN99_data_in(2) <= VN126_data_out(1);
    CN99_sign_in(2) <= VN126_sign_out(1);
    CN99_data_in(3) <= VN198_data_out(1);
    CN99_sign_in(3) <= VN198_sign_out(1);
    CN99_data_in(4) <= VN261_data_out(1);
    CN99_sign_in(4) <= VN261_sign_out(1);
    CN99_data_in(5) <= VN285_data_out(1);
    CN99_sign_in(5) <= VN285_sign_out(1);
    CN99_data_in(6) <= VN376_data_out(1);
    CN99_sign_in(6) <= VN376_sign_out(1);
    CN99_data_in(7) <= VN402_data_out(1);
    CN99_sign_in(7) <= VN402_sign_out(1);
    CN99_data_in(8) <= VN467_data_out(1);
    CN99_sign_in(8) <= VN467_sign_out(1);
    CN99_data_in(9) <= VN540_data_out(1);
    CN99_sign_in(9) <= VN540_sign_out(1);
    CN99_data_in(10) <= VN612_data_out(1);
    CN99_sign_in(10) <= VN612_sign_out(1);
    CN99_data_in(11) <= VN635_data_out(1);
    CN99_sign_in(11) <= VN635_sign_out(1);
    CN99_data_in(12) <= VN715_data_out(1);
    CN99_sign_in(12) <= VN715_sign_out(1);
    CN99_data_in(13) <= VN750_data_out(1);
    CN99_sign_in(13) <= VN750_sign_out(1);
    CN99_data_in(14) <= VN793_data_out(1);
    CN99_sign_in(14) <= VN793_sign_out(1);
    CN99_data_in(15) <= VN834_data_out(1);
    CN99_sign_in(15) <= VN834_sign_out(1);
    CN99_data_in(16) <= VN925_data_out(1);
    CN99_sign_in(16) <= VN925_sign_out(1);
    CN99_data_in(17) <= VN968_data_out(1);
    CN99_sign_in(17) <= VN968_sign_out(1);
    CN99_data_in(18) <= VN1026_data_out(1);
    CN99_sign_in(18) <= VN1026_sign_out(1);
    CN99_data_in(19) <= VN1096_data_out(1);
    CN99_sign_in(19) <= VN1096_sign_out(1);
    CN99_data_in(20) <= VN1140_data_out(1);
    CN99_sign_in(20) <= VN1140_sign_out(1);
    CN99_data_in(21) <= VN1238_data_out(1);
    CN99_sign_in(21) <= VN1238_sign_out(1);
    CN99_data_in(22) <= VN1290_data_out(1);
    CN99_sign_in(22) <= VN1290_sign_out(1);
    CN99_data_in(23) <= VN1355_data_out(1);
    CN99_sign_in(23) <= VN1355_sign_out(1);
    CN99_data_in(24) <= VN1395_data_out(1);
    CN99_sign_in(24) <= VN1395_sign_out(1);
    CN99_data_in(25) <= VN1558_data_out(1);
    CN99_sign_in(25) <= VN1558_sign_out(1);
    CN99_data_in(26) <= VN1564_data_out(1);
    CN99_sign_in(26) <= VN1564_sign_out(1);
    CN99_data_in(27) <= VN1592_data_out(1);
    CN99_sign_in(27) <= VN1592_sign_out(1);
    CN99_data_in(28) <= VN1626_data_out(1);
    CN99_sign_in(28) <= VN1626_sign_out(1);
    CN99_data_in(29) <= VN1649_data_out(1);
    CN99_sign_in(29) <= VN1649_sign_out(1);
    CN99_data_in(30) <= VN1691_data_out(1);
    CN99_sign_in(30) <= VN1691_sign_out(1);
    CN99_data_in(31) <= VN1748_data_out(1);
    CN99_sign_in(31) <= VN1748_sign_out(1);
    CN100_data_in(0) <= VN18_data_out(1);
    CN100_sign_in(0) <= VN18_sign_out(1);
    CN100_data_in(1) <= VN94_data_out(1);
    CN100_sign_in(1) <= VN94_sign_out(1);
    CN100_data_in(2) <= VN120_data_out(1);
    CN100_sign_in(2) <= VN120_sign_out(1);
    CN100_data_in(3) <= VN178_data_out(1);
    CN100_sign_in(3) <= VN178_sign_out(1);
    CN100_data_in(4) <= VN250_data_out(1);
    CN100_sign_in(4) <= VN250_sign_out(1);
    CN100_data_in(5) <= VN295_data_out(1);
    CN100_sign_in(5) <= VN295_sign_out(1);
    CN100_data_in(6) <= VN349_data_out(1);
    CN100_sign_in(6) <= VN349_sign_out(1);
    CN100_data_in(7) <= VN444_data_out(1);
    CN100_sign_in(7) <= VN444_sign_out(1);
    CN100_data_in(8) <= VN492_data_out(1);
    CN100_sign_in(8) <= VN492_sign_out(1);
    CN100_data_in(9) <= VN541_data_out(1);
    CN100_sign_in(9) <= VN541_sign_out(1);
    CN100_data_in(10) <= VN578_data_out(1);
    CN100_sign_in(10) <= VN578_sign_out(1);
    CN100_data_in(11) <= VN692_data_out(1);
    CN100_sign_in(11) <= VN692_sign_out(1);
    CN100_data_in(12) <= VN770_data_out(1);
    CN100_sign_in(12) <= VN770_sign_out(1);
    CN100_data_in(13) <= VN782_data_out(1);
    CN100_sign_in(13) <= VN782_sign_out(1);
    CN100_data_in(14) <= VN840_data_out(1);
    CN100_sign_in(14) <= VN840_sign_out(1);
    CN100_data_in(15) <= VN941_data_out(1);
    CN100_sign_in(15) <= VN941_sign_out(1);
    CN100_data_in(16) <= VN983_data_out(1);
    CN100_sign_in(16) <= VN983_sign_out(1);
    CN100_data_in(17) <= VN1050_data_out(1);
    CN100_sign_in(17) <= VN1050_sign_out(1);
    CN100_data_in(18) <= VN1071_data_out(1);
    CN100_sign_in(18) <= VN1071_sign_out(1);
    CN100_data_in(19) <= VN1163_data_out(1);
    CN100_sign_in(19) <= VN1163_sign_out(1);
    CN100_data_in(20) <= VN1220_data_out(1);
    CN100_sign_in(20) <= VN1220_sign_out(1);
    CN100_data_in(21) <= VN1241_data_out(1);
    CN100_sign_in(21) <= VN1241_sign_out(1);
    CN100_data_in(22) <= VN1301_data_out(1);
    CN100_sign_in(22) <= VN1301_sign_out(1);
    CN100_data_in(23) <= VN1335_data_out(1);
    CN100_sign_in(23) <= VN1335_sign_out(1);
    CN100_data_in(24) <= VN1417_data_out(1);
    CN100_sign_in(24) <= VN1417_sign_out(1);
    CN100_data_in(25) <= VN1441_data_out(1);
    CN100_sign_in(25) <= VN1441_sign_out(1);
    CN100_data_in(26) <= VN1519_data_out(1);
    CN100_sign_in(26) <= VN1519_sign_out(1);
    CN100_data_in(27) <= VN1602_data_out(1);
    CN100_sign_in(27) <= VN1602_sign_out(1);
    CN100_data_in(28) <= VN1627_data_out(1);
    CN100_sign_in(28) <= VN1627_sign_out(1);
    CN100_data_in(29) <= VN1671_data_out(1);
    CN100_sign_in(29) <= VN1671_sign_out(1);
    CN100_data_in(30) <= VN1778_data_out(1);
    CN100_sign_in(30) <= VN1778_sign_out(1);
    CN100_data_in(31) <= VN1825_data_out(1);
    CN100_sign_in(31) <= VN1825_sign_out(1);
    CN101_data_in(0) <= VN17_data_out(1);
    CN101_sign_in(0) <= VN17_sign_out(1);
    CN101_data_in(1) <= VN58_data_out(1);
    CN101_sign_in(1) <= VN58_sign_out(1);
    CN101_data_in(2) <= VN123_data_out(1);
    CN101_sign_in(2) <= VN123_sign_out(1);
    CN101_data_in(3) <= VN211_data_out(1);
    CN101_sign_in(3) <= VN211_sign_out(1);
    CN101_data_in(4) <= VN273_data_out(1);
    CN101_sign_in(4) <= VN273_sign_out(1);
    CN101_data_in(5) <= VN289_data_out(1);
    CN101_sign_in(5) <= VN289_sign_out(1);
    CN101_data_in(6) <= VN346_data_out(1);
    CN101_sign_in(6) <= VN346_sign_out(1);
    CN101_data_in(7) <= VN420_data_out(1);
    CN101_sign_in(7) <= VN420_sign_out(1);
    CN101_data_in(8) <= VN517_data_out(1);
    CN101_sign_in(8) <= VN517_sign_out(1);
    CN101_data_in(9) <= VN603_data_out(1);
    CN101_sign_in(9) <= VN603_sign_out(1);
    CN101_data_in(10) <= VN684_data_out(1);
    CN101_sign_in(10) <= VN684_sign_out(1);
    CN101_data_in(11) <= VN724_data_out(1);
    CN101_sign_in(11) <= VN724_sign_out(1);
    CN101_data_in(12) <= VN823_data_out(1);
    CN101_sign_in(12) <= VN823_sign_out(1);
    CN101_data_in(13) <= VN830_data_out(1);
    CN101_sign_in(13) <= VN830_sign_out(1);
    CN101_data_in(14) <= VN879_data_out(1);
    CN101_sign_in(14) <= VN879_sign_out(1);
    CN101_data_in(15) <= VN889_data_out(1);
    CN101_sign_in(15) <= VN889_sign_out(1);
    CN101_data_in(16) <= VN954_data_out(1);
    CN101_sign_in(16) <= VN954_sign_out(1);
    CN101_data_in(17) <= VN1357_data_out(1);
    CN101_sign_in(17) <= VN1357_sign_out(1);
    CN101_data_in(18) <= VN1472_data_out(1);
    CN101_sign_in(18) <= VN1472_sign_out(1);
    CN101_data_in(19) <= VN1488_data_out(1);
    CN101_sign_in(19) <= VN1488_sign_out(1);
    CN101_data_in(20) <= VN1508_data_out(1);
    CN101_sign_in(20) <= VN1508_sign_out(1);
    CN101_data_in(21) <= VN1516_data_out(1);
    CN101_sign_in(21) <= VN1516_sign_out(1);
    CN101_data_in(22) <= VN1525_data_out(1);
    CN101_sign_in(22) <= VN1525_sign_out(1);
    CN101_data_in(23) <= VN1674_data_out(1);
    CN101_sign_in(23) <= VN1674_sign_out(1);
    CN101_data_in(24) <= VN1710_data_out(1);
    CN101_sign_in(24) <= VN1710_sign_out(1);
    CN101_data_in(25) <= VN1831_data_out(1);
    CN101_sign_in(25) <= VN1831_sign_out(1);
    CN101_data_in(26) <= VN1840_data_out(1);
    CN101_sign_in(26) <= VN1840_sign_out(1);
    CN101_data_in(27) <= VN1850_data_out(1);
    CN101_sign_in(27) <= VN1850_sign_out(1);
    CN101_data_in(28) <= VN1884_data_out(1);
    CN101_sign_in(28) <= VN1884_sign_out(1);
    CN101_data_in(29) <= VN1912_data_out(1);
    CN101_sign_in(29) <= VN1912_sign_out(1);
    CN101_data_in(30) <= VN1997_data_out(1);
    CN101_sign_in(30) <= VN1997_sign_out(1);
    CN101_data_in(31) <= VN2002_data_out(1);
    CN101_sign_in(31) <= VN2002_sign_out(1);
    CN102_data_in(0) <= VN16_data_out(1);
    CN102_sign_in(0) <= VN16_sign_out(1);
    CN102_data_in(1) <= VN59_data_out(1);
    CN102_sign_in(1) <= VN59_sign_out(1);
    CN102_data_in(2) <= VN113_data_out(1);
    CN102_sign_in(2) <= VN113_sign_out(1);
    CN102_data_in(3) <= VN214_data_out(1);
    CN102_sign_in(3) <= VN214_sign_out(1);
    CN102_data_in(4) <= VN226_data_out(1);
    CN102_sign_in(4) <= VN226_sign_out(1);
    CN102_data_in(5) <= VN361_data_out(1);
    CN102_sign_in(5) <= VN361_sign_out(1);
    CN102_data_in(6) <= VN440_data_out(1);
    CN102_sign_in(6) <= VN440_sign_out(1);
    CN102_data_in(7) <= VN472_data_out(1);
    CN102_sign_in(7) <= VN472_sign_out(1);
    CN102_data_in(8) <= VN510_data_out(1);
    CN102_sign_in(8) <= VN510_sign_out(1);
    CN102_data_in(9) <= VN589_data_out(1);
    CN102_sign_in(9) <= VN589_sign_out(1);
    CN102_data_in(10) <= VN621_data_out(1);
    CN102_sign_in(10) <= VN621_sign_out(1);
    CN102_data_in(11) <= VN702_data_out(1);
    CN102_sign_in(11) <= VN702_sign_out(1);
    CN102_data_in(12) <= VN774_data_out(1);
    CN102_sign_in(12) <= VN774_sign_out(1);
    CN102_data_in(13) <= VN881_data_out(1);
    CN102_sign_in(13) <= VN881_sign_out(1);
    CN102_data_in(14) <= VN991_data_out(1);
    CN102_sign_in(14) <= VN991_sign_out(1);
    CN102_data_in(15) <= VN1005_data_out(1);
    CN102_sign_in(15) <= VN1005_sign_out(1);
    CN102_data_in(16) <= VN1098_data_out(1);
    CN102_sign_in(16) <= VN1098_sign_out(1);
    CN102_data_in(17) <= VN1139_data_out(1);
    CN102_sign_in(17) <= VN1139_sign_out(1);
    CN102_data_in(18) <= VN1285_data_out(1);
    CN102_sign_in(18) <= VN1285_sign_out(1);
    CN102_data_in(19) <= VN1477_data_out(1);
    CN102_sign_in(19) <= VN1477_sign_out(1);
    CN102_data_in(20) <= VN1502_data_out(1);
    CN102_sign_in(20) <= VN1502_sign_out(1);
    CN102_data_in(21) <= VN1631_data_out(1);
    CN102_sign_in(21) <= VN1631_sign_out(1);
    CN102_data_in(22) <= VN1666_data_out(1);
    CN102_sign_in(22) <= VN1666_sign_out(1);
    CN102_data_in(23) <= VN1713_data_out(1);
    CN102_sign_in(23) <= VN1713_sign_out(1);
    CN102_data_in(24) <= VN1798_data_out(1);
    CN102_sign_in(24) <= VN1798_sign_out(1);
    CN102_data_in(25) <= VN1844_data_out(1);
    CN102_sign_in(25) <= VN1844_sign_out(1);
    CN102_data_in(26) <= VN1890_data_out(1);
    CN102_sign_in(26) <= VN1890_sign_out(1);
    CN102_data_in(27) <= VN1906_data_out(1);
    CN102_sign_in(27) <= VN1906_sign_out(1);
    CN102_data_in(28) <= VN1989_data_out(1);
    CN102_sign_in(28) <= VN1989_sign_out(1);
    CN102_data_in(29) <= VN2004_data_out(1);
    CN102_sign_in(29) <= VN2004_sign_out(1);
    CN102_data_in(30) <= VN2023_data_out(1);
    CN102_sign_in(30) <= VN2023_sign_out(1);
    CN102_data_in(31) <= VN2027_data_out(1);
    CN102_sign_in(31) <= VN2027_sign_out(1);
    CN103_data_in(0) <= VN15_data_out(1);
    CN103_sign_in(0) <= VN15_sign_out(1);
    CN103_data_in(1) <= VN93_data_out(1);
    CN103_sign_in(1) <= VN93_sign_out(1);
    CN103_data_in(2) <= VN151_data_out(1);
    CN103_sign_in(2) <= VN151_sign_out(1);
    CN103_data_in(3) <= VN200_data_out(1);
    CN103_sign_in(3) <= VN200_sign_out(1);
    CN103_data_in(4) <= VN265_data_out(1);
    CN103_sign_in(4) <= VN265_sign_out(1);
    CN103_data_in(5) <= VN284_data_out(1);
    CN103_sign_in(5) <= VN284_sign_out(1);
    CN103_data_in(6) <= VN354_data_out(1);
    CN103_sign_in(6) <= VN354_sign_out(1);
    CN103_data_in(7) <= VN410_data_out(1);
    CN103_sign_in(7) <= VN410_sign_out(1);
    CN103_data_in(8) <= VN488_data_out(1);
    CN103_sign_in(8) <= VN488_sign_out(1);
    CN103_data_in(9) <= VN525_data_out(1);
    CN103_sign_in(9) <= VN525_sign_out(1);
    CN103_data_in(10) <= VN614_data_out(1);
    CN103_sign_in(10) <= VN614_sign_out(1);
    CN103_data_in(11) <= VN642_data_out(1);
    CN103_sign_in(11) <= VN642_sign_out(1);
    CN103_data_in(12) <= VN706_data_out(1);
    CN103_sign_in(12) <= VN706_sign_out(1);
    CN103_data_in(13) <= VN802_data_out(1);
    CN103_sign_in(13) <= VN802_sign_out(1);
    CN103_data_in(14) <= VN852_data_out(1);
    CN103_sign_in(14) <= VN852_sign_out(1);
    CN103_data_in(15) <= VN888_data_out(1);
    CN103_sign_in(15) <= VN888_sign_out(1);
    CN103_data_in(16) <= VN956_data_out(1);
    CN103_sign_in(16) <= VN956_sign_out(1);
    CN103_data_in(17) <= VN1022_data_out(1);
    CN103_sign_in(17) <= VN1022_sign_out(1);
    CN103_data_in(18) <= VN1062_data_out(1);
    CN103_sign_in(18) <= VN1062_sign_out(1);
    CN103_data_in(19) <= VN1131_data_out(1);
    CN103_sign_in(19) <= VN1131_sign_out(1);
    CN103_data_in(20) <= VN1197_data_out(1);
    CN103_sign_in(20) <= VN1197_sign_out(1);
    CN103_data_in(21) <= VN1236_data_out(1);
    CN103_sign_in(21) <= VN1236_sign_out(1);
    CN103_data_in(22) <= VN1326_data_out(1);
    CN103_sign_in(22) <= VN1326_sign_out(1);
    CN103_data_in(23) <= VN1366_data_out(1);
    CN103_sign_in(23) <= VN1366_sign_out(1);
    CN103_data_in(24) <= VN1538_data_out(1);
    CN103_sign_in(24) <= VN1538_sign_out(1);
    CN103_data_in(25) <= VN1553_data_out(1);
    CN103_sign_in(25) <= VN1553_sign_out(1);
    CN103_data_in(26) <= VN1573_data_out(1);
    CN103_sign_in(26) <= VN1573_sign_out(1);
    CN103_data_in(27) <= VN1604_data_out(1);
    CN103_sign_in(27) <= VN1604_sign_out(1);
    CN103_data_in(28) <= VN1642_data_out(1);
    CN103_sign_in(28) <= VN1642_sign_out(1);
    CN103_data_in(29) <= VN1650_data_out(1);
    CN103_sign_in(29) <= VN1650_sign_out(1);
    CN103_data_in(30) <= VN1712_data_out(1);
    CN103_sign_in(30) <= VN1712_sign_out(1);
    CN103_data_in(31) <= VN1749_data_out(1);
    CN103_sign_in(31) <= VN1749_sign_out(1);
    CN104_data_in(0) <= VN14_data_out(1);
    CN104_sign_in(0) <= VN14_sign_out(1);
    CN104_data_in(1) <= VN86_data_out(1);
    CN104_sign_in(1) <= VN86_sign_out(1);
    CN104_data_in(2) <= VN133_data_out(1);
    CN104_sign_in(2) <= VN133_sign_out(1);
    CN104_data_in(3) <= VN179_data_out(1);
    CN104_sign_in(3) <= VN179_sign_out(1);
    CN104_data_in(4) <= VN267_data_out(1);
    CN104_sign_in(4) <= VN267_sign_out(1);
    CN104_data_in(5) <= VN317_data_out(1);
    CN104_sign_in(5) <= VN317_sign_out(1);
    CN104_data_in(6) <= VN388_data_out(1);
    CN104_sign_in(6) <= VN388_sign_out(1);
    CN104_data_in(7) <= VN396_data_out(1);
    CN104_sign_in(7) <= VN396_sign_out(1);
    CN104_data_in(8) <= VN464_data_out(1);
    CN104_sign_in(8) <= VN464_sign_out(1);
    CN104_data_in(9) <= VN530_data_out(1);
    CN104_sign_in(9) <= VN530_sign_out(1);
    CN104_data_in(10) <= VN605_data_out(1);
    CN104_sign_in(10) <= VN605_sign_out(1);
    CN104_data_in(11) <= VN640_data_out(1);
    CN104_sign_in(11) <= VN640_sign_out(1);
    CN104_data_in(12) <= VN769_data_out(1);
    CN104_sign_in(12) <= VN769_sign_out(1);
    CN104_data_in(13) <= VN811_data_out(1);
    CN104_sign_in(13) <= VN811_sign_out(1);
    CN104_data_in(14) <= VN832_data_out(1);
    CN104_sign_in(14) <= VN832_sign_out(1);
    CN104_data_in(15) <= VN939_data_out(1);
    CN104_sign_in(15) <= VN939_sign_out(1);
    CN104_data_in(16) <= VN970_data_out(1);
    CN104_sign_in(16) <= VN970_sign_out(1);
    CN104_data_in(17) <= VN1043_data_out(1);
    CN104_sign_in(17) <= VN1043_sign_out(1);
    CN104_data_in(18) <= VN1080_data_out(1);
    CN104_sign_in(18) <= VN1080_sign_out(1);
    CN104_data_in(19) <= VN1149_data_out(1);
    CN104_sign_in(19) <= VN1149_sign_out(1);
    CN104_data_in(20) <= VN1204_data_out(1);
    CN104_sign_in(20) <= VN1204_sign_out(1);
    CN104_data_in(21) <= VN1274_data_out(1);
    CN104_sign_in(21) <= VN1274_sign_out(1);
    CN104_data_in(22) <= VN1312_data_out(1);
    CN104_sign_in(22) <= VN1312_sign_out(1);
    CN104_data_in(23) <= VN1454_data_out(1);
    CN104_sign_in(23) <= VN1454_sign_out(1);
    CN104_data_in(24) <= VN1470_data_out(1);
    CN104_sign_in(24) <= VN1470_sign_out(1);
    CN104_data_in(25) <= VN1480_data_out(1);
    CN104_sign_in(25) <= VN1480_sign_out(1);
    CN104_data_in(26) <= VN1489_data_out(1);
    CN104_sign_in(26) <= VN1489_sign_out(1);
    CN104_data_in(27) <= VN1498_data_out(1);
    CN104_sign_in(27) <= VN1498_sign_out(1);
    CN104_data_in(28) <= VN1533_data_out(1);
    CN104_sign_in(28) <= VN1533_sign_out(1);
    CN104_data_in(29) <= VN1663_data_out(1);
    CN104_sign_in(29) <= VN1663_sign_out(1);
    CN104_data_in(30) <= VN1714_data_out(1);
    CN104_sign_in(30) <= VN1714_sign_out(1);
    CN104_data_in(31) <= VN1750_data_out(1);
    CN104_sign_in(31) <= VN1750_sign_out(1);
    CN105_data_in(0) <= VN13_data_out(1);
    CN105_sign_in(0) <= VN13_sign_out(1);
    CN105_data_in(1) <= VN146_data_out(1);
    CN105_sign_in(1) <= VN146_sign_out(1);
    CN105_data_in(2) <= VN197_data_out(1);
    CN105_sign_in(2) <= VN197_sign_out(1);
    CN105_data_in(3) <= VN237_data_out(1);
    CN105_sign_in(3) <= VN237_sign_out(1);
    CN105_data_in(4) <= VN300_data_out(1);
    CN105_sign_in(4) <= VN300_sign_out(1);
    CN105_data_in(5) <= VN338_data_out(1);
    CN105_sign_in(5) <= VN338_sign_out(1);
    CN105_data_in(6) <= VN422_data_out(1);
    CN105_sign_in(6) <= VN422_sign_out(1);
    CN105_data_in(7) <= VN462_data_out(1);
    CN105_sign_in(7) <= VN462_sign_out(1);
    CN105_data_in(8) <= VN593_data_out(1);
    CN105_sign_in(8) <= VN593_sign_out(1);
    CN105_data_in(9) <= VN705_data_out(1);
    CN105_sign_in(9) <= VN705_sign_out(1);
    CN105_data_in(10) <= VN737_data_out(1);
    CN105_sign_in(10) <= VN737_sign_out(1);
    CN105_data_in(11) <= VN806_data_out(1);
    CN105_sign_in(11) <= VN806_sign_out(1);
    CN105_data_in(12) <= VN844_data_out(1);
    CN105_sign_in(12) <= VN844_sign_out(1);
    CN105_data_in(13) <= VN922_data_out(1);
    CN105_sign_in(13) <= VN922_sign_out(1);
    CN105_data_in(14) <= VN966_data_out(1);
    CN105_sign_in(14) <= VN966_sign_out(1);
    CN105_data_in(15) <= VN1044_data_out(1);
    CN105_sign_in(15) <= VN1044_sign_out(1);
    CN105_data_in(16) <= VN1089_data_out(1);
    CN105_sign_in(16) <= VN1089_sign_out(1);
    CN105_data_in(17) <= VN1172_data_out(1);
    CN105_sign_in(17) <= VN1172_sign_out(1);
    CN105_data_in(18) <= VN1225_data_out(1);
    CN105_sign_in(18) <= VN1225_sign_out(1);
    CN105_data_in(19) <= VN1351_data_out(1);
    CN105_sign_in(19) <= VN1351_sign_out(1);
    CN105_data_in(20) <= VN1418_data_out(1);
    CN105_sign_in(20) <= VN1418_sign_out(1);
    CN105_data_in(21) <= VN1428_data_out(1);
    CN105_sign_in(21) <= VN1428_sign_out(1);
    CN105_data_in(22) <= VN1443_data_out(1);
    CN105_sign_in(22) <= VN1443_sign_out(1);
    CN105_data_in(23) <= VN1497_data_out(1);
    CN105_sign_in(23) <= VN1497_sign_out(1);
    CN105_data_in(24) <= VN1526_data_out(1);
    CN105_sign_in(24) <= VN1526_sign_out(1);
    CN105_data_in(25) <= VN1709_data_out(1);
    CN105_sign_in(25) <= VN1709_sign_out(1);
    CN105_data_in(26) <= VN1783_data_out(1);
    CN105_sign_in(26) <= VN1783_sign_out(1);
    CN105_data_in(27) <= VN1806_data_out(1);
    CN105_sign_in(27) <= VN1806_sign_out(1);
    CN105_data_in(28) <= VN1966_data_out(1);
    CN105_sign_in(28) <= VN1966_sign_out(1);
    CN105_data_in(29) <= VN2012_data_out(1);
    CN105_sign_in(29) <= VN2012_sign_out(1);
    CN105_data_in(30) <= VN2044_data_out(1);
    CN105_sign_in(30) <= VN2044_sign_out(1);
    CN105_data_in(31) <= VN2046_data_out(1);
    CN105_sign_in(31) <= VN2046_sign_out(1);
    CN106_data_in(0) <= VN12_data_out(1);
    CN106_sign_in(0) <= VN12_sign_out(1);
    CN106_data_in(1) <= VN157_data_out(1);
    CN106_sign_in(1) <= VN157_sign_out(1);
    CN106_data_in(2) <= VN223_data_out(1);
    CN106_sign_in(2) <= VN223_sign_out(1);
    CN106_data_in(3) <= VN272_data_out(1);
    CN106_sign_in(3) <= VN272_sign_out(1);
    CN106_data_in(4) <= VN312_data_out(1);
    CN106_sign_in(4) <= VN312_sign_out(1);
    CN106_data_in(5) <= VN333_data_out(1);
    CN106_sign_in(5) <= VN333_sign_out(1);
    CN106_data_in(6) <= VN412_data_out(1);
    CN106_sign_in(6) <= VN412_sign_out(1);
    CN106_data_in(7) <= VN529_data_out(1);
    CN106_sign_in(7) <= VN529_sign_out(1);
    CN106_data_in(8) <= VN610_data_out(1);
    CN106_sign_in(8) <= VN610_sign_out(1);
    CN106_data_in(9) <= VN700_data_out(1);
    CN106_sign_in(9) <= VN700_sign_out(1);
    CN106_data_in(10) <= VN744_data_out(1);
    CN106_sign_in(10) <= VN744_sign_out(1);
    CN106_data_in(11) <= VN812_data_out(1);
    CN106_sign_in(11) <= VN812_sign_out(1);
    CN106_data_in(12) <= VN853_data_out(1);
    CN106_sign_in(12) <= VN853_sign_out(1);
    CN106_data_in(13) <= VN929_data_out(1);
    CN106_sign_in(13) <= VN929_sign_out(1);
    CN106_data_in(14) <= VN986_data_out(1);
    CN106_sign_in(14) <= VN986_sign_out(1);
    CN106_data_in(15) <= VN1021_data_out(1);
    CN106_sign_in(15) <= VN1021_sign_out(1);
    CN106_data_in(16) <= VN1085_data_out(1);
    CN106_sign_in(16) <= VN1085_sign_out(1);
    CN106_data_in(17) <= VN1170_data_out(1);
    CN106_sign_in(17) <= VN1170_sign_out(1);
    CN106_data_in(18) <= VN1246_data_out(1);
    CN106_sign_in(18) <= VN1246_sign_out(1);
    CN106_data_in(19) <= VN1280_data_out(1);
    CN106_sign_in(19) <= VN1280_sign_out(1);
    CN106_data_in(20) <= VN1295_data_out(1);
    CN106_sign_in(20) <= VN1295_sign_out(1);
    CN106_data_in(21) <= VN1352_data_out(1);
    CN106_sign_in(21) <= VN1352_sign_out(1);
    CN106_data_in(22) <= VN1394_data_out(1);
    CN106_sign_in(22) <= VN1394_sign_out(1);
    CN106_data_in(23) <= VN1514_data_out(1);
    CN106_sign_in(23) <= VN1514_sign_out(1);
    CN106_data_in(24) <= VN1594_data_out(1);
    CN106_sign_in(24) <= VN1594_sign_out(1);
    CN106_data_in(25) <= VN1637_data_out(1);
    CN106_sign_in(25) <= VN1637_sign_out(1);
    CN106_data_in(26) <= VN1803_data_out(1);
    CN106_sign_in(26) <= VN1803_sign_out(1);
    CN106_data_in(27) <= VN1807_data_out(1);
    CN106_sign_in(27) <= VN1807_sign_out(1);
    CN106_data_in(28) <= VN1885_data_out(1);
    CN106_sign_in(28) <= VN1885_sign_out(1);
    CN106_data_in(29) <= VN1938_data_out(1);
    CN106_sign_in(29) <= VN1938_sign_out(1);
    CN106_data_in(30) <= VN1953_data_out(1);
    CN106_sign_in(30) <= VN1953_sign_out(1);
    CN106_data_in(31) <= VN1963_data_out(1);
    CN106_sign_in(31) <= VN1963_sign_out(1);
    CN107_data_in(0) <= VN110_data_out(1);
    CN107_sign_in(0) <= VN110_sign_out(1);
    CN107_data_in(1) <= VN127_data_out(1);
    CN107_sign_in(1) <= VN127_sign_out(1);
    CN107_data_in(2) <= VN207_data_out(1);
    CN107_sign_in(2) <= VN207_sign_out(1);
    CN107_data_in(3) <= VN230_data_out(1);
    CN107_sign_in(3) <= VN230_sign_out(1);
    CN107_data_in(4) <= VN323_data_out(1);
    CN107_sign_in(4) <= VN323_sign_out(1);
    CN107_data_in(5) <= VN335_data_out(1);
    CN107_sign_in(5) <= VN335_sign_out(1);
    CN107_data_in(6) <= VN469_data_out(1);
    CN107_sign_in(6) <= VN469_sign_out(1);
    CN107_data_in(7) <= VN586_data_out(1);
    CN107_sign_in(7) <= VN586_sign_out(1);
    CN107_data_in(8) <= VN656_data_out(1);
    CN107_sign_in(8) <= VN656_sign_out(1);
    CN107_data_in(9) <= VN681_data_out(1);
    CN107_sign_in(9) <= VN681_sign_out(1);
    CN107_data_in(10) <= VN728_data_out(1);
    CN107_sign_in(10) <= VN728_sign_out(1);
    CN107_data_in(11) <= VN801_data_out(1);
    CN107_sign_in(11) <= VN801_sign_out(1);
    CN107_data_in(12) <= VN880_data_out(1);
    CN107_sign_in(12) <= VN880_sign_out(1);
    CN107_data_in(13) <= VN895_data_out(1);
    CN107_sign_in(13) <= VN895_sign_out(1);
    CN107_data_in(14) <= VN949_data_out(1);
    CN107_sign_in(14) <= VN949_sign_out(1);
    CN107_data_in(15) <= VN1153_data_out(1);
    CN107_sign_in(15) <= VN1153_sign_out(1);
    CN107_data_in(16) <= VN1202_data_out(1);
    CN107_sign_in(16) <= VN1202_sign_out(1);
    CN107_data_in(17) <= VN1244_data_out(1);
    CN107_sign_in(17) <= VN1244_sign_out(1);
    CN107_data_in(18) <= VN1302_data_out(1);
    CN107_sign_in(18) <= VN1302_sign_out(1);
    CN107_data_in(19) <= VN1333_data_out(1);
    CN107_sign_in(19) <= VN1333_sign_out(1);
    CN107_data_in(20) <= VN1415_data_out(1);
    CN107_sign_in(20) <= VN1415_sign_out(1);
    CN107_data_in(21) <= VN1445_data_out(1);
    CN107_sign_in(21) <= VN1445_sign_out(1);
    CN107_data_in(22) <= VN1729_data_out(1);
    CN107_sign_in(22) <= VN1729_sign_out(1);
    CN107_data_in(23) <= VN1793_data_out(1);
    CN107_sign_in(23) <= VN1793_sign_out(1);
    CN107_data_in(24) <= VN1797_data_out(1);
    CN107_sign_in(24) <= VN1797_sign_out(1);
    CN107_data_in(25) <= VN1817_data_out(1);
    CN107_sign_in(25) <= VN1817_sign_out(1);
    CN107_data_in(26) <= VN1835_data_out(1);
    CN107_sign_in(26) <= VN1835_sign_out(1);
    CN107_data_in(27) <= VN1889_data_out(1);
    CN107_sign_in(27) <= VN1889_sign_out(1);
    CN107_data_in(28) <= VN1977_data_out(1);
    CN107_sign_in(28) <= VN1977_sign_out(1);
    CN107_data_in(29) <= VN1981_data_out(1);
    CN107_sign_in(29) <= VN1981_sign_out(1);
    CN107_data_in(30) <= VN2045_data_out(1);
    CN107_sign_in(30) <= VN2045_sign_out(1);
    CN107_data_in(31) <= VN2047_data_out(1);
    CN107_sign_in(31) <= VN2047_sign_out(1);
    CN108_data_in(0) <= VN11_data_out(1);
    CN108_sign_in(0) <= VN11_sign_out(1);
    CN108_data_in(1) <= VN105_data_out(1);
    CN108_sign_in(1) <= VN105_sign_out(1);
    CN108_data_in(2) <= VN115_data_out(1);
    CN108_sign_in(2) <= VN115_sign_out(1);
    CN108_data_in(3) <= VN181_data_out(1);
    CN108_sign_in(3) <= VN181_sign_out(1);
    CN108_data_in(4) <= VN238_data_out(1);
    CN108_sign_in(4) <= VN238_sign_out(1);
    CN108_data_in(5) <= VN296_data_out(1);
    CN108_sign_in(5) <= VN296_sign_out(1);
    CN108_data_in(6) <= VN385_data_out(1);
    CN108_sign_in(6) <= VN385_sign_out(1);
    CN108_data_in(7) <= VN418_data_out(1);
    CN108_sign_in(7) <= VN418_sign_out(1);
    CN108_data_in(8) <= VN500_data_out(1);
    CN108_sign_in(8) <= VN500_sign_out(1);
    CN108_data_in(9) <= VN508_data_out(1);
    CN108_sign_in(9) <= VN508_sign_out(1);
    CN108_data_in(10) <= VN583_data_out(1);
    CN108_sign_in(10) <= VN583_sign_out(1);
    CN108_data_in(11) <= VN643_data_out(1);
    CN108_sign_in(11) <= VN643_sign_out(1);
    CN108_data_in(12) <= VN689_data_out(1);
    CN108_sign_in(12) <= VN689_sign_out(1);
    CN108_data_in(13) <= VN730_data_out(1);
    CN108_sign_in(13) <= VN730_sign_out(1);
    CN108_data_in(14) <= VN826_data_out(1);
    CN108_sign_in(14) <= VN826_sign_out(1);
    CN108_data_in(15) <= VN839_data_out(1);
    CN108_sign_in(15) <= VN839_sign_out(1);
    CN108_data_in(16) <= VN893_data_out(1);
    CN108_sign_in(16) <= VN893_sign_out(1);
    CN108_data_in(17) <= VN950_data_out(1);
    CN108_sign_in(17) <= VN950_sign_out(1);
    CN108_data_in(18) <= VN1029_data_out(1);
    CN108_sign_in(18) <= VN1029_sign_out(1);
    CN108_data_in(19) <= VN1108_data_out(1);
    CN108_sign_in(19) <= VN1108_sign_out(1);
    CN108_data_in(20) <= VN1147_data_out(1);
    CN108_sign_in(20) <= VN1147_sign_out(1);
    CN108_data_in(21) <= VN1184_data_out(1);
    CN108_sign_in(21) <= VN1184_sign_out(1);
    CN108_data_in(22) <= VN1299_data_out(1);
    CN108_sign_in(22) <= VN1299_sign_out(1);
    CN108_data_in(23) <= VN1376_data_out(1);
    CN108_sign_in(23) <= VN1376_sign_out(1);
    CN108_data_in(24) <= VN1471_data_out(1);
    CN108_sign_in(24) <= VN1471_sign_out(1);
    CN108_data_in(25) <= VN1523_data_out(1);
    CN108_sign_in(25) <= VN1523_sign_out(1);
    CN108_data_in(26) <= VN1548_data_out(1);
    CN108_sign_in(26) <= VN1548_sign_out(1);
    CN108_data_in(27) <= VN1595_data_out(1);
    CN108_sign_in(27) <= VN1595_sign_out(1);
    CN108_data_in(28) <= VN1644_data_out(1);
    CN108_sign_in(28) <= VN1644_sign_out(1);
    CN108_data_in(29) <= VN1683_data_out(1);
    CN108_sign_in(29) <= VN1683_sign_out(1);
    CN108_data_in(30) <= VN1717_data_out(1);
    CN108_sign_in(30) <= VN1717_sign_out(1);
    CN108_data_in(31) <= VN1751_data_out(1);
    CN108_sign_in(31) <= VN1751_sign_out(1);
    CN109_data_in(0) <= VN10_data_out(1);
    CN109_sign_in(0) <= VN10_sign_out(1);
    CN109_data_in(1) <= VN100_data_out(1);
    CN109_sign_in(1) <= VN100_sign_out(1);
    CN109_data_in(2) <= VN160_data_out(1);
    CN109_sign_in(2) <= VN160_sign_out(1);
    CN109_data_in(3) <= VN171_data_out(1);
    CN109_sign_in(3) <= VN171_sign_out(1);
    CN109_data_in(4) <= VN266_data_out(1);
    CN109_sign_in(4) <= VN266_sign_out(1);
    CN109_data_in(5) <= VN362_data_out(1);
    CN109_sign_in(5) <= VN362_sign_out(1);
    CN109_data_in(6) <= VN454_data_out(1);
    CN109_sign_in(6) <= VN454_sign_out(1);
    CN109_data_in(7) <= VN598_data_out(1);
    CN109_sign_in(7) <= VN598_sign_out(1);
    CN109_data_in(8) <= VN711_data_out(1);
    CN109_sign_in(8) <= VN711_sign_out(1);
    CN109_data_in(9) <= VN754_data_out(1);
    CN109_sign_in(9) <= VN754_sign_out(1);
    CN109_data_in(10) <= VN778_data_out(1);
    CN109_sign_in(10) <= VN778_sign_out(1);
    CN109_data_in(11) <= VN927_data_out(1);
    CN109_sign_in(11) <= VN927_sign_out(1);
    CN109_data_in(12) <= VN985_data_out(1);
    CN109_sign_in(12) <= VN985_sign_out(1);
    CN109_data_in(13) <= VN1129_data_out(1);
    CN109_sign_in(13) <= VN1129_sign_out(1);
    CN109_data_in(14) <= VN1169_data_out(1);
    CN109_sign_in(14) <= VN1169_sign_out(1);
    CN109_data_in(15) <= VN1186_data_out(1);
    CN109_sign_in(15) <= VN1186_sign_out(1);
    CN109_data_in(16) <= VN1258_data_out(1);
    CN109_sign_in(16) <= VN1258_sign_out(1);
    CN109_data_in(17) <= VN1303_data_out(1);
    CN109_sign_in(17) <= VN1303_sign_out(1);
    CN109_data_in(18) <= VN1337_data_out(1);
    CN109_sign_in(18) <= VN1337_sign_out(1);
    CN109_data_in(19) <= VN1588_data_out(1);
    CN109_sign_in(19) <= VN1588_sign_out(1);
    CN109_data_in(20) <= VN1615_data_out(1);
    CN109_sign_in(20) <= VN1615_sign_out(1);
    CN109_data_in(21) <= VN1672_data_out(1);
    CN109_sign_in(21) <= VN1672_sign_out(1);
    CN109_data_in(22) <= VN1732_data_out(1);
    CN109_sign_in(22) <= VN1732_sign_out(1);
    CN109_data_in(23) <= VN1734_data_out(1);
    CN109_sign_in(23) <= VN1734_sign_out(1);
    CN109_data_in(24) <= VN1767_data_out(1);
    CN109_sign_in(24) <= VN1767_sign_out(1);
    CN109_data_in(25) <= VN1858_data_out(1);
    CN109_sign_in(25) <= VN1858_sign_out(1);
    CN109_data_in(26) <= VN1893_data_out(1);
    CN109_sign_in(26) <= VN1893_sign_out(1);
    CN109_data_in(27) <= VN1927_data_out(1);
    CN109_sign_in(27) <= VN1927_sign_out(1);
    CN109_data_in(28) <= VN1939_data_out(1);
    CN109_sign_in(28) <= VN1939_sign_out(1);
    CN109_data_in(29) <= VN2007_data_out(1);
    CN109_sign_in(29) <= VN2007_sign_out(1);
    CN109_data_in(30) <= VN2029_data_out(1);
    CN109_sign_in(30) <= VN2029_sign_out(1);
    CN109_data_in(31) <= VN2042_data_out(1);
    CN109_sign_in(31) <= VN2042_sign_out(1);
    CN110_data_in(0) <= VN9_data_out(1);
    CN110_sign_in(0) <= VN9_sign_out(1);
    CN110_data_in(1) <= VN83_data_out(1);
    CN110_sign_in(1) <= VN83_sign_out(1);
    CN110_data_in(2) <= VN118_data_out(1);
    CN110_sign_in(2) <= VN118_sign_out(1);
    CN110_data_in(3) <= VN212_data_out(1);
    CN110_sign_in(3) <= VN212_sign_out(1);
    CN110_data_in(4) <= VN225_data_out(1);
    CN110_sign_in(4) <= VN225_sign_out(1);
    CN110_data_in(5) <= VN326_data_out(1);
    CN110_sign_in(5) <= VN326_sign_out(1);
    CN110_data_in(6) <= VN345_data_out(1);
    CN110_sign_in(6) <= VN345_sign_out(1);
    CN110_data_in(7) <= VN446_data_out(1);
    CN110_sign_in(7) <= VN446_sign_out(1);
    CN110_data_in(8) <= VN504_data_out(1);
    CN110_sign_in(8) <= VN504_sign_out(1);
    CN110_data_in(9) <= VN536_data_out(1);
    CN110_sign_in(9) <= VN536_sign_out(1);
    CN110_data_in(10) <= VN591_data_out(1);
    CN110_sign_in(10) <= VN591_sign_out(1);
    CN110_data_in(11) <= VN639_data_out(1);
    CN110_sign_in(11) <= VN639_sign_out(1);
    CN110_data_in(12) <= VN710_data_out(1);
    CN110_sign_in(12) <= VN710_sign_out(1);
    CN110_data_in(13) <= VN736_data_out(1);
    CN110_sign_in(13) <= VN736_sign_out(1);
    CN110_data_in(14) <= VN816_data_out(1);
    CN110_sign_in(14) <= VN816_sign_out(1);
    CN110_data_in(15) <= VN847_data_out(1);
    CN110_sign_in(15) <= VN847_sign_out(1);
    CN110_data_in(16) <= VN909_data_out(1);
    CN110_sign_in(16) <= VN909_sign_out(1);
    CN110_data_in(17) <= VN977_data_out(1);
    CN110_sign_in(17) <= VN977_sign_out(1);
    CN110_data_in(18) <= VN1107_data_out(1);
    CN110_sign_in(18) <= VN1107_sign_out(1);
    CN110_data_in(19) <= VN1136_data_out(1);
    CN110_sign_in(19) <= VN1136_sign_out(1);
    CN110_data_in(20) <= VN1165_data_out(1);
    CN110_sign_in(20) <= VN1165_sign_out(1);
    CN110_data_in(21) <= VN1173_data_out(1);
    CN110_sign_in(21) <= VN1173_sign_out(1);
    CN110_data_in(22) <= VN1261_data_out(1);
    CN110_sign_in(22) <= VN1261_sign_out(1);
    CN110_data_in(23) <= VN1294_data_out(1);
    CN110_sign_in(23) <= VN1294_sign_out(1);
    CN110_data_in(24) <= VN1341_data_out(1);
    CN110_sign_in(24) <= VN1341_sign_out(1);
    CN110_data_in(25) <= VN1439_data_out(1);
    CN110_sign_in(25) <= VN1439_sign_out(1);
    CN110_data_in(26) <= VN1458_data_out(1);
    CN110_sign_in(26) <= VN1458_sign_out(1);
    CN110_data_in(27) <= VN1494_data_out(1);
    CN110_sign_in(27) <= VN1494_sign_out(1);
    CN110_data_in(28) <= VN1505_data_out(1);
    CN110_sign_in(28) <= VN1505_sign_out(1);
    CN110_data_in(29) <= VN1628_data_out(1);
    CN110_sign_in(29) <= VN1628_sign_out(1);
    CN110_data_in(30) <= VN1704_data_out(1);
    CN110_sign_in(30) <= VN1704_sign_out(1);
    CN110_data_in(31) <= VN1752_data_out(1);
    CN110_sign_in(31) <= VN1752_sign_out(1);
    CN111_data_in(0) <= VN8_data_out(1);
    CN111_sign_in(0) <= VN8_sign_out(1);
    CN111_data_in(1) <= VN90_data_out(1);
    CN111_sign_in(1) <= VN90_sign_out(1);
    CN111_data_in(2) <= VN138_data_out(1);
    CN111_sign_in(2) <= VN138_sign_out(1);
    CN111_data_in(3) <= VN177_data_out(1);
    CN111_sign_in(3) <= VN177_sign_out(1);
    CN111_data_in(4) <= VN252_data_out(1);
    CN111_sign_in(4) <= VN252_sign_out(1);
    CN111_data_in(5) <= VN287_data_out(1);
    CN111_sign_in(5) <= VN287_sign_out(1);
    CN111_data_in(6) <= VN357_data_out(1);
    CN111_sign_in(6) <= VN357_sign_out(1);
    CN111_data_in(7) <= VN405_data_out(1);
    CN111_sign_in(7) <= VN405_sign_out(1);
    CN111_data_in(8) <= VN451_data_out(1);
    CN111_sign_in(8) <= VN451_sign_out(1);
    CN111_data_in(9) <= VN534_data_out(1);
    CN111_sign_in(9) <= VN534_sign_out(1);
    CN111_data_in(10) <= VN567_data_out(1);
    CN111_sign_in(10) <= VN567_sign_out(1);
    CN111_data_in(11) <= VN665_data_out(1);
    CN111_sign_in(11) <= VN665_sign_out(1);
    CN111_data_in(12) <= VN687_data_out(1);
    CN111_sign_in(12) <= VN687_sign_out(1);
    CN111_data_in(13) <= VN747_data_out(1);
    CN111_sign_in(13) <= VN747_sign_out(1);
    CN111_data_in(14) <= VN818_data_out(1);
    CN111_sign_in(14) <= VN818_sign_out(1);
    CN111_data_in(15) <= VN868_data_out(1);
    CN111_sign_in(15) <= VN868_sign_out(1);
    CN111_data_in(16) <= VN911_data_out(1);
    CN111_sign_in(16) <= VN911_sign_out(1);
    CN111_data_in(17) <= VN994_data_out(1);
    CN111_sign_in(17) <= VN994_sign_out(1);
    CN111_data_in(18) <= VN1033_data_out(1);
    CN111_sign_in(18) <= VN1033_sign_out(1);
    CN111_data_in(19) <= VN1092_data_out(1);
    CN111_sign_in(19) <= VN1092_sign_out(1);
    CN111_data_in(20) <= VN1159_data_out(1);
    CN111_sign_in(20) <= VN1159_sign_out(1);
    CN111_data_in(21) <= VN1203_data_out(1);
    CN111_sign_in(21) <= VN1203_sign_out(1);
    CN111_data_in(22) <= VN1218_data_out(1);
    CN111_sign_in(22) <= VN1218_sign_out(1);
    CN111_data_in(23) <= VN1247_data_out(1);
    CN111_sign_in(23) <= VN1247_sign_out(1);
    CN111_data_in(24) <= VN1314_data_out(1);
    CN111_sign_in(24) <= VN1314_sign_out(1);
    CN111_data_in(25) <= VN1390_data_out(1);
    CN111_sign_in(25) <= VN1390_sign_out(1);
    CN111_data_in(26) <= VN1465_data_out(1);
    CN111_sign_in(26) <= VN1465_sign_out(1);
    CN111_data_in(27) <= VN1536_data_out(1);
    CN111_sign_in(27) <= VN1536_sign_out(1);
    CN111_data_in(28) <= VN1550_data_out(1);
    CN111_sign_in(28) <= VN1550_sign_out(1);
    CN111_data_in(29) <= VN1668_data_out(1);
    CN111_sign_in(29) <= VN1668_sign_out(1);
    CN111_data_in(30) <= VN1782_data_out(1);
    CN111_sign_in(30) <= VN1782_sign_out(1);
    CN111_data_in(31) <= VN1826_data_out(1);
    CN111_sign_in(31) <= VN1826_sign_out(1);
    CN112_data_in(0) <= VN7_data_out(1);
    CN112_sign_in(0) <= VN7_sign_out(1);
    CN112_data_in(1) <= VN54_data_out(1);
    CN112_sign_in(1) <= VN54_sign_out(1);
    CN112_data_in(2) <= VN148_data_out(1);
    CN112_sign_in(2) <= VN148_sign_out(1);
    CN112_data_in(3) <= VN205_data_out(1);
    CN112_sign_in(3) <= VN205_sign_out(1);
    CN112_data_in(4) <= VN233_data_out(1);
    CN112_sign_in(4) <= VN233_sign_out(1);
    CN112_data_in(5) <= VN305_data_out(1);
    CN112_sign_in(5) <= VN305_sign_out(1);
    CN112_data_in(6) <= VN369_data_out(1);
    CN112_sign_in(6) <= VN369_sign_out(1);
    CN112_data_in(7) <= VN398_data_out(1);
    CN112_sign_in(7) <= VN398_sign_out(1);
    CN112_data_in(8) <= VN497_data_out(1);
    CN112_sign_in(8) <= VN497_sign_out(1);
    CN112_data_in(9) <= VN513_data_out(1);
    CN112_sign_in(9) <= VN513_sign_out(1);
    CN112_data_in(10) <= VN577_data_out(1);
    CN112_sign_in(10) <= VN577_sign_out(1);
    CN112_data_in(11) <= VN652_data_out(1);
    CN112_sign_in(11) <= VN652_sign_out(1);
    CN112_data_in(12) <= VN669_data_out(1);
    CN112_sign_in(12) <= VN669_sign_out(1);
    CN112_data_in(13) <= VN755_data_out(1);
    CN112_sign_in(13) <= VN755_sign_out(1);
    CN112_data_in(14) <= VN788_data_out(1);
    CN112_sign_in(14) <= VN788_sign_out(1);
    CN112_data_in(15) <= VN882_data_out(1);
    CN112_sign_in(15) <= VN882_sign_out(1);
    CN112_data_in(16) <= VN896_data_out(1);
    CN112_sign_in(16) <= VN896_sign_out(1);
    CN112_data_in(17) <= VN999_data_out(1);
    CN112_sign_in(17) <= VN999_sign_out(1);
    CN112_data_in(18) <= VN1028_data_out(1);
    CN112_sign_in(18) <= VN1028_sign_out(1);
    CN112_data_in(19) <= VN1060_data_out(1);
    CN112_sign_in(19) <= VN1060_sign_out(1);
    CN112_data_in(20) <= VN1094_data_out(1);
    CN112_sign_in(20) <= VN1094_sign_out(1);
    CN112_data_in(21) <= VN1157_data_out(1);
    CN112_sign_in(21) <= VN1157_sign_out(1);
    CN112_data_in(22) <= VN1321_data_out(1);
    CN112_sign_in(22) <= VN1321_sign_out(1);
    CN112_data_in(23) <= VN1340_data_out(1);
    CN112_sign_in(23) <= VN1340_sign_out(1);
    CN112_data_in(24) <= VN1473_data_out(1);
    CN112_sign_in(24) <= VN1473_sign_out(1);
    CN112_data_in(25) <= VN1518_data_out(1);
    CN112_sign_in(25) <= VN1518_sign_out(1);
    CN112_data_in(26) <= VN1524_data_out(1);
    CN112_sign_in(26) <= VN1524_sign_out(1);
    CN112_data_in(27) <= VN1598_data_out(1);
    CN112_sign_in(27) <= VN1598_sign_out(1);
    CN112_data_in(28) <= VN1640_data_out(1);
    CN112_sign_in(28) <= VN1640_sign_out(1);
    CN112_data_in(29) <= VN1667_data_out(1);
    CN112_sign_in(29) <= VN1667_sign_out(1);
    CN112_data_in(30) <= VN1698_data_out(1);
    CN112_sign_in(30) <= VN1698_sign_out(1);
    CN112_data_in(31) <= VN1753_data_out(1);
    CN112_sign_in(31) <= VN1753_sign_out(1);
    CN113_data_in(0) <= VN6_data_out(1);
    CN113_sign_in(0) <= VN6_sign_out(1);
    CN113_data_in(1) <= VN108_data_out(1);
    CN113_sign_in(1) <= VN108_sign_out(1);
    CN113_data_in(2) <= VN143_data_out(1);
    CN113_sign_in(2) <= VN143_sign_out(1);
    CN113_data_in(3) <= VN202_data_out(1);
    CN113_sign_in(3) <= VN202_sign_out(1);
    CN113_data_in(4) <= VN253_data_out(1);
    CN113_sign_in(4) <= VN253_sign_out(1);
    CN113_data_in(5) <= VN314_data_out(1);
    CN113_sign_in(5) <= VN314_sign_out(1);
    CN113_data_in(6) <= VN339_data_out(1);
    CN113_sign_in(6) <= VN339_sign_out(1);
    CN113_data_in(7) <= VN429_data_out(1);
    CN113_sign_in(7) <= VN429_sign_out(1);
    CN113_data_in(8) <= VN550_data_out(1);
    CN113_sign_in(8) <= VN550_sign_out(1);
    CN113_data_in(9) <= VN570_data_out(1);
    CN113_sign_in(9) <= VN570_sign_out(1);
    CN113_data_in(10) <= VN622_data_out(1);
    CN113_sign_in(10) <= VN622_sign_out(1);
    CN113_data_in(11) <= VN671_data_out(1);
    CN113_sign_in(11) <= VN671_sign_out(1);
    CN113_data_in(12) <= VN729_data_out(1);
    CN113_sign_in(12) <= VN729_sign_out(1);
    CN113_data_in(13) <= VN824_data_out(1);
    CN113_sign_in(13) <= VN824_sign_out(1);
    CN113_data_in(14) <= VN878_data_out(1);
    CN113_sign_in(14) <= VN878_sign_out(1);
    CN113_data_in(15) <= VN928_data_out(1);
    CN113_sign_in(15) <= VN928_sign_out(1);
    CN113_data_in(16) <= VN1011_data_out(1);
    CN113_sign_in(16) <= VN1011_sign_out(1);
    CN113_data_in(17) <= VN1066_data_out(1);
    CN113_sign_in(17) <= VN1066_sign_out(1);
    CN113_data_in(18) <= VN1134_data_out(1);
    CN113_sign_in(18) <= VN1134_sign_out(1);
    CN113_data_in(19) <= VN1194_data_out(1);
    CN113_sign_in(19) <= VN1194_sign_out(1);
    CN113_data_in(20) <= VN1243_data_out(1);
    CN113_sign_in(20) <= VN1243_sign_out(1);
    CN113_data_in(21) <= VN1305_data_out(1);
    CN113_sign_in(21) <= VN1305_sign_out(1);
    CN113_data_in(22) <= VN1329_data_out(1);
    CN113_sign_in(22) <= VN1329_sign_out(1);
    CN113_data_in(23) <= VN1393_data_out(1);
    CN113_sign_in(23) <= VN1393_sign_out(1);
    CN113_data_in(24) <= VN1440_data_out(1);
    CN113_sign_in(24) <= VN1440_sign_out(1);
    CN113_data_in(25) <= VN1503_data_out(1);
    CN113_sign_in(25) <= VN1503_sign_out(1);
    CN113_data_in(26) <= VN1610_data_out(1);
    CN113_sign_in(26) <= VN1610_sign_out(1);
    CN113_data_in(27) <= VN1677_data_out(1);
    CN113_sign_in(27) <= VN1677_sign_out(1);
    CN113_data_in(28) <= VN1728_data_out(1);
    CN113_sign_in(28) <= VN1728_sign_out(1);
    CN113_data_in(29) <= VN1737_data_out(1);
    CN113_sign_in(29) <= VN1737_sign_out(1);
    CN113_data_in(30) <= VN1794_data_out(1);
    CN113_sign_in(30) <= VN1794_sign_out(1);
    CN113_data_in(31) <= VN1827_data_out(1);
    CN113_sign_in(31) <= VN1827_sign_out(1);
    CN114_data_in(0) <= VN5_data_out(1);
    CN114_sign_in(0) <= VN5_sign_out(1);
    CN114_data_in(1) <= VN88_data_out(1);
    CN114_sign_in(1) <= VN88_sign_out(1);
    CN114_data_in(2) <= VN149_data_out(1);
    CN114_sign_in(2) <= VN149_sign_out(1);
    CN114_data_in(3) <= VN216_data_out(1);
    CN114_sign_in(3) <= VN216_sign_out(1);
    CN114_data_in(4) <= VN268_data_out(1);
    CN114_sign_in(4) <= VN268_sign_out(1);
    CN114_data_in(5) <= VN309_data_out(1);
    CN114_sign_in(5) <= VN309_sign_out(1);
    CN114_data_in(6) <= VN387_data_out(1);
    CN114_sign_in(6) <= VN387_sign_out(1);
    CN114_data_in(7) <= VN439_data_out(1);
    CN114_sign_in(7) <= VN439_sign_out(1);
    CN114_data_in(8) <= VN461_data_out(1);
    CN114_sign_in(8) <= VN461_sign_out(1);
    CN114_data_in(9) <= VN553_data_out(1);
    CN114_sign_in(9) <= VN553_sign_out(1);
    CN114_data_in(10) <= VN574_data_out(1);
    CN114_sign_in(10) <= VN574_sign_out(1);
    CN114_data_in(11) <= VN667_data_out(1);
    CN114_sign_in(11) <= VN667_sign_out(1);
    CN114_data_in(12) <= VN712_data_out(1);
    CN114_sign_in(12) <= VN712_sign_out(1);
    CN114_data_in(13) <= VN743_data_out(1);
    CN114_sign_in(13) <= VN743_sign_out(1);
    CN114_data_in(14) <= VN781_data_out(1);
    CN114_sign_in(14) <= VN781_sign_out(1);
    CN114_data_in(15) <= VN842_data_out(1);
    CN114_sign_in(15) <= VN842_sign_out(1);
    CN114_data_in(16) <= VN892_data_out(1);
    CN114_sign_in(16) <= VN892_sign_out(1);
    CN114_data_in(17) <= VN998_data_out(1);
    CN114_sign_in(17) <= VN998_sign_out(1);
    CN114_data_in(18) <= VN1018_data_out(1);
    CN114_sign_in(18) <= VN1018_sign_out(1);
    CN114_data_in(19) <= VN1099_data_out(1);
    CN114_sign_in(19) <= VN1099_sign_out(1);
    CN114_data_in(20) <= VN1180_data_out(1);
    CN114_sign_in(20) <= VN1180_sign_out(1);
    CN114_data_in(21) <= VN1271_data_out(1);
    CN114_sign_in(21) <= VN1271_sign_out(1);
    CN114_data_in(22) <= VN1307_data_out(1);
    CN114_sign_in(22) <= VN1307_sign_out(1);
    CN114_data_in(23) <= VN1373_data_out(1);
    CN114_sign_in(23) <= VN1373_sign_out(1);
    CN114_data_in(24) <= VN1422_data_out(1);
    CN114_sign_in(24) <= VN1422_sign_out(1);
    CN114_data_in(25) <= VN1429_data_out(1);
    CN114_sign_in(25) <= VN1429_sign_out(1);
    CN114_data_in(26) <= VN1486_data_out(1);
    CN114_sign_in(26) <= VN1486_sign_out(1);
    CN114_data_in(27) <= VN1555_data_out(1);
    CN114_sign_in(27) <= VN1555_sign_out(1);
    CN114_data_in(28) <= VN1611_data_out(1);
    CN114_sign_in(28) <= VN1611_sign_out(1);
    CN114_data_in(29) <= VN1736_data_out(1);
    CN114_sign_in(29) <= VN1736_sign_out(1);
    CN114_data_in(30) <= VN1809_data_out(1);
    CN114_sign_in(30) <= VN1809_sign_out(1);
    CN114_data_in(31) <= VN1828_data_out(1);
    CN114_sign_in(31) <= VN1828_sign_out(1);
    CN115_data_in(0) <= VN4_data_out(1);
    CN115_sign_in(0) <= VN4_sign_out(1);
    CN115_data_in(1) <= VN68_data_out(1);
    CN115_sign_in(1) <= VN68_sign_out(1);
    CN115_data_in(2) <= VN137_data_out(1);
    CN115_sign_in(2) <= VN137_sign_out(1);
    CN115_data_in(3) <= VN209_data_out(1);
    CN115_sign_in(3) <= VN209_sign_out(1);
    CN115_data_in(4) <= VN264_data_out(1);
    CN115_sign_in(4) <= VN264_sign_out(1);
    CN115_data_in(5) <= VN315_data_out(1);
    CN115_sign_in(5) <= VN315_sign_out(1);
    CN115_data_in(6) <= VN372_data_out(1);
    CN115_sign_in(6) <= VN372_sign_out(1);
    CN115_data_in(7) <= VN433_data_out(1);
    CN115_sign_in(7) <= VN433_sign_out(1);
    CN115_data_in(8) <= VN473_data_out(1);
    CN115_sign_in(8) <= VN473_sign_out(1);
    CN115_data_in(9) <= VN537_data_out(1);
    CN115_sign_in(9) <= VN537_sign_out(1);
    CN115_data_in(10) <= VN564_data_out(1);
    CN115_sign_in(10) <= VN564_sign_out(1);
    CN115_data_in(11) <= VN654_data_out(1);
    CN115_sign_in(11) <= VN654_sign_out(1);
    CN115_data_in(12) <= VN688_data_out(1);
    CN115_sign_in(12) <= VN688_sign_out(1);
    CN115_data_in(13) <= VN771_data_out(1);
    CN115_sign_in(13) <= VN771_sign_out(1);
    CN115_data_in(14) <= VN789_data_out(1);
    CN115_sign_in(14) <= VN789_sign_out(1);
    CN115_data_in(15) <= VN864_data_out(1);
    CN115_sign_in(15) <= VN864_sign_out(1);
    CN115_data_in(16) <= VN920_data_out(1);
    CN115_sign_in(16) <= VN920_sign_out(1);
    CN115_data_in(17) <= VN992_data_out(1);
    CN115_sign_in(17) <= VN992_sign_out(1);
    CN115_data_in(18) <= VN1039_data_out(1);
    CN115_sign_in(18) <= VN1039_sign_out(1);
    CN115_data_in(19) <= VN1111_data_out(1);
    CN115_sign_in(19) <= VN1111_sign_out(1);
    CN115_data_in(20) <= VN1117_data_out(1);
    CN115_sign_in(20) <= VN1117_sign_out(1);
    CN115_data_in(21) <= VN1205_data_out(1);
    CN115_sign_in(21) <= VN1205_sign_out(1);
    CN115_data_in(22) <= VN1222_data_out(1);
    CN115_sign_in(22) <= VN1222_sign_out(1);
    CN115_data_in(23) <= VN1255_data_out(1);
    CN115_sign_in(23) <= VN1255_sign_out(1);
    CN115_data_in(24) <= VN1380_data_out(1);
    CN115_sign_in(24) <= VN1380_sign_out(1);
    CN115_data_in(25) <= VN1420_data_out(1);
    CN115_sign_in(25) <= VN1420_sign_out(1);
    CN115_data_in(26) <= VN1469_data_out(1);
    CN115_sign_in(26) <= VN1469_sign_out(1);
    CN115_data_in(27) <= VN1530_data_out(1);
    CN115_sign_in(27) <= VN1530_sign_out(1);
    CN115_data_in(28) <= VN1605_data_out(1);
    CN115_sign_in(28) <= VN1605_sign_out(1);
    CN115_data_in(29) <= VN1639_data_out(1);
    CN115_sign_in(29) <= VN1639_sign_out(1);
    CN115_data_in(30) <= VN1654_data_out(1);
    CN115_sign_in(30) <= VN1654_sign_out(1);
    CN115_data_in(31) <= VN1754_data_out(1);
    CN115_sign_in(31) <= VN1754_sign_out(1);
    CN116_data_in(0) <= VN71_data_out(1);
    CN116_sign_in(0) <= VN71_sign_out(1);
    CN116_data_in(1) <= VN163_data_out(1);
    CN116_sign_in(1) <= VN163_sign_out(1);
    CN116_data_in(2) <= VN187_data_out(1);
    CN116_sign_in(2) <= VN187_sign_out(1);
    CN116_data_in(3) <= VN228_data_out(1);
    CN116_sign_in(3) <= VN228_sign_out(1);
    CN116_data_in(4) <= VN304_data_out(1);
    CN116_sign_in(4) <= VN304_sign_out(1);
    CN116_data_in(5) <= VN390_data_out(1);
    CN116_sign_in(5) <= VN390_sign_out(1);
    CN116_data_in(6) <= VN437_data_out(1);
    CN116_sign_in(6) <= VN437_sign_out(1);
    CN116_data_in(7) <= VN483_data_out(1);
    CN116_sign_in(7) <= VN483_sign_out(1);
    CN116_data_in(8) <= VN514_data_out(1);
    CN116_sign_in(8) <= VN514_sign_out(1);
    CN116_data_in(9) <= VN599_data_out(1);
    CN116_sign_in(9) <= VN599_sign_out(1);
    CN116_data_in(10) <= VN620_data_out(1);
    CN116_sign_in(10) <= VN620_sign_out(1);
    CN116_data_in(11) <= VN709_data_out(1);
    CN116_sign_in(11) <= VN709_sign_out(1);
    CN116_data_in(12) <= VN749_data_out(1);
    CN116_sign_in(12) <= VN749_sign_out(1);
    CN116_data_in(13) <= VN817_data_out(1);
    CN116_sign_in(13) <= VN817_sign_out(1);
    CN116_data_in(14) <= VN905_data_out(1);
    CN116_sign_in(14) <= VN905_sign_out(1);
    CN116_data_in(15) <= VN974_data_out(1);
    CN116_sign_in(15) <= VN974_sign_out(1);
    CN116_data_in(16) <= VN1037_data_out(1);
    CN116_sign_in(16) <= VN1037_sign_out(1);
    CN116_data_in(17) <= VN1067_data_out(1);
    CN116_sign_in(17) <= VN1067_sign_out(1);
    CN116_data_in(18) <= VN1160_data_out(1);
    CN116_sign_in(18) <= VN1160_sign_out(1);
    CN116_data_in(19) <= VN1196_data_out(1);
    CN116_sign_in(19) <= VN1196_sign_out(1);
    CN116_data_in(20) <= VN1224_data_out(1);
    CN116_sign_in(20) <= VN1224_sign_out(1);
    CN116_data_in(21) <= VN1226_data_out(1);
    CN116_sign_in(21) <= VN1226_sign_out(1);
    CN116_data_in(22) <= VN1347_data_out(1);
    CN116_sign_in(22) <= VN1347_sign_out(1);
    CN116_data_in(23) <= VN1386_data_out(1);
    CN116_sign_in(23) <= VN1386_sign_out(1);
    CN116_data_in(24) <= VN1542_data_out(1);
    CN116_sign_in(24) <= VN1542_sign_out(1);
    CN116_data_in(25) <= VN1632_data_out(1);
    CN116_sign_in(25) <= VN1632_sign_out(1);
    CN116_data_in(26) <= VN1662_data_out(1);
    CN116_sign_in(26) <= VN1662_sign_out(1);
    CN116_data_in(27) <= VN1785_data_out(1);
    CN116_sign_in(27) <= VN1785_sign_out(1);
    CN116_data_in(28) <= VN1947_data_out(1);
    CN116_sign_in(28) <= VN1947_sign_out(1);
    CN116_data_in(29) <= VN1998_data_out(1);
    CN116_sign_in(29) <= VN1998_sign_out(1);
    CN116_data_in(30) <= VN2024_data_out(1);
    CN116_sign_in(30) <= VN2024_sign_out(1);
    CN116_data_in(31) <= VN2035_data_out(1);
    CN116_sign_in(31) <= VN2035_sign_out(1);
    CN117_data_in(0) <= VN3_data_out(1);
    CN117_sign_in(0) <= VN3_sign_out(1);
    CN117_data_in(1) <= VN55_data_out(1);
    CN117_sign_in(1) <= VN55_sign_out(1);
    CN117_data_in(2) <= VN111_data_out(1);
    CN117_sign_in(2) <= VN111_sign_out(1);
    CN117_data_in(3) <= VN196_data_out(1);
    CN117_sign_in(3) <= VN196_sign_out(1);
    CN117_data_in(4) <= VN426_data_out(1);
    CN117_sign_in(4) <= VN426_sign_out(1);
    CN117_data_in(5) <= VN455_data_out(1);
    CN117_sign_in(5) <= VN455_sign_out(1);
    CN117_data_in(6) <= VN533_data_out(1);
    CN117_sign_in(6) <= VN533_sign_out(1);
    CN117_data_in(7) <= VN648_data_out(1);
    CN117_sign_in(7) <= VN648_sign_out(1);
    CN117_data_in(8) <= VN679_data_out(1);
    CN117_sign_in(8) <= VN679_sign_out(1);
    CN117_data_in(9) <= VN841_data_out(1);
    CN117_sign_in(9) <= VN841_sign_out(1);
    CN117_data_in(10) <= VN930_data_out(1);
    CN117_sign_in(10) <= VN930_sign_out(1);
    CN117_data_in(11) <= VN981_data_out(1);
    CN117_sign_in(11) <= VN981_sign_out(1);
    CN117_data_in(12) <= VN1016_data_out(1);
    CN117_sign_in(12) <= VN1016_sign_out(1);
    CN117_data_in(13) <= VN1093_data_out(1);
    CN117_sign_in(13) <= VN1093_sign_out(1);
    CN117_data_in(14) <= VN1135_data_out(1);
    CN117_sign_in(14) <= VN1135_sign_out(1);
    CN117_data_in(15) <= VN1185_data_out(1);
    CN117_sign_in(15) <= VN1185_sign_out(1);
    CN117_data_in(16) <= VN1273_data_out(1);
    CN117_sign_in(16) <= VN1273_sign_out(1);
    CN117_data_in(17) <= VN1325_data_out(1);
    CN117_sign_in(17) <= VN1325_sign_out(1);
    CN117_data_in(18) <= VN1345_data_out(1);
    CN117_sign_in(18) <= VN1345_sign_out(1);
    CN117_data_in(19) <= VN1449_data_out(1);
    CN117_sign_in(19) <= VN1449_sign_out(1);
    CN117_data_in(20) <= VN1537_data_out(1);
    CN117_sign_in(20) <= VN1537_sign_out(1);
    CN117_data_in(21) <= VN1576_data_out(1);
    CN117_sign_in(21) <= VN1576_sign_out(1);
    CN117_data_in(22) <= VN1657_data_out(1);
    CN117_sign_in(22) <= VN1657_sign_out(1);
    CN117_data_in(23) <= VN1701_data_out(1);
    CN117_sign_in(23) <= VN1701_sign_out(1);
    CN117_data_in(24) <= VN1808_data_out(1);
    CN117_sign_in(24) <= VN1808_sign_out(1);
    CN117_data_in(25) <= VN1864_data_out(1);
    CN117_sign_in(25) <= VN1864_sign_out(1);
    CN117_data_in(26) <= VN1877_data_out(1);
    CN117_sign_in(26) <= VN1877_sign_out(1);
    CN117_data_in(27) <= VN1913_data_out(1);
    CN117_sign_in(27) <= VN1913_sign_out(1);
    CN117_data_in(28) <= VN1931_data_out(1);
    CN117_sign_in(28) <= VN1931_sign_out(1);
    CN117_data_in(29) <= VN1934_data_out(1);
    CN117_sign_in(29) <= VN1934_sign_out(1);
    CN117_data_in(30) <= VN1965_data_out(1);
    CN117_sign_in(30) <= VN1965_sign_out(1);
    CN117_data_in(31) <= VN1974_data_out(1);
    CN117_sign_in(31) <= VN1974_sign_out(1);
    CN118_data_in(0) <= VN2_data_out(1);
    CN118_sign_in(0) <= VN2_sign_out(1);
    CN118_data_in(1) <= VN89_data_out(1);
    CN118_sign_in(1) <= VN89_sign_out(1);
    CN118_data_in(2) <= VN152_data_out(1);
    CN118_sign_in(2) <= VN152_sign_out(1);
    CN118_data_in(3) <= VN249_data_out(1);
    CN118_sign_in(3) <= VN249_sign_out(1);
    CN118_data_in(4) <= VN282_data_out(1);
    CN118_sign_in(4) <= VN282_sign_out(1);
    CN118_data_in(5) <= VN359_data_out(1);
    CN118_sign_in(5) <= VN359_sign_out(1);
    CN118_data_in(6) <= VN406_data_out(1);
    CN118_sign_in(6) <= VN406_sign_out(1);
    CN118_data_in(7) <= VN499_data_out(1);
    CN118_sign_in(7) <= VN499_sign_out(1);
    CN118_data_in(8) <= VN506_data_out(1);
    CN118_sign_in(8) <= VN506_sign_out(1);
    CN118_data_in(9) <= VN594_data_out(1);
    CN118_sign_in(9) <= VN594_sign_out(1);
    CN118_data_in(10) <= VN645_data_out(1);
    CN118_sign_in(10) <= VN645_sign_out(1);
    CN118_data_in(11) <= VN803_data_out(1);
    CN118_sign_in(11) <= VN803_sign_out(1);
    CN118_data_in(12) <= VN833_data_out(1);
    CN118_sign_in(12) <= VN833_sign_out(1);
    CN118_data_in(13) <= VN945_data_out(1);
    CN118_sign_in(13) <= VN945_sign_out(1);
    CN118_data_in(14) <= VN1053_data_out(1);
    CN118_sign_in(14) <= VN1053_sign_out(1);
    CN118_data_in(15) <= VN1106_data_out(1);
    CN118_sign_in(15) <= VN1106_sign_out(1);
    CN118_data_in(16) <= VN1156_data_out(1);
    CN118_sign_in(16) <= VN1156_sign_out(1);
    CN118_data_in(17) <= VN1201_data_out(1);
    CN118_sign_in(17) <= VN1201_sign_out(1);
    CN118_data_in(18) <= VN1259_data_out(1);
    CN118_sign_in(18) <= VN1259_sign_out(1);
    CN118_data_in(19) <= VN1281_data_out(1);
    CN118_sign_in(19) <= VN1281_sign_out(1);
    CN118_data_in(20) <= VN1378_data_out(1);
    CN118_sign_in(20) <= VN1378_sign_out(1);
    CN118_data_in(21) <= VN1403_data_out(1);
    CN118_sign_in(21) <= VN1403_sign_out(1);
    CN118_data_in(22) <= VN1433_data_out(1);
    CN118_sign_in(22) <= VN1433_sign_out(1);
    CN118_data_in(23) <= VN1492_data_out(1);
    CN118_sign_in(23) <= VN1492_sign_out(1);
    CN118_data_in(24) <= VN1531_data_out(1);
    CN118_sign_in(24) <= VN1531_sign_out(1);
    CN118_data_in(25) <= VN1599_data_out(1);
    CN118_sign_in(25) <= VN1599_sign_out(1);
    CN118_data_in(26) <= VN1660_data_out(1);
    CN118_sign_in(26) <= VN1660_sign_out(1);
    CN118_data_in(27) <= VN1711_data_out(1);
    CN118_sign_in(27) <= VN1711_sign_out(1);
    CN118_data_in(28) <= VN1873_data_out(1);
    CN118_sign_in(28) <= VN1873_sign_out(1);
    CN118_data_in(29) <= VN1924_data_out(1);
    CN118_sign_in(29) <= VN1924_sign_out(1);
    CN118_data_in(30) <= VN1984_data_out(1);
    CN118_sign_in(30) <= VN1984_sign_out(1);
    CN118_data_in(31) <= VN1985_data_out(1);
    CN118_sign_in(31) <= VN1985_sign_out(1);
    CN119_data_in(0) <= VN1_data_out(1);
    CN119_sign_in(0) <= VN1_sign_out(1);
    CN119_data_in(1) <= VN107_data_out(1);
    CN119_sign_in(1) <= VN107_sign_out(1);
    CN119_data_in(2) <= VN154_data_out(1);
    CN119_sign_in(2) <= VN154_sign_out(1);
    CN119_data_in(3) <= VN227_data_out(1);
    CN119_sign_in(3) <= VN227_sign_out(1);
    CN119_data_in(4) <= VN319_data_out(1);
    CN119_sign_in(4) <= VN319_sign_out(1);
    CN119_data_in(5) <= VN445_data_out(1);
    CN119_sign_in(5) <= VN445_sign_out(1);
    CN119_data_in(6) <= VN546_data_out(1);
    CN119_sign_in(6) <= VN546_sign_out(1);
    CN119_data_in(7) <= VN604_data_out(1);
    CN119_sign_in(7) <= VN604_sign_out(1);
    CN119_data_in(8) <= VN659_data_out(1);
    CN119_sign_in(8) <= VN659_sign_out(1);
    CN119_data_in(9) <= VN727_data_out(1);
    CN119_sign_in(9) <= VN727_sign_out(1);
    CN119_data_in(10) <= VN784_data_out(1);
    CN119_sign_in(10) <= VN784_sign_out(1);
    CN119_data_in(11) <= VN851_data_out(1);
    CN119_sign_in(11) <= VN851_sign_out(1);
    CN119_data_in(12) <= VN1002_data_out(1);
    CN119_sign_in(12) <= VN1002_sign_out(1);
    CN119_data_in(13) <= VN1056_data_out(1);
    CN119_sign_in(13) <= VN1056_sign_out(1);
    CN119_data_in(14) <= VN1081_data_out(1);
    CN119_sign_in(14) <= VN1081_sign_out(1);
    CN119_data_in(15) <= VN1126_data_out(1);
    CN119_sign_in(15) <= VN1126_sign_out(1);
    CN119_data_in(16) <= VN1306_data_out(1);
    CN119_sign_in(16) <= VN1306_sign_out(1);
    CN119_data_in(17) <= VN1359_data_out(1);
    CN119_sign_in(17) <= VN1359_sign_out(1);
    CN119_data_in(18) <= VN1413_data_out(1);
    CN119_sign_in(18) <= VN1413_sign_out(1);
    CN119_data_in(19) <= VN1427_data_out(1);
    CN119_sign_in(19) <= VN1427_sign_out(1);
    CN119_data_in(20) <= VN1464_data_out(1);
    CN119_sign_in(20) <= VN1464_sign_out(1);
    CN119_data_in(21) <= VN1522_data_out(1);
    CN119_sign_in(21) <= VN1522_sign_out(1);
    CN119_data_in(22) <= VN1648_data_out(1);
    CN119_sign_in(22) <= VN1648_sign_out(1);
    CN119_data_in(23) <= VN1688_data_out(1);
    CN119_sign_in(23) <= VN1688_sign_out(1);
    CN119_data_in(24) <= VN1800_data_out(1);
    CN119_sign_in(24) <= VN1800_sign_out(1);
    CN119_data_in(25) <= VN1879_data_out(1);
    CN119_sign_in(25) <= VN1879_sign_out(1);
    CN119_data_in(26) <= VN1941_data_out(1);
    CN119_sign_in(26) <= VN1941_sign_out(1);
    CN119_data_in(27) <= VN1942_data_out(1);
    CN119_sign_in(27) <= VN1942_sign_out(1);
    CN119_data_in(28) <= VN1945_data_out(1);
    CN119_sign_in(28) <= VN1945_sign_out(1);
    CN119_data_in(29) <= VN1955_data_out(1);
    CN119_sign_in(29) <= VN1955_sign_out(1);
    CN119_data_in(30) <= VN1969_data_out(1);
    CN119_sign_in(30) <= VN1969_sign_out(1);
    CN119_data_in(31) <= VN1975_data_out(1);
    CN119_sign_in(31) <= VN1975_sign_out(1);
    CN120_data_in(0) <= VN0_data_out(1);
    CN120_sign_in(0) <= VN0_sign_out(1);
    CN120_data_in(1) <= VN80_data_out(1);
    CN120_sign_in(1) <= VN80_sign_out(1);
    CN120_data_in(2) <= VN321_data_out(1);
    CN120_sign_in(2) <= VN321_sign_out(1);
    CN120_data_in(3) <= VN360_data_out(1);
    CN120_sign_in(3) <= VN360_sign_out(1);
    CN120_data_in(4) <= VN401_data_out(1);
    CN120_sign_in(4) <= VN401_sign_out(1);
    CN120_data_in(5) <= VN502_data_out(1);
    CN120_sign_in(5) <= VN502_sign_out(1);
    CN120_data_in(6) <= VN515_data_out(1);
    CN120_sign_in(6) <= VN515_sign_out(1);
    CN120_data_in(7) <= VN653_data_out(1);
    CN120_sign_in(7) <= VN653_sign_out(1);
    CN120_data_in(8) <= VN745_data_out(1);
    CN120_sign_in(8) <= VN745_sign_out(1);
    CN120_data_in(9) <= VN805_data_out(1);
    CN120_sign_in(9) <= VN805_sign_out(1);
    CN120_data_in(10) <= VN855_data_out(1);
    CN120_sign_in(10) <= VN855_sign_out(1);
    CN120_data_in(11) <= VN980_data_out(1);
    CN120_sign_in(11) <= VN980_sign_out(1);
    CN120_data_in(12) <= VN1040_data_out(1);
    CN120_sign_in(12) <= VN1040_sign_out(1);
    CN120_data_in(13) <= VN1061_data_out(1);
    CN120_sign_in(13) <= VN1061_sign_out(1);
    CN120_data_in(14) <= VN1252_data_out(1);
    CN120_sign_in(14) <= VN1252_sign_out(1);
    CN120_data_in(15) <= VN1320_data_out(1);
    CN120_sign_in(15) <= VN1320_sign_out(1);
    CN120_data_in(16) <= VN1362_data_out(1);
    CN120_sign_in(16) <= VN1362_sign_out(1);
    CN120_data_in(17) <= VN1407_data_out(1);
    CN120_sign_in(17) <= VN1407_sign_out(1);
    CN120_data_in(18) <= VN1491_data_out(1);
    CN120_sign_in(18) <= VN1491_sign_out(1);
    CN120_data_in(19) <= VN1562_data_out(1);
    CN120_sign_in(19) <= VN1562_sign_out(1);
    CN120_data_in(20) <= VN1589_data_out(1);
    CN120_sign_in(20) <= VN1589_sign_out(1);
    CN120_data_in(21) <= VN1716_data_out(1);
    CN120_sign_in(21) <= VN1716_sign_out(1);
    CN120_data_in(22) <= VN1726_data_out(1);
    CN120_sign_in(22) <= VN1726_sign_out(1);
    CN120_data_in(23) <= VN1780_data_out(1);
    CN120_sign_in(23) <= VN1780_sign_out(1);
    CN120_data_in(24) <= VN1790_data_out(1);
    CN120_sign_in(24) <= VN1790_sign_out(1);
    CN120_data_in(25) <= VN1852_data_out(1);
    CN120_sign_in(25) <= VN1852_sign_out(1);
    CN120_data_in(26) <= VN1862_data_out(1);
    CN120_sign_in(26) <= VN1862_sign_out(1);
    CN120_data_in(27) <= VN1899_data_out(1);
    CN120_sign_in(27) <= VN1899_sign_out(1);
    CN120_data_in(28) <= VN1904_data_out(1);
    CN120_sign_in(28) <= VN1904_sign_out(1);
    CN120_data_in(29) <= VN1958_data_out(1);
    CN120_sign_in(29) <= VN1958_sign_out(1);
    CN120_data_in(30) <= VN2006_data_out(1);
    CN120_sign_in(30) <= VN2006_sign_out(1);
    CN120_data_in(31) <= VN2009_data_out(1);
    CN120_sign_in(31) <= VN2009_sign_out(1);
    CN121_data_in(0) <= VN64_data_out(1);
    CN121_sign_in(0) <= VN64_sign_out(1);
    CN121_data_in(1) <= VN161_data_out(1);
    CN121_sign_in(1) <= VN161_sign_out(1);
    CN121_data_in(2) <= VN217_data_out(1);
    CN121_sign_in(2) <= VN217_sign_out(1);
    CN121_data_in(3) <= VN236_data_out(1);
    CN121_sign_in(3) <= VN236_sign_out(1);
    CN121_data_in(4) <= VN291_data_out(1);
    CN121_sign_in(4) <= VN291_sign_out(1);
    CN121_data_in(5) <= VN350_data_out(1);
    CN121_sign_in(5) <= VN350_sign_out(1);
    CN121_data_in(6) <= VN411_data_out(1);
    CN121_sign_in(6) <= VN411_sign_out(1);
    CN121_data_in(7) <= VN466_data_out(1);
    CN121_sign_in(7) <= VN466_sign_out(1);
    CN121_data_in(8) <= VN566_data_out(1);
    CN121_sign_in(8) <= VN566_sign_out(1);
    CN121_data_in(9) <= VN628_data_out(1);
    CN121_sign_in(9) <= VN628_sign_out(1);
    CN121_data_in(10) <= VN670_data_out(1);
    CN121_sign_in(10) <= VN670_sign_out(1);
    CN121_data_in(11) <= VN767_data_out(1);
    CN121_sign_in(11) <= VN767_sign_out(1);
    CN121_data_in(12) <= VN819_data_out(1);
    CN121_sign_in(12) <= VN819_sign_out(1);
    CN121_data_in(13) <= VN901_data_out(1);
    CN121_sign_in(13) <= VN901_sign_out(1);
    CN121_data_in(14) <= VN959_data_out(1);
    CN121_sign_in(14) <= VN959_sign_out(1);
    CN121_data_in(15) <= VN1017_data_out(1);
    CN121_sign_in(15) <= VN1017_sign_out(1);
    CN121_data_in(16) <= VN1083_data_out(1);
    CN121_sign_in(16) <= VN1083_sign_out(1);
    CN121_data_in(17) <= VN1137_data_out(1);
    CN121_sign_in(17) <= VN1137_sign_out(1);
    CN121_data_in(18) <= VN1189_data_out(1);
    CN121_sign_in(18) <= VN1189_sign_out(1);
    CN121_data_in(19) <= VN1223_data_out(1);
    CN121_sign_in(19) <= VN1223_sign_out(1);
    CN121_data_in(20) <= VN1249_data_out(1);
    CN121_sign_in(20) <= VN1249_sign_out(1);
    CN121_data_in(21) <= VN1296_data_out(1);
    CN121_sign_in(21) <= VN1296_sign_out(1);
    CN121_data_in(22) <= VN1348_data_out(1);
    CN121_sign_in(22) <= VN1348_sign_out(1);
    CN121_data_in(23) <= VN1411_data_out(1);
    CN121_sign_in(23) <= VN1411_sign_out(1);
    CN121_data_in(24) <= VN1479_data_out(1);
    CN121_sign_in(24) <= VN1479_sign_out(1);
    CN121_data_in(25) <= VN1501_data_out(1);
    CN121_sign_in(25) <= VN1501_sign_out(1);
    CN121_data_in(26) <= VN1572_data_out(1);
    CN121_sign_in(26) <= VN1572_sign_out(1);
    CN121_data_in(27) <= VN1646_data_out(1);
    CN121_sign_in(27) <= VN1646_sign_out(1);
    CN121_data_in(28) <= VN1696_data_out(1);
    CN121_sign_in(28) <= VN1696_sign_out(1);
    CN121_data_in(29) <= VN1723_data_out(1);
    CN121_sign_in(29) <= VN1723_sign_out(1);
    CN121_data_in(30) <= VN1766_data_out(1);
    CN121_sign_in(30) <= VN1766_sign_out(1);
    CN121_data_in(31) <= VN1829_data_out(1);
    CN121_sign_in(31) <= VN1829_sign_out(1);
    CN122_data_in(0) <= VN91_data_out(1);
    CN122_sign_in(0) <= VN91_sign_out(1);
    CN122_data_in(1) <= VN114_data_out(1);
    CN122_sign_in(1) <= VN114_sign_out(1);
    CN122_data_in(2) <= VN201_data_out(1);
    CN122_sign_in(2) <= VN201_sign_out(1);
    CN122_data_in(3) <= VN241_data_out(1);
    CN122_sign_in(3) <= VN241_sign_out(1);
    CN122_data_in(4) <= VN327_data_out(1);
    CN122_sign_in(4) <= VN327_sign_out(1);
    CN122_data_in(5) <= VN375_data_out(1);
    CN122_sign_in(5) <= VN375_sign_out(1);
    CN122_data_in(6) <= VN475_data_out(1);
    CN122_sign_in(6) <= VN475_sign_out(1);
    CN122_data_in(7) <= VN551_data_out(1);
    CN122_sign_in(7) <= VN551_sign_out(1);
    CN122_data_in(8) <= VN607_data_out(1);
    CN122_sign_in(8) <= VN607_sign_out(1);
    CN122_data_in(9) <= VN637_data_out(1);
    CN122_sign_in(9) <= VN637_sign_out(1);
    CN122_data_in(10) <= VN686_data_out(1);
    CN122_sign_in(10) <= VN686_sign_out(1);
    CN122_data_in(11) <= VN768_data_out(1);
    CN122_sign_in(11) <= VN768_sign_out(1);
    CN122_data_in(12) <= VN815_data_out(1);
    CN122_sign_in(12) <= VN815_sign_out(1);
    CN122_data_in(13) <= VN898_data_out(1);
    CN122_sign_in(13) <= VN898_sign_out(1);
    CN122_data_in(14) <= VN962_data_out(1);
    CN122_sign_in(14) <= VN962_sign_out(1);
    CN122_data_in(15) <= VN1036_data_out(1);
    CN122_sign_in(15) <= VN1036_sign_out(1);
    CN122_data_in(16) <= VN1128_data_out(1);
    CN122_sign_in(16) <= VN1128_sign_out(1);
    CN122_data_in(17) <= VN1182_data_out(1);
    CN122_sign_in(17) <= VN1182_sign_out(1);
    CN122_data_in(18) <= VN1264_data_out(1);
    CN122_sign_in(18) <= VN1264_sign_out(1);
    CN122_data_in(19) <= VN1328_data_out(1);
    CN122_sign_in(19) <= VN1328_sign_out(1);
    CN122_data_in(20) <= VN1379_data_out(1);
    CN122_sign_in(20) <= VN1379_sign_out(1);
    CN122_data_in(21) <= VN1400_data_out(1);
    CN122_sign_in(21) <= VN1400_sign_out(1);
    CN122_data_in(22) <= VN1565_data_out(1);
    CN122_sign_in(22) <= VN1565_sign_out(1);
    CN122_data_in(23) <= VN1673_data_out(1);
    CN122_sign_in(23) <= VN1673_sign_out(1);
    CN122_data_in(24) <= VN1760_data_out(1);
    CN122_sign_in(24) <= VN1760_sign_out(1);
    CN122_data_in(25) <= VN1771_data_out(1);
    CN122_sign_in(25) <= VN1771_sign_out(1);
    CN122_data_in(26) <= VN1774_data_out(1);
    CN122_sign_in(26) <= VN1774_sign_out(1);
    CN122_data_in(27) <= VN1789_data_out(1);
    CN122_sign_in(27) <= VN1789_sign_out(1);
    CN122_data_in(28) <= VN1865_data_out(1);
    CN122_sign_in(28) <= VN1865_sign_out(1);
    CN122_data_in(29) <= VN1928_data_out(1);
    CN122_sign_in(29) <= VN1928_sign_out(1);
    CN122_data_in(30) <= VN1990_data_out(1);
    CN122_sign_in(30) <= VN1990_sign_out(1);
    CN122_data_in(31) <= VN1991_data_out(1);
    CN122_sign_in(31) <= VN1991_sign_out(1);
    CN123_data_in(0) <= VN82_data_out(1);
    CN123_sign_in(0) <= VN82_sign_out(1);
    CN123_data_in(1) <= VN122_data_out(1);
    CN123_sign_in(1) <= VN122_sign_out(1);
    CN123_data_in(2) <= VN213_data_out(1);
    CN123_sign_in(2) <= VN213_sign_out(1);
    CN123_data_in(3) <= VN279_data_out(1);
    CN123_sign_in(3) <= VN279_sign_out(1);
    CN123_data_in(4) <= VN382_data_out(1);
    CN123_sign_in(4) <= VN382_sign_out(1);
    CN123_data_in(5) <= VN428_data_out(1);
    CN123_sign_in(5) <= VN428_sign_out(1);
    CN123_data_in(6) <= VN470_data_out(1);
    CN123_sign_in(6) <= VN470_sign_out(1);
    CN123_data_in(7) <= VN512_data_out(1);
    CN123_sign_in(7) <= VN512_sign_out(1);
    CN123_data_in(8) <= VN569_data_out(1);
    CN123_sign_in(8) <= VN569_sign_out(1);
    CN123_data_in(9) <= VN630_data_out(1);
    CN123_sign_in(9) <= VN630_sign_out(1);
    CN123_data_in(10) <= VN716_data_out(1);
    CN123_sign_in(10) <= VN716_sign_out(1);
    CN123_data_in(11) <= VN849_data_out(1);
    CN123_sign_in(11) <= VN849_sign_out(1);
    CN123_data_in(12) <= VN914_data_out(1);
    CN123_sign_in(12) <= VN914_sign_out(1);
    CN123_data_in(13) <= VN946_data_out(1);
    CN123_sign_in(13) <= VN946_sign_out(1);
    CN123_data_in(14) <= VN1008_data_out(1);
    CN123_sign_in(14) <= VN1008_sign_out(1);
    CN123_data_in(15) <= VN1091_data_out(1);
    CN123_sign_in(15) <= VN1091_sign_out(1);
    CN123_data_in(16) <= VN1110_data_out(1);
    CN123_sign_in(16) <= VN1110_sign_out(1);
    CN123_data_in(17) <= VN1115_data_out(1);
    CN123_sign_in(17) <= VN1115_sign_out(1);
    CN123_data_in(18) <= VN1297_data_out(1);
    CN123_sign_in(18) <= VN1297_sign_out(1);
    CN123_data_in(19) <= VN1344_data_out(1);
    CN123_sign_in(19) <= VN1344_sign_out(1);
    CN123_data_in(20) <= VN1543_data_out(1);
    CN123_sign_in(20) <= VN1543_sign_out(1);
    CN123_data_in(21) <= VN1569_data_out(1);
    CN123_sign_in(21) <= VN1569_sign_out(1);
    CN123_data_in(22) <= VN1600_data_out(1);
    CN123_sign_in(22) <= VN1600_sign_out(1);
    CN123_data_in(23) <= VN1636_data_out(1);
    CN123_sign_in(23) <= VN1636_sign_out(1);
    CN123_data_in(24) <= VN1682_data_out(1);
    CN123_sign_in(24) <= VN1682_sign_out(1);
    CN123_data_in(25) <= VN1722_data_out(1);
    CN123_sign_in(25) <= VN1722_sign_out(1);
    CN123_data_in(26) <= VN1814_data_out(1);
    CN123_sign_in(26) <= VN1814_sign_out(1);
    CN123_data_in(27) <= VN1838_data_out(1);
    CN123_sign_in(27) <= VN1838_sign_out(1);
    CN123_data_in(28) <= VN1868_data_out(1);
    CN123_sign_in(28) <= VN1868_sign_out(1);
    CN123_data_in(29) <= VN1876_data_out(1);
    CN123_sign_in(29) <= VN1876_sign_out(1);
    CN123_data_in(30) <= VN1987_data_out(1);
    CN123_sign_in(30) <= VN1987_sign_out(1);
    CN123_data_in(31) <= VN1988_data_out(1);
    CN123_sign_in(31) <= VN1988_sign_out(1);
    CN124_data_in(0) <= VN69_data_out(1);
    CN124_sign_in(0) <= VN69_sign_out(1);
    CN124_data_in(1) <= VN153_data_out(1);
    CN124_sign_in(1) <= VN153_sign_out(1);
    CN124_data_in(2) <= VN240_data_out(1);
    CN124_sign_in(2) <= VN240_sign_out(1);
    CN124_data_in(3) <= VN292_data_out(1);
    CN124_sign_in(3) <= VN292_sign_out(1);
    CN124_data_in(4) <= VN364_data_out(1);
    CN124_sign_in(4) <= VN364_sign_out(1);
    CN124_data_in(5) <= VN414_data_out(1);
    CN124_sign_in(5) <= VN414_sign_out(1);
    CN124_data_in(6) <= VN476_data_out(1);
    CN124_sign_in(6) <= VN476_sign_out(1);
    CN124_data_in(7) <= VN542_data_out(1);
    CN124_sign_in(7) <= VN542_sign_out(1);
    CN124_data_in(8) <= VN634_data_out(1);
    CN124_sign_in(8) <= VN634_sign_out(1);
    CN124_data_in(9) <= VN886_data_out(1);
    CN124_sign_in(9) <= VN886_sign_out(1);
    CN124_data_in(10) <= VN907_data_out(1);
    CN124_sign_in(10) <= VN907_sign_out(1);
    CN124_data_in(11) <= VN1049_data_out(1);
    CN124_sign_in(11) <= VN1049_sign_out(1);
    CN124_data_in(12) <= VN1109_data_out(1);
    CN124_sign_in(12) <= VN1109_sign_out(1);
    CN124_data_in(13) <= VN1133_data_out(1);
    CN124_sign_in(13) <= VN1133_sign_out(1);
    CN124_data_in(14) <= VN1234_data_out(1);
    CN124_sign_in(14) <= VN1234_sign_out(1);
    CN124_data_in(15) <= VN1308_data_out(1);
    CN124_sign_in(15) <= VN1308_sign_out(1);
    CN124_data_in(16) <= VN1370_data_out(1);
    CN124_sign_in(16) <= VN1370_sign_out(1);
    CN124_data_in(17) <= VN1419_data_out(1);
    CN124_sign_in(17) <= VN1419_sign_out(1);
    CN124_data_in(18) <= VN1457_data_out(1);
    CN124_sign_in(18) <= VN1457_sign_out(1);
    CN124_data_in(19) <= VN1597_data_out(1);
    CN124_sign_in(19) <= VN1597_sign_out(1);
    CN124_data_in(20) <= VN1608_data_out(1);
    CN124_sign_in(20) <= VN1608_sign_out(1);
    CN124_data_in(21) <= VN1721_data_out(1);
    CN124_sign_in(21) <= VN1721_sign_out(1);
    CN124_data_in(22) <= VN1795_data_out(1);
    CN124_sign_in(22) <= VN1795_sign_out(1);
    CN124_data_in(23) <= VN1821_data_out(1);
    CN124_sign_in(23) <= VN1821_sign_out(1);
    CN124_data_in(24) <= VN1843_data_out(1);
    CN124_sign_in(24) <= VN1843_sign_out(1);
    CN124_data_in(25) <= VN1856_data_out(1);
    CN124_sign_in(25) <= VN1856_sign_out(1);
    CN124_data_in(26) <= VN1898_data_out(1);
    CN124_sign_in(26) <= VN1898_sign_out(1);
    CN124_data_in(27) <= VN1910_data_out(1);
    CN124_sign_in(27) <= VN1910_sign_out(1);
    CN124_data_in(28) <= VN1932_data_out(1);
    CN124_sign_in(28) <= VN1932_sign_out(1);
    CN124_data_in(29) <= VN1962_data_out(1);
    CN124_sign_in(29) <= VN1962_sign_out(1);
    CN124_data_in(30) <= VN1970_data_out(1);
    CN124_sign_in(30) <= VN1970_sign_out(1);
    CN124_data_in(31) <= VN1976_data_out(1);
    CN124_sign_in(31) <= VN1976_sign_out(1);
    CN125_data_in(0) <= VN87_data_out(1);
    CN125_sign_in(0) <= VN87_sign_out(1);
    CN125_data_in(1) <= VN169_data_out(1);
    CN125_sign_in(1) <= VN169_sign_out(1);
    CN125_data_in(2) <= VN320_data_out(1);
    CN125_sign_in(2) <= VN320_sign_out(1);
    CN125_data_in(3) <= VN366_data_out(1);
    CN125_sign_in(3) <= VN366_sign_out(1);
    CN125_data_in(4) <= VN431_data_out(1);
    CN125_sign_in(4) <= VN431_sign_out(1);
    CN125_data_in(5) <= VN465_data_out(1);
    CN125_sign_in(5) <= VN465_sign_out(1);
    CN125_data_in(6) <= VN539_data_out(1);
    CN125_sign_in(6) <= VN539_sign_out(1);
    CN125_data_in(7) <= VN596_data_out(1);
    CN125_sign_in(7) <= VN596_sign_out(1);
    CN125_data_in(8) <= VN625_data_out(1);
    CN125_sign_in(8) <= VN625_sign_out(1);
    CN125_data_in(9) <= VN753_data_out(1);
    CN125_sign_in(9) <= VN753_sign_out(1);
    CN125_data_in(10) <= VN800_data_out(1);
    CN125_sign_in(10) <= VN800_sign_out(1);
    CN125_data_in(11) <= VN837_data_out(1);
    CN125_sign_in(11) <= VN837_sign_out(1);
    CN125_data_in(12) <= VN936_data_out(1);
    CN125_sign_in(12) <= VN936_sign_out(1);
    CN125_data_in(13) <= VN1001_data_out(1);
    CN125_sign_in(13) <= VN1001_sign_out(1);
    CN125_data_in(14) <= VN1019_data_out(1);
    CN125_sign_in(14) <= VN1019_sign_out(1);
    CN125_data_in(15) <= VN1078_data_out(1);
    CN125_sign_in(15) <= VN1078_sign_out(1);
    CN125_data_in(16) <= VN1113_data_out(1);
    CN125_sign_in(16) <= VN1113_sign_out(1);
    CN125_data_in(17) <= VN1304_data_out(1);
    CN125_sign_in(17) <= VN1304_sign_out(1);
    CN125_data_in(18) <= VN1356_data_out(1);
    CN125_sign_in(18) <= VN1356_sign_out(1);
    CN125_data_in(19) <= VN1434_data_out(1);
    CN125_sign_in(19) <= VN1434_sign_out(1);
    CN125_data_in(20) <= VN1493_data_out(1);
    CN125_sign_in(20) <= VN1493_sign_out(1);
    CN125_data_in(21) <= VN1510_data_out(1);
    CN125_sign_in(21) <= VN1510_sign_out(1);
    CN125_data_in(22) <= VN1539_data_out(1);
    CN125_sign_in(22) <= VN1539_sign_out(1);
    CN125_data_in(23) <= VN1692_data_out(1);
    CN125_sign_in(23) <= VN1692_sign_out(1);
    CN125_data_in(24) <= VN1719_data_out(1);
    CN125_sign_in(24) <= VN1719_sign_out(1);
    CN125_data_in(25) <= VN1738_data_out(1);
    CN125_sign_in(25) <= VN1738_sign_out(1);
    CN125_data_in(26) <= VN1784_data_out(1);
    CN125_sign_in(26) <= VN1784_sign_out(1);
    CN125_data_in(27) <= VN1816_data_out(1);
    CN125_sign_in(27) <= VN1816_sign_out(1);
    CN125_data_in(28) <= VN1859_data_out(1);
    CN125_sign_in(28) <= VN1859_sign_out(1);
    CN125_data_in(29) <= VN1896_data_out(1);
    CN125_sign_in(29) <= VN1896_sign_out(1);
    CN125_data_in(30) <= VN1959_data_out(1);
    CN125_sign_in(30) <= VN1959_sign_out(1);
    CN125_data_in(31) <= VN1964_data_out(1);
    CN125_sign_in(31) <= VN1964_sign_out(1);
    CN126_data_in(0) <= VN60_data_out(1);
    CN126_sign_in(0) <= VN60_sign_out(1);
    CN126_data_in(1) <= VN139_data_out(1);
    CN126_sign_in(1) <= VN139_sign_out(1);
    CN126_data_in(2) <= VN186_data_out(1);
    CN126_sign_in(2) <= VN186_sign_out(1);
    CN126_data_in(3) <= VN271_data_out(1);
    CN126_sign_in(3) <= VN271_sign_out(1);
    CN126_data_in(4) <= VN281_data_out(1);
    CN126_sign_in(4) <= VN281_sign_out(1);
    CN126_data_in(5) <= VN334_data_out(1);
    CN126_sign_in(5) <= VN334_sign_out(1);
    CN126_data_in(6) <= VN394_data_out(1);
    CN126_sign_in(6) <= VN394_sign_out(1);
    CN126_data_in(7) <= VN487_data_out(1);
    CN126_sign_in(7) <= VN487_sign_out(1);
    CN126_data_in(8) <= VN555_data_out(1);
    CN126_sign_in(8) <= VN555_sign_out(1);
    CN126_data_in(9) <= VN660_data_out(1);
    CN126_sign_in(9) <= VN660_sign_out(1);
    CN126_data_in(10) <= VN720_data_out(1);
    CN126_sign_in(10) <= VN720_sign_out(1);
    CN126_data_in(11) <= VN758_data_out(1);
    CN126_sign_in(11) <= VN758_sign_out(1);
    CN126_data_in(12) <= VN779_data_out(1);
    CN126_sign_in(12) <= VN779_sign_out(1);
    CN126_data_in(13) <= VN860_data_out(1);
    CN126_sign_in(13) <= VN860_sign_out(1);
    CN126_data_in(14) <= VN890_data_out(1);
    CN126_sign_in(14) <= VN890_sign_out(1);
    CN126_data_in(15) <= VN971_data_out(1);
    CN126_sign_in(15) <= VN971_sign_out(1);
    CN126_data_in(16) <= VN1010_data_out(1);
    CN126_sign_in(16) <= VN1010_sign_out(1);
    CN126_data_in(17) <= VN1079_data_out(1);
    CN126_sign_in(17) <= VN1079_sign_out(1);
    CN126_data_in(18) <= VN1162_data_out(1);
    CN126_sign_in(18) <= VN1162_sign_out(1);
    CN126_data_in(19) <= VN1237_data_out(1);
    CN126_sign_in(19) <= VN1237_sign_out(1);
    CN126_data_in(20) <= VN1276_data_out(1);
    CN126_sign_in(20) <= VN1276_sign_out(1);
    CN126_data_in(21) <= VN1323_data_out(1);
    CN126_sign_in(21) <= VN1323_sign_out(1);
    CN126_data_in(22) <= VN1334_data_out(1);
    CN126_sign_in(22) <= VN1334_sign_out(1);
    CN126_data_in(23) <= VN1381_data_out(1);
    CN126_sign_in(23) <= VN1381_sign_out(1);
    CN126_data_in(24) <= VN1515_data_out(1);
    CN126_sign_in(24) <= VN1515_sign_out(1);
    CN126_data_in(25) <= VN1549_data_out(1);
    CN126_sign_in(25) <= VN1549_sign_out(1);
    CN126_data_in(26) <= VN1586_data_out(1);
    CN126_sign_in(26) <= VN1586_sign_out(1);
    CN126_data_in(27) <= VN1635_data_out(1);
    CN126_sign_in(27) <= VN1635_sign_out(1);
    CN126_data_in(28) <= VN1720_data_out(1);
    CN126_sign_in(28) <= VN1720_sign_out(1);
    CN126_data_in(29) <= VN1757_data_out(1);
    CN126_sign_in(29) <= VN1757_sign_out(1);
    CN126_data_in(30) <= VN1764_data_out(1);
    CN126_sign_in(30) <= VN1764_sign_out(1);
    CN126_data_in(31) <= VN1830_data_out(1);
    CN126_sign_in(31) <= VN1830_sign_out(1);
    CN127_data_in(0) <= VN52_data_out(1);
    CN127_sign_in(0) <= VN52_sign_out(1);
    CN127_data_in(1) <= VN57_data_out(1);
    CN127_sign_in(1) <= VN57_sign_out(1);
    CN127_data_in(2) <= VN117_data_out(1);
    CN127_sign_in(2) <= VN117_sign_out(1);
    CN127_data_in(3) <= VN173_data_out(1);
    CN127_sign_in(3) <= VN173_sign_out(1);
    CN127_data_in(4) <= VN277_data_out(1);
    CN127_sign_in(4) <= VN277_sign_out(1);
    CN127_data_in(5) <= VN306_data_out(1);
    CN127_sign_in(5) <= VN306_sign_out(1);
    CN127_data_in(6) <= VN373_data_out(1);
    CN127_sign_in(6) <= VN373_sign_out(1);
    CN127_data_in(7) <= VN403_data_out(1);
    CN127_sign_in(7) <= VN403_sign_out(1);
    CN127_data_in(8) <= VN494_data_out(1);
    CN127_sign_in(8) <= VN494_sign_out(1);
    CN127_data_in(9) <= VN548_data_out(1);
    CN127_sign_in(9) <= VN548_sign_out(1);
    CN127_data_in(10) <= VN597_data_out(1);
    CN127_sign_in(10) <= VN597_sign_out(1);
    CN127_data_in(11) <= VN644_data_out(1);
    CN127_sign_in(11) <= VN644_sign_out(1);
    CN127_data_in(12) <= VN697_data_out(1);
    CN127_sign_in(12) <= VN697_sign_out(1);
    CN127_data_in(13) <= VN825_data_out(1);
    CN127_sign_in(13) <= VN825_sign_out(1);
    CN127_data_in(14) <= VN858_data_out(1);
    CN127_sign_in(14) <= VN858_sign_out(1);
    CN127_data_in(15) <= VN940_data_out(1);
    CN127_sign_in(15) <= VN940_sign_out(1);
    CN127_data_in(16) <= VN955_data_out(1);
    CN127_sign_in(16) <= VN955_sign_out(1);
    CN127_data_in(17) <= VN1054_data_out(1);
    CN127_sign_in(17) <= VN1054_sign_out(1);
    CN127_data_in(18) <= VN1120_data_out(1);
    CN127_sign_in(18) <= VN1120_sign_out(1);
    CN127_data_in(19) <= VN1210_data_out(1);
    CN127_sign_in(19) <= VN1210_sign_out(1);
    CN127_data_in(20) <= VN1221_data_out(1);
    CN127_sign_in(20) <= VN1221_sign_out(1);
    CN127_data_in(21) <= VN1240_data_out(1);
    CN127_sign_in(21) <= VN1240_sign_out(1);
    CN127_data_in(22) <= VN1292_data_out(1);
    CN127_sign_in(22) <= VN1292_sign_out(1);
    CN127_data_in(23) <= VN1372_data_out(1);
    CN127_sign_in(23) <= VN1372_sign_out(1);
    CN127_data_in(24) <= VN1414_data_out(1);
    CN127_sign_in(24) <= VN1414_sign_out(1);
    CN127_data_in(25) <= VN1430_data_out(1);
    CN127_sign_in(25) <= VN1430_sign_out(1);
    CN127_data_in(26) <= VN1499_data_out(1);
    CN127_sign_in(26) <= VN1499_sign_out(1);
    CN127_data_in(27) <= VN1506_data_out(1);
    CN127_sign_in(27) <= VN1506_sign_out(1);
    CN127_data_in(28) <= VN1587_data_out(1);
    CN127_sign_in(28) <= VN1587_sign_out(1);
    CN127_data_in(29) <= VN1618_data_out(1);
    CN127_sign_in(29) <= VN1618_sign_out(1);
    CN127_data_in(30) <= VN1706_data_out(1);
    CN127_sign_in(30) <= VN1706_sign_out(1);
    CN127_data_in(31) <= VN1755_data_out(1);
    CN127_sign_in(31) <= VN1755_sign_out(1);
    CN128_data_in(0) <= VN53_data_out(2);
    CN128_sign_in(0) <= VN53_sign_out(2);
    CN128_data_in(1) <= VN108_data_out(2);
    CN128_sign_in(1) <= VN108_sign_out(2);
    CN128_data_in(2) <= VN129_data_out(2);
    CN128_sign_in(2) <= VN129_sign_out(2);
    CN128_data_in(3) <= VN198_data_out(2);
    CN128_sign_in(3) <= VN198_sign_out(2);
    CN128_data_in(4) <= VN244_data_out(2);
    CN128_sign_in(4) <= VN244_sign_out(2);
    CN128_data_in(5) <= VN298_data_out(2);
    CN128_sign_in(5) <= VN298_sign_out(2);
    CN128_data_in(6) <= VN341_data_out(2);
    CN128_sign_in(6) <= VN341_sign_out(2);
    CN128_data_in(7) <= VN391_data_out(2);
    CN128_sign_in(7) <= VN391_sign_out(2);
    CN128_data_in(8) <= VN441_data_out(2);
    CN128_sign_in(8) <= VN441_sign_out(2);
    CN128_data_in(9) <= VN457_data_out(2);
    CN128_sign_in(9) <= VN457_sign_out(2);
    CN128_data_in(10) <= VN534_data_out(2);
    CN128_sign_in(10) <= VN534_sign_out(2);
    CN128_data_in(11) <= VN579_data_out(2);
    CN128_sign_in(11) <= VN579_sign_out(2);
    CN128_data_in(12) <= VN640_data_out(2);
    CN128_sign_in(12) <= VN640_sign_out(2);
    CN128_data_in(13) <= VN710_data_out(2);
    CN128_sign_in(13) <= VN710_sign_out(2);
    CN128_data_in(14) <= VN762_data_out(2);
    CN128_sign_in(14) <= VN762_sign_out(2);
    CN128_data_in(15) <= VN795_data_out(2);
    CN128_sign_in(15) <= VN795_sign_out(2);
    CN128_data_in(16) <= VN858_data_out(2);
    CN128_sign_in(16) <= VN858_sign_out(2);
    CN128_data_in(17) <= VN893_data_out(2);
    CN128_sign_in(17) <= VN893_sign_out(2);
    CN128_data_in(18) <= VN1002_data_out(2);
    CN128_sign_in(18) <= VN1002_sign_out(2);
    CN128_data_in(19) <= VN1037_data_out(2);
    CN128_sign_in(19) <= VN1037_sign_out(2);
    CN128_data_in(20) <= VN1073_data_out(2);
    CN128_sign_in(20) <= VN1073_sign_out(2);
    CN128_data_in(21) <= VN1157_data_out(2);
    CN128_sign_in(21) <= VN1157_sign_out(2);
    CN128_data_in(22) <= VN1170_data_out(2);
    CN128_sign_in(22) <= VN1170_sign_out(2);
    CN128_data_in(23) <= VN1244_data_out(2);
    CN128_sign_in(23) <= VN1244_sign_out(2);
    CN128_data_in(24) <= VN1286_data_out(2);
    CN128_sign_in(24) <= VN1286_sign_out(2);
    CN128_data_in(25) <= VN1345_data_out(2);
    CN128_sign_in(25) <= VN1345_sign_out(2);
    CN128_data_in(26) <= VN1493_data_out(2);
    CN128_sign_in(26) <= VN1493_sign_out(2);
    CN128_data_in(27) <= VN1573_data_out(2);
    CN128_sign_in(27) <= VN1573_sign_out(2);
    CN128_data_in(28) <= VN1581_data_out(2);
    CN128_sign_in(28) <= VN1581_sign_out(2);
    CN128_data_in(29) <= VN1707_data_out(2);
    CN128_sign_in(29) <= VN1707_sign_out(2);
    CN128_data_in(30) <= VN1781_data_out(2);
    CN128_sign_in(30) <= VN1781_sign_out(2);
    CN128_data_in(31) <= VN1831_data_out(2);
    CN128_sign_in(31) <= VN1831_sign_out(2);
    CN129_data_in(0) <= VN51_data_out(2);
    CN129_sign_in(0) <= VN51_sign_out(2);
    CN129_data_in(1) <= VN56_data_out(2);
    CN129_sign_in(1) <= VN56_sign_out(2);
    CN129_data_in(2) <= VN116_data_out(2);
    CN129_sign_in(2) <= VN116_sign_out(2);
    CN129_data_in(3) <= VN172_data_out(2);
    CN129_sign_in(3) <= VN172_sign_out(2);
    CN129_data_in(4) <= VN276_data_out(2);
    CN129_sign_in(4) <= VN276_sign_out(2);
    CN129_data_in(5) <= VN305_data_out(2);
    CN129_sign_in(5) <= VN305_sign_out(2);
    CN129_data_in(6) <= VN372_data_out(2);
    CN129_sign_in(6) <= VN372_sign_out(2);
    CN129_data_in(7) <= VN402_data_out(2);
    CN129_sign_in(7) <= VN402_sign_out(2);
    CN129_data_in(8) <= VN493_data_out(2);
    CN129_sign_in(8) <= VN493_sign_out(2);
    CN129_data_in(9) <= VN547_data_out(2);
    CN129_sign_in(9) <= VN547_sign_out(2);
    CN129_data_in(10) <= VN596_data_out(2);
    CN129_sign_in(10) <= VN596_sign_out(2);
    CN129_data_in(11) <= VN643_data_out(2);
    CN129_sign_in(11) <= VN643_sign_out(2);
    CN129_data_in(12) <= VN696_data_out(2);
    CN129_sign_in(12) <= VN696_sign_out(2);
    CN129_data_in(13) <= VN824_data_out(2);
    CN129_sign_in(13) <= VN824_sign_out(2);
    CN129_data_in(14) <= VN857_data_out(2);
    CN129_sign_in(14) <= VN857_sign_out(2);
    CN129_data_in(15) <= VN939_data_out(2);
    CN129_sign_in(15) <= VN939_sign_out(2);
    CN129_data_in(16) <= VN954_data_out(2);
    CN129_sign_in(16) <= VN954_sign_out(2);
    CN129_data_in(17) <= VN1053_data_out(2);
    CN129_sign_in(17) <= VN1053_sign_out(2);
    CN129_data_in(18) <= VN1107_data_out(2);
    CN129_sign_in(18) <= VN1107_sign_out(2);
    CN129_data_in(19) <= VN1119_data_out(2);
    CN129_sign_in(19) <= VN1119_sign_out(2);
    CN129_data_in(20) <= VN1209_data_out(2);
    CN129_sign_in(20) <= VN1209_sign_out(2);
    CN129_data_in(21) <= VN1220_data_out(2);
    CN129_sign_in(21) <= VN1220_sign_out(2);
    CN129_data_in(22) <= VN1291_data_out(2);
    CN129_sign_in(22) <= VN1291_sign_out(2);
    CN129_data_in(23) <= VN1371_data_out(2);
    CN129_sign_in(23) <= VN1371_sign_out(2);
    CN129_data_in(24) <= VN1413_data_out(2);
    CN129_sign_in(24) <= VN1413_sign_out(2);
    CN129_data_in(25) <= VN1429_data_out(2);
    CN129_sign_in(25) <= VN1429_sign_out(2);
    CN129_data_in(26) <= VN1499_data_out(2);
    CN129_sign_in(26) <= VN1499_sign_out(2);
    CN129_data_in(27) <= VN1586_data_out(2);
    CN129_sign_in(27) <= VN1586_sign_out(2);
    CN129_data_in(28) <= VN1617_data_out(2);
    CN129_sign_in(28) <= VN1617_sign_out(2);
    CN129_data_in(29) <= VN1655_data_out(2);
    CN129_sign_in(29) <= VN1655_sign_out(2);
    CN129_data_in(30) <= VN1705_data_out(2);
    CN129_sign_in(30) <= VN1705_sign_out(2);
    CN129_data_in(31) <= VN1756_data_out(2);
    CN129_sign_in(31) <= VN1756_sign_out(2);
    CN130_data_in(0) <= VN50_data_out(2);
    CN130_sign_in(0) <= VN50_sign_out(2);
    CN130_data_in(1) <= VN73_data_out(2);
    CN130_sign_in(1) <= VN73_sign_out(2);
    CN130_data_in(2) <= VN140_data_out(2);
    CN130_sign_in(2) <= VN140_sign_out(2);
    CN130_data_in(3) <= VN188_data_out(2);
    CN130_sign_in(3) <= VN188_sign_out(2);
    CN130_data_in(4) <= VN245_data_out(2);
    CN130_sign_in(4) <= VN245_sign_out(2);
    CN130_data_in(5) <= VN285_data_out(2);
    CN130_sign_in(5) <= VN285_sign_out(2);
    CN130_data_in(6) <= VN385_data_out(2);
    CN130_sign_in(6) <= VN385_sign_out(2);
    CN130_data_in(7) <= VN398_data_out(2);
    CN130_sign_in(7) <= VN398_sign_out(2);
    CN130_data_in(8) <= VN477_data_out(2);
    CN130_sign_in(8) <= VN477_sign_out(2);
    CN130_data_in(9) <= VN520_data_out(2);
    CN130_sign_in(9) <= VN520_sign_out(2);
    CN130_data_in(10) <= VN586_data_out(2);
    CN130_sign_in(10) <= VN586_sign_out(2);
    CN130_data_in(11) <= VN654_data_out(2);
    CN130_sign_in(11) <= VN654_sign_out(2);
    CN130_data_in(12) <= VN706_data_out(2);
    CN130_sign_in(12) <= VN706_sign_out(2);
    CN130_data_in(13) <= VN756_data_out(2);
    CN130_sign_in(13) <= VN756_sign_out(2);
    CN130_data_in(14) <= VN786_data_out(2);
    CN130_sign_in(14) <= VN786_sign_out(2);
    CN130_data_in(15) <= VN835_data_out(2);
    CN130_sign_in(15) <= VN835_sign_out(2);
    CN130_data_in(16) <= VN981_data_out(2);
    CN130_sign_in(16) <= VN981_sign_out(2);
    CN130_data_in(17) <= VN1014_data_out(2);
    CN130_sign_in(17) <= VN1014_sign_out(2);
    CN130_data_in(18) <= VN1099_data_out(2);
    CN130_sign_in(18) <= VN1099_sign_out(2);
    CN130_data_in(19) <= VN1189_data_out(2);
    CN130_sign_in(19) <= VN1189_sign_out(2);
    CN130_data_in(20) <= VN1230_data_out(2);
    CN130_sign_in(20) <= VN1230_sign_out(2);
    CN130_data_in(21) <= VN1292_data_out(2);
    CN130_sign_in(21) <= VN1292_sign_out(2);
    CN130_data_in(22) <= VN1359_data_out(2);
    CN130_sign_in(22) <= VN1359_sign_out(2);
    CN130_data_in(23) <= VN1401_data_out(2);
    CN130_sign_in(23) <= VN1401_sign_out(2);
    CN130_data_in(24) <= VN1439_data_out(2);
    CN130_sign_in(24) <= VN1439_sign_out(2);
    CN130_data_in(25) <= VN1465_data_out(2);
    CN130_sign_in(25) <= VN1465_sign_out(2);
    CN130_data_in(26) <= VN1513_data_out(2);
    CN130_sign_in(26) <= VN1513_sign_out(2);
    CN130_data_in(27) <= VN1556_data_out(2);
    CN130_sign_in(27) <= VN1556_sign_out(2);
    CN130_data_in(28) <= VN1620_data_out(2);
    CN130_sign_in(28) <= VN1620_sign_out(2);
    CN130_data_in(29) <= VN1718_data_out(2);
    CN130_sign_in(29) <= VN1718_sign_out(2);
    CN130_data_in(30) <= VN1773_data_out(2);
    CN130_sign_in(30) <= VN1773_sign_out(2);
    CN130_data_in(31) <= VN1832_data_out(2);
    CN130_sign_in(31) <= VN1832_sign_out(2);
    CN131_data_in(0) <= VN65_data_out(2);
    CN131_sign_in(0) <= VN65_sign_out(2);
    CN131_data_in(1) <= VN154_data_out(2);
    CN131_sign_in(1) <= VN154_sign_out(2);
    CN131_data_in(2) <= VN206_data_out(2);
    CN131_sign_in(2) <= VN206_sign_out(2);
    CN131_data_in(3) <= VN243_data_out(2);
    CN131_sign_in(3) <= VN243_sign_out(2);
    CN131_data_in(4) <= VN307_data_out(2);
    CN131_sign_in(4) <= VN307_sign_out(2);
    CN131_data_in(5) <= VN334_data_out(2);
    CN131_sign_in(5) <= VN334_sign_out(2);
    CN131_data_in(6) <= VN403_data_out(2);
    CN131_sign_in(6) <= VN403_sign_out(2);
    CN131_data_in(7) <= VN479_data_out(2);
    CN131_sign_in(7) <= VN479_sign_out(2);
    CN131_data_in(8) <= VN530_data_out(2);
    CN131_sign_in(8) <= VN530_sign_out(2);
    CN131_data_in(9) <= VN608_data_out(2);
    CN131_sign_in(9) <= VN608_sign_out(2);
    CN131_data_in(10) <= VN665_data_out(2);
    CN131_sign_in(10) <= VN665_sign_out(2);
    CN131_data_in(11) <= VN700_data_out(2);
    CN131_sign_in(11) <= VN700_sign_out(2);
    CN131_data_in(12) <= VN750_data_out(2);
    CN131_sign_in(12) <= VN750_sign_out(2);
    CN131_data_in(13) <= VN791_data_out(2);
    CN131_sign_in(13) <= VN791_sign_out(2);
    CN131_data_in(14) <= VN870_data_out(2);
    CN131_sign_in(14) <= VN870_sign_out(2);
    CN131_data_in(15) <= VN887_data_out(2);
    CN131_sign_in(15) <= VN887_sign_out(2);
    CN131_data_in(16) <= VN932_data_out(2);
    CN131_sign_in(16) <= VN932_sign_out(2);
    CN131_data_in(17) <= VN972_data_out(2);
    CN131_sign_in(17) <= VN972_sign_out(2);
    CN131_data_in(18) <= VN1044_data_out(2);
    CN131_sign_in(18) <= VN1044_sign_out(2);
    CN131_data_in(19) <= VN1064_data_out(2);
    CN131_sign_in(19) <= VN1064_sign_out(2);
    CN131_data_in(20) <= VN1143_data_out(2);
    CN131_sign_in(20) <= VN1143_sign_out(2);
    CN131_data_in(21) <= VN1173_data_out(2);
    CN131_sign_in(21) <= VN1173_sign_out(2);
    CN131_data_in(22) <= VN1264_data_out(2);
    CN131_sign_in(22) <= VN1264_sign_out(2);
    CN131_data_in(23) <= VN1321_data_out(2);
    CN131_sign_in(23) <= VN1321_sign_out(2);
    CN131_data_in(24) <= VN1377_data_out(2);
    CN131_sign_in(24) <= VN1377_sign_out(2);
    CN131_data_in(25) <= VN1551_data_out(2);
    CN131_sign_in(25) <= VN1551_sign_out(2);
    CN131_data_in(26) <= VN1572_data_out(2);
    CN131_sign_in(26) <= VN1572_sign_out(2);
    CN131_data_in(27) <= VN1605_data_out(2);
    CN131_sign_in(27) <= VN1605_sign_out(2);
    CN131_data_in(28) <= VN1608_data_out(2);
    CN131_sign_in(28) <= VN1608_sign_out(2);
    CN131_data_in(29) <= VN1674_data_out(2);
    CN131_sign_in(29) <= VN1674_sign_out(2);
    CN131_data_in(30) <= VN1792_data_out(2);
    CN131_sign_in(30) <= VN1792_sign_out(2);
    CN131_data_in(31) <= VN1833_data_out(2);
    CN131_sign_in(31) <= VN1833_sign_out(2);
    CN132_data_in(0) <= VN49_data_out(2);
    CN132_sign_in(0) <= VN49_sign_out(2);
    CN132_data_in(1) <= VN151_data_out(2);
    CN132_sign_in(1) <= VN151_sign_out(2);
    CN132_data_in(2) <= VN214_data_out(2);
    CN132_sign_in(2) <= VN214_sign_out(2);
    CN132_data_in(3) <= VN274_data_out(2);
    CN132_sign_in(3) <= VN274_sign_out(2);
    CN132_data_in(4) <= VN321_data_out(2);
    CN132_sign_in(4) <= VN321_sign_out(2);
    CN132_data_in(5) <= VN364_data_out(2);
    CN132_sign_in(5) <= VN364_sign_out(2);
    CN132_data_in(6) <= VN448_data_out(2);
    CN132_sign_in(6) <= VN448_sign_out(2);
    CN132_data_in(7) <= VN615_data_out(2);
    CN132_sign_in(7) <= VN615_sign_out(2);
    CN132_data_in(8) <= VN637_data_out(2);
    CN132_sign_in(8) <= VN637_sign_out(2);
    CN132_data_in(9) <= VN704_data_out(2);
    CN132_sign_in(9) <= VN704_sign_out(2);
    CN132_data_in(10) <= VN733_data_out(2);
    CN132_sign_in(10) <= VN733_sign_out(2);
    CN132_data_in(11) <= VN873_data_out(2);
    CN132_sign_in(11) <= VN873_sign_out(2);
    CN132_data_in(12) <= VN914_data_out(2);
    CN132_sign_in(12) <= VN914_sign_out(2);
    CN132_data_in(13) <= VN959_data_out(2);
    CN132_sign_in(13) <= VN959_sign_out(2);
    CN132_data_in(14) <= VN1041_data_out(2);
    CN132_sign_in(14) <= VN1041_sign_out(2);
    CN132_data_in(15) <= VN1185_data_out(2);
    CN132_sign_in(15) <= VN1185_sign_out(2);
    CN132_data_in(16) <= VN1247_data_out(2);
    CN132_sign_in(16) <= VN1247_sign_out(2);
    CN132_data_in(17) <= VN1352_data_out(2);
    CN132_sign_in(17) <= VN1352_sign_out(2);
    CN132_data_in(18) <= VN1404_data_out(2);
    CN132_sign_in(18) <= VN1404_sign_out(2);
    CN132_data_in(19) <= VN1482_data_out(2);
    CN132_sign_in(19) <= VN1482_sign_out(2);
    CN132_data_in(20) <= VN1500_data_out(2);
    CN132_sign_in(20) <= VN1500_sign_out(2);
    CN132_data_in(21) <= VN1560_data_out(2);
    CN132_sign_in(21) <= VN1560_sign_out(2);
    CN132_data_in(22) <= VN1635_data_out(2);
    CN132_sign_in(22) <= VN1635_sign_out(2);
    CN132_data_in(23) <= VN1778_data_out(2);
    CN132_sign_in(23) <= VN1778_sign_out(2);
    CN132_data_in(24) <= VN1809_data_out(2);
    CN132_sign_in(24) <= VN1809_sign_out(2);
    CN132_data_in(25) <= VN1940_data_out(2);
    CN132_sign_in(25) <= VN1940_sign_out(2);
    CN132_data_in(26) <= VN1947_data_out(2);
    CN132_sign_in(26) <= VN1947_sign_out(2);
    CN132_data_in(27) <= VN1982_data_out(2);
    CN132_sign_in(27) <= VN1982_sign_out(2);
    CN132_data_in(28) <= VN2017_data_out(2);
    CN132_sign_in(28) <= VN2017_sign_out(2);
    CN132_data_in(29) <= VN2042_data_out(2);
    CN132_sign_in(29) <= VN2042_sign_out(2);
    CN132_data_in(30) <= VN2044_data_out(2);
    CN132_sign_in(30) <= VN2044_sign_out(2);
    CN132_data_in(31) <= VN2047_data_out(2);
    CN132_sign_in(31) <= VN2047_sign_out(2);
    CN133_data_in(0) <= VN48_data_out(2);
    CN133_sign_in(0) <= VN48_sign_out(2);
    CN133_data_in(1) <= VN209_data_out(2);
    CN133_sign_in(1) <= VN209_sign_out(2);
    CN133_data_in(2) <= VN255_data_out(2);
    CN133_sign_in(2) <= VN255_sign_out(2);
    CN133_data_in(3) <= VN317_data_out(2);
    CN133_sign_in(3) <= VN317_sign_out(2);
    CN133_data_in(4) <= VN380_data_out(2);
    CN133_sign_in(4) <= VN380_sign_out(2);
    CN133_data_in(5) <= VN416_data_out(2);
    CN133_sign_in(5) <= VN416_sign_out(2);
    CN133_data_in(6) <= VN527_data_out(2);
    CN133_sign_in(6) <= VN527_sign_out(2);
    CN133_data_in(7) <= VN600_data_out(2);
    CN133_sign_in(7) <= VN600_sign_out(2);
    CN133_data_in(8) <= VN626_data_out(2);
    CN133_sign_in(8) <= VN626_sign_out(2);
    CN133_data_in(9) <= VN693_data_out(2);
    CN133_sign_in(9) <= VN693_sign_out(2);
    CN133_data_in(10) <= VN740_data_out(2);
    CN133_sign_in(10) <= VN740_sign_out(2);
    CN133_data_in(11) <= VN790_data_out(2);
    CN133_sign_in(11) <= VN790_sign_out(2);
    CN133_data_in(12) <= VN860_data_out(2);
    CN133_sign_in(12) <= VN860_sign_out(2);
    CN133_data_in(13) <= VN896_data_out(2);
    CN133_sign_in(13) <= VN896_sign_out(2);
    CN133_data_in(14) <= VN978_data_out(2);
    CN133_sign_in(14) <= VN978_sign_out(2);
    CN133_data_in(15) <= VN1058_data_out(2);
    CN133_sign_in(15) <= VN1058_sign_out(2);
    CN133_data_in(16) <= VN1147_data_out(2);
    CN133_sign_in(16) <= VN1147_sign_out(2);
    CN133_data_in(17) <= VN1194_data_out(2);
    CN133_sign_in(17) <= VN1194_sign_out(2);
    CN133_data_in(18) <= VN1259_data_out(2);
    CN133_sign_in(18) <= VN1259_sign_out(2);
    CN133_data_in(19) <= VN1349_data_out(2);
    CN133_sign_in(19) <= VN1349_sign_out(2);
    CN133_data_in(20) <= VN1423_data_out(2);
    CN133_sign_in(20) <= VN1423_sign_out(2);
    CN133_data_in(21) <= VN1441_data_out(2);
    CN133_sign_in(21) <= VN1441_sign_out(2);
    CN133_data_in(22) <= VN1509_data_out(2);
    CN133_sign_in(22) <= VN1509_sign_out(2);
    CN133_data_in(23) <= VN1528_data_out(2);
    CN133_sign_in(23) <= VN1528_sign_out(2);
    CN133_data_in(24) <= VN1555_data_out(2);
    CN133_sign_in(24) <= VN1555_sign_out(2);
    CN133_data_in(25) <= VN1577_data_out(2);
    CN133_sign_in(25) <= VN1577_sign_out(2);
    CN133_data_in(26) <= VN1675_data_out(2);
    CN133_sign_in(26) <= VN1675_sign_out(2);
    CN133_data_in(27) <= VN1878_data_out(2);
    CN133_sign_in(27) <= VN1878_sign_out(2);
    CN133_data_in(28) <= VN1929_data_out(2);
    CN133_sign_in(28) <= VN1929_sign_out(2);
    CN133_data_in(29) <= VN1938_data_out(2);
    CN133_sign_in(29) <= VN1938_sign_out(2);
    CN133_data_in(30) <= VN1945_data_out(2);
    CN133_sign_in(30) <= VN1945_sign_out(2);
    CN133_data_in(31) <= VN1952_data_out(2);
    CN133_sign_in(31) <= VN1952_sign_out(2);
    CN134_data_in(0) <= VN47_data_out(2);
    CN134_sign_in(0) <= VN47_sign_out(2);
    CN134_data_in(1) <= VN100_data_out(2);
    CN134_sign_in(1) <= VN100_sign_out(2);
    CN134_data_in(2) <= VN134_data_out(2);
    CN134_sign_in(2) <= VN134_sign_out(2);
    CN134_data_in(3) <= VN258_data_out(2);
    CN134_sign_in(3) <= VN258_sign_out(2);
    CN134_data_in(4) <= VN423_data_out(2);
    CN134_sign_in(4) <= VN423_sign_out(2);
    CN134_data_in(5) <= VN497_data_out(2);
    CN134_sign_in(5) <= VN497_sign_out(2);
    CN134_data_in(6) <= VN518_data_out(2);
    CN134_sign_in(6) <= VN518_sign_out(2);
    CN134_data_in(7) <= VN763_data_out(2);
    CN134_sign_in(7) <= VN763_sign_out(2);
    CN134_data_in(8) <= VN950_data_out(2);
    CN134_sign_in(8) <= VN950_sign_out(2);
    CN134_data_in(9) <= VN1050_data_out(2);
    CN134_sign_in(9) <= VN1050_sign_out(2);
    CN134_data_in(10) <= VN1068_data_out(2);
    CN134_sign_in(10) <= VN1068_sign_out(2);
    CN134_data_in(11) <= VN1151_data_out(2);
    CN134_sign_in(11) <= VN1151_sign_out(2);
    CN134_data_in(12) <= VN1271_data_out(2);
    CN134_sign_in(12) <= VN1271_sign_out(2);
    CN134_data_in(13) <= VN1281_data_out(2);
    CN134_sign_in(13) <= VN1281_sign_out(2);
    CN134_data_in(14) <= VN1284_data_out(2);
    CN134_sign_in(14) <= VN1284_sign_out(2);
    CN134_data_in(15) <= VN1607_data_out(2);
    CN134_sign_in(15) <= VN1607_sign_out(2);
    CN134_data_in(16) <= VN1628_data_out(2);
    CN134_sign_in(16) <= VN1628_sign_out(2);
    CN134_data_in(17) <= VN1668_data_out(2);
    CN134_sign_in(17) <= VN1668_sign_out(2);
    CN134_data_in(18) <= VN1694_data_out(2);
    CN134_sign_in(18) <= VN1694_sign_out(2);
    CN134_data_in(19) <= VN1750_data_out(2);
    CN134_sign_in(19) <= VN1750_sign_out(2);
    CN134_data_in(20) <= VN1787_data_out(2);
    CN134_sign_in(20) <= VN1787_sign_out(2);
    CN134_data_in(21) <= VN1850_data_out(2);
    CN134_sign_in(21) <= VN1850_sign_out(2);
    CN134_data_in(22) <= VN1856_data_out(2);
    CN134_sign_in(22) <= VN1856_sign_out(2);
    CN134_data_in(23) <= VN1869_data_out(2);
    CN134_sign_in(23) <= VN1869_sign_out(2);
    CN134_data_in(24) <= VN1880_data_out(2);
    CN134_sign_in(24) <= VN1880_sign_out(2);
    CN134_data_in(25) <= VN1941_data_out(2);
    CN134_sign_in(25) <= VN1941_sign_out(2);
    CN134_data_in(26) <= VN1964_data_out(2);
    CN134_sign_in(26) <= VN1964_sign_out(2);
    CN134_data_in(27) <= VN1965_data_out(2);
    CN134_sign_in(27) <= VN1965_sign_out(2);
    CN134_data_in(28) <= VN2001_data_out(2);
    CN134_sign_in(28) <= VN2001_sign_out(2);
    CN134_data_in(29) <= VN2008_data_out(2);
    CN134_sign_in(29) <= VN2008_sign_out(2);
    CN134_data_in(30) <= VN2014_data_out(2);
    CN134_sign_in(30) <= VN2014_sign_out(2);
    CN134_data_in(31) <= VN2023_data_out(2);
    CN134_sign_in(31) <= VN2023_sign_out(2);
    CN135_data_in(0) <= VN46_data_out(2);
    CN135_sign_in(0) <= VN46_sign_out(2);
    CN135_data_in(1) <= VN103_data_out(2);
    CN135_sign_in(1) <= VN103_sign_out(2);
    CN135_data_in(2) <= VN135_data_out(2);
    CN135_sign_in(2) <= VN135_sign_out(2);
    CN135_data_in(3) <= VN205_data_out(2);
    CN135_sign_in(3) <= VN205_sign_out(2);
    CN135_data_in(4) <= VN388_data_out(2);
    CN135_sign_in(4) <= VN388_sign_out(2);
    CN135_data_in(5) <= VN449_data_out(2);
    CN135_sign_in(5) <= VN449_sign_out(2);
    CN135_data_in(6) <= VN555_data_out(2);
    CN135_sign_in(6) <= VN555_sign_out(2);
    CN135_data_in(7) <= VN571_data_out(2);
    CN135_sign_in(7) <= VN571_sign_out(2);
    CN135_data_in(8) <= VN712_data_out(2);
    CN135_sign_in(8) <= VN712_sign_out(2);
    CN135_data_in(9) <= VN761_data_out(2);
    CN135_sign_in(9) <= VN761_sign_out(2);
    CN135_data_in(10) <= VN821_data_out(2);
    CN135_sign_in(10) <= VN821_sign_out(2);
    CN135_data_in(11) <= VN920_data_out(2);
    CN135_sign_in(11) <= VN920_sign_out(2);
    CN135_data_in(12) <= VN947_data_out(2);
    CN135_sign_in(12) <= VN947_sign_out(2);
    CN135_data_in(13) <= VN1062_data_out(2);
    CN135_sign_in(13) <= VN1062_sign_out(2);
    CN135_data_in(14) <= VN1140_data_out(2);
    CN135_sign_in(14) <= VN1140_sign_out(2);
    CN135_data_in(15) <= VN1211_data_out(2);
    CN135_sign_in(15) <= VN1211_sign_out(2);
    CN135_data_in(16) <= VN1357_data_out(2);
    CN135_sign_in(16) <= VN1357_sign_out(2);
    CN135_data_in(17) <= VN1387_data_out(2);
    CN135_sign_in(17) <= VN1387_sign_out(2);
    CN135_data_in(18) <= VN1447_data_out(2);
    CN135_sign_in(18) <= VN1447_sign_out(2);
    CN135_data_in(19) <= VN1487_data_out(2);
    CN135_sign_in(19) <= VN1487_sign_out(2);
    CN135_data_in(20) <= VN1532_data_out(2);
    CN135_sign_in(20) <= VN1532_sign_out(2);
    CN135_data_in(21) <= VN1537_data_out(2);
    CN135_sign_in(21) <= VN1537_sign_out(2);
    CN135_data_in(22) <= VN1686_data_out(2);
    CN135_sign_in(22) <= VN1686_sign_out(2);
    CN135_data_in(23) <= VN1816_data_out(2);
    CN135_sign_in(23) <= VN1816_sign_out(2);
    CN135_data_in(24) <= VN1817_data_out(2);
    CN135_sign_in(24) <= VN1817_sign_out(2);
    CN135_data_in(25) <= VN1824_data_out(2);
    CN135_sign_in(25) <= VN1824_sign_out(2);
    CN135_data_in(26) <= VN1846_data_out(2);
    CN135_sign_in(26) <= VN1846_sign_out(2);
    CN135_data_in(27) <= VN1851_data_out(2);
    CN135_sign_in(27) <= VN1851_sign_out(2);
    CN135_data_in(28) <= VN1886_data_out(2);
    CN135_sign_in(28) <= VN1886_sign_out(2);
    CN135_data_in(29) <= VN1994_data_out(2);
    CN135_sign_in(29) <= VN1994_sign_out(2);
    CN135_data_in(30) <= VN2005_data_out(2);
    CN135_sign_in(30) <= VN2005_sign_out(2);
    CN135_data_in(31) <= VN2010_data_out(2);
    CN135_sign_in(31) <= VN2010_sign_out(2);
    CN136_data_in(0) <= VN45_data_out(2);
    CN136_sign_in(0) <= VN45_sign_out(2);
    CN136_data_in(1) <= VN94_data_out(2);
    CN136_sign_in(1) <= VN94_sign_out(2);
    CN136_data_in(2) <= VN111_data_out(2);
    CN136_sign_in(2) <= VN111_sign_out(2);
    CN136_data_in(3) <= VN175_data_out(2);
    CN136_sign_in(3) <= VN175_sign_out(2);
    CN136_data_in(4) <= VN275_data_out(2);
    CN136_sign_in(4) <= VN275_sign_out(2);
    CN136_data_in(5) <= VN301_data_out(2);
    CN136_sign_in(5) <= VN301_sign_out(2);
    CN136_data_in(6) <= VN352_data_out(2);
    CN136_sign_in(6) <= VN352_sign_out(2);
    CN136_data_in(7) <= VN408_data_out(2);
    CN136_sign_in(7) <= VN408_sign_out(2);
    CN136_data_in(8) <= VN478_data_out(2);
    CN136_sign_in(8) <= VN478_sign_out(2);
    CN136_data_in(9) <= VN537_data_out(2);
    CN136_sign_in(9) <= VN537_sign_out(2);
    CN136_data_in(10) <= VN607_data_out(2);
    CN136_sign_in(10) <= VN607_sign_out(2);
    CN136_data_in(11) <= VN649_data_out(2);
    CN136_sign_in(11) <= VN649_sign_out(2);
    CN136_data_in(12) <= VN670_data_out(2);
    CN136_sign_in(12) <= VN670_sign_out(2);
    CN136_data_in(13) <= VN738_data_out(2);
    CN136_sign_in(13) <= VN738_sign_out(2);
    CN136_data_in(14) <= VN827_data_out(2);
    CN136_sign_in(14) <= VN827_sign_out(2);
    CN136_data_in(15) <= VN882_data_out(2);
    CN136_sign_in(15) <= VN882_sign_out(2);
    CN136_data_in(16) <= VN890_data_out(2);
    CN136_sign_in(16) <= VN890_sign_out(2);
    CN136_data_in(17) <= VN1097_data_out(2);
    CN136_sign_in(17) <= VN1097_sign_out(2);
    CN136_data_in(18) <= VN1120_data_out(2);
    CN136_sign_in(18) <= VN1120_sign_out(2);
    CN136_data_in(19) <= VN1197_data_out(2);
    CN136_sign_in(19) <= VN1197_sign_out(2);
    CN136_data_in(20) <= VN1232_data_out(2);
    CN136_sign_in(20) <= VN1232_sign_out(2);
    CN136_data_in(21) <= VN1283_data_out(2);
    CN136_sign_in(21) <= VN1283_sign_out(2);
    CN136_data_in(22) <= VN1451_data_out(2);
    CN136_sign_in(22) <= VN1451_sign_out(2);
    CN136_data_in(23) <= VN1480_data_out(2);
    CN136_sign_in(23) <= VN1480_sign_out(2);
    CN136_data_in(24) <= VN1540_data_out(2);
    CN136_sign_in(24) <= VN1540_sign_out(2);
    CN136_data_in(25) <= VN1636_data_out(2);
    CN136_sign_in(25) <= VN1636_sign_out(2);
    CN136_data_in(26) <= VN1777_data_out(2);
    CN136_sign_in(26) <= VN1777_sign_out(2);
    CN136_data_in(27) <= VN1845_data_out(2);
    CN136_sign_in(27) <= VN1845_sign_out(2);
    CN136_data_in(28) <= VN1894_data_out(2);
    CN136_sign_in(28) <= VN1894_sign_out(2);
    CN136_data_in(29) <= VN1939_data_out(2);
    CN136_sign_in(29) <= VN1939_sign_out(2);
    CN136_data_in(30) <= VN1949_data_out(2);
    CN136_sign_in(30) <= VN1949_sign_out(2);
    CN136_data_in(31) <= VN1953_data_out(2);
    CN136_sign_in(31) <= VN1953_sign_out(2);
    CN137_data_in(0) <= VN44_data_out(2);
    CN137_sign_in(0) <= VN44_sign_out(2);
    CN137_data_in(1) <= VN74_data_out(2);
    CN137_sign_in(1) <= VN74_sign_out(2);
    CN137_data_in(2) <= VN161_data_out(2);
    CN137_sign_in(2) <= VN161_sign_out(2);
    CN137_data_in(3) <= VN182_data_out(2);
    CN137_sign_in(3) <= VN182_sign_out(2);
    CN137_data_in(4) <= VN242_data_out(2);
    CN137_sign_in(4) <= VN242_sign_out(2);
    CN137_data_in(5) <= VN282_data_out(2);
    CN137_sign_in(5) <= VN282_sign_out(2);
    CN137_data_in(6) <= VN366_data_out(2);
    CN137_sign_in(6) <= VN366_sign_out(2);
    CN137_data_in(7) <= VN434_data_out(2);
    CN137_sign_in(7) <= VN434_sign_out(2);
    CN137_data_in(8) <= VN492_data_out(2);
    CN137_sign_in(8) <= VN492_sign_out(2);
    CN137_data_in(9) <= VN551_data_out(2);
    CN137_sign_in(9) <= VN551_sign_out(2);
    CN137_data_in(10) <= VN564_data_out(2);
    CN137_sign_in(10) <= VN564_sign_out(2);
    CN137_data_in(11) <= VN656_data_out(2);
    CN137_sign_in(11) <= VN656_sign_out(2);
    CN137_data_in(12) <= VN679_data_out(2);
    CN137_sign_in(12) <= VN679_sign_out(2);
    CN137_data_in(13) <= VN774_data_out(2);
    CN137_sign_in(13) <= VN774_sign_out(2);
    CN137_data_in(14) <= VN796_data_out(2);
    CN137_sign_in(14) <= VN796_sign_out(2);
    CN137_data_in(15) <= VN934_data_out(2);
    CN137_sign_in(15) <= VN934_sign_out(2);
    CN137_data_in(16) <= VN956_data_out(2);
    CN137_sign_in(16) <= VN956_sign_out(2);
    CN137_data_in(17) <= VN1028_data_out(2);
    CN137_sign_in(17) <= VN1028_sign_out(2);
    CN137_data_in(18) <= VN1103_data_out(2);
    CN137_sign_in(18) <= VN1103_sign_out(2);
    CN137_data_in(19) <= VN1160_data_out(2);
    CN137_sign_in(19) <= VN1160_sign_out(2);
    CN137_data_in(20) <= VN1213_data_out(2);
    CN137_sign_in(20) <= VN1213_sign_out(2);
    CN137_data_in(21) <= VN1274_data_out(2);
    CN137_sign_in(21) <= VN1274_sign_out(2);
    CN137_data_in(22) <= VN1341_data_out(2);
    CN137_sign_in(22) <= VN1341_sign_out(2);
    CN137_data_in(23) <= VN1422_data_out(2);
    CN137_sign_in(23) <= VN1422_sign_out(2);
    CN137_data_in(24) <= VN1427_data_out(2);
    CN137_sign_in(24) <= VN1427_sign_out(2);
    CN137_data_in(25) <= VN1526_data_out(2);
    CN137_sign_in(25) <= VN1526_sign_out(2);
    CN137_data_in(26) <= VN1678_data_out(2);
    CN137_sign_in(26) <= VN1678_sign_out(2);
    CN137_data_in(27) <= VN1693_data_out(2);
    CN137_sign_in(27) <= VN1693_sign_out(2);
    CN137_data_in(28) <= VN1724_data_out(2);
    CN137_sign_in(28) <= VN1724_sign_out(2);
    CN137_data_in(29) <= VN1731_data_out(2);
    CN137_sign_in(29) <= VN1731_sign_out(2);
    CN137_data_in(30) <= VN1893_data_out(2);
    CN137_sign_in(30) <= VN1893_sign_out(2);
    CN137_data_in(31) <= VN1909_data_out(2);
    CN137_sign_in(31) <= VN1909_sign_out(2);
    CN138_data_in(0) <= VN43_data_out(2);
    CN138_sign_in(0) <= VN43_sign_out(2);
    CN138_data_in(1) <= VN55_data_out(2);
    CN138_sign_in(1) <= VN55_sign_out(2);
    CN138_data_in(2) <= VN120_data_out(2);
    CN138_sign_in(2) <= VN120_sign_out(2);
    CN138_data_in(3) <= VN218_data_out(2);
    CN138_sign_in(3) <= VN218_sign_out(2);
    CN138_data_in(4) <= VN268_data_out(2);
    CN138_sign_in(4) <= VN268_sign_out(2);
    CN138_data_in(5) <= VN327_data_out(2);
    CN138_sign_in(5) <= VN327_sign_out(2);
    CN138_data_in(6) <= VN362_data_out(2);
    CN138_sign_in(6) <= VN362_sign_out(2);
    CN138_data_in(7) <= VN414_data_out(2);
    CN138_sign_in(7) <= VN414_sign_out(2);
    CN138_data_in(8) <= VN466_data_out(2);
    CN138_sign_in(8) <= VN466_sign_out(2);
    CN138_data_in(9) <= VN506_data_out(2);
    CN138_sign_in(9) <= VN506_sign_out(2);
    CN138_data_in(10) <= VN572_data_out(2);
    CN138_sign_in(10) <= VN572_sign_out(2);
    CN138_data_in(11) <= VN653_data_out(2);
    CN138_sign_in(11) <= VN653_sign_out(2);
    CN138_data_in(12) <= VN707_data_out(2);
    CN138_sign_in(12) <= VN707_sign_out(2);
    CN138_data_in(13) <= VN776_data_out(2);
    CN138_sign_in(13) <= VN776_sign_out(2);
    CN138_data_in(14) <= VN794_data_out(2);
    CN138_sign_in(14) <= VN794_sign_out(2);
    CN138_data_in(15) <= VN837_data_out(2);
    CN138_sign_in(15) <= VN837_sign_out(2);
    CN138_data_in(16) <= VN922_data_out(2);
    CN138_sign_in(16) <= VN922_sign_out(2);
    CN138_data_in(17) <= VN989_data_out(2);
    CN138_sign_in(17) <= VN989_sign_out(2);
    CN138_data_in(18) <= VN1031_data_out(2);
    CN138_sign_in(18) <= VN1031_sign_out(2);
    CN138_data_in(19) <= VN1074_data_out(2);
    CN138_sign_in(19) <= VN1074_sign_out(2);
    CN138_data_in(20) <= VN1115_data_out(2);
    CN138_sign_in(20) <= VN1115_sign_out(2);
    CN138_data_in(21) <= VN1177_data_out(2);
    CN138_sign_in(21) <= VN1177_sign_out(2);
    CN138_data_in(22) <= VN1310_data_out(2);
    CN138_sign_in(22) <= VN1310_sign_out(2);
    CN138_data_in(23) <= VN1431_data_out(2);
    CN138_sign_in(23) <= VN1431_sign_out(2);
    CN138_data_in(24) <= VN1450_data_out(2);
    CN138_sign_in(24) <= VN1450_sign_out(2);
    CN138_data_in(25) <= VN1461_data_out(2);
    CN138_sign_in(25) <= VN1461_sign_out(2);
    CN138_data_in(26) <= VN1618_data_out(2);
    CN138_sign_in(26) <= VN1618_sign_out(2);
    CN138_data_in(27) <= VN1680_data_out(2);
    CN138_sign_in(27) <= VN1680_sign_out(2);
    CN138_data_in(28) <= VN1712_data_out(2);
    CN138_sign_in(28) <= VN1712_sign_out(2);
    CN138_data_in(29) <= VN1744_data_out(2);
    CN138_sign_in(29) <= VN1744_sign_out(2);
    CN138_data_in(30) <= VN1794_data_out(2);
    CN138_sign_in(30) <= VN1794_sign_out(2);
    CN138_data_in(31) <= VN1834_data_out(2);
    CN138_sign_in(31) <= VN1834_sign_out(2);
    CN139_data_in(0) <= VN42_data_out(2);
    CN139_sign_in(0) <= VN42_sign_out(2);
    CN139_data_in(1) <= VN69_data_out(2);
    CN139_sign_in(1) <= VN69_sign_out(2);
    CN139_data_in(2) <= VN124_data_out(2);
    CN139_sign_in(2) <= VN124_sign_out(2);
    CN139_data_in(3) <= VN220_data_out(2);
    CN139_sign_in(3) <= VN220_sign_out(2);
    CN139_data_in(4) <= VN252_data_out(2);
    CN139_sign_in(4) <= VN252_sign_out(2);
    CN139_data_in(5) <= VN289_data_out(2);
    CN139_sign_in(5) <= VN289_sign_out(2);
    CN139_data_in(6) <= VN383_data_out(2);
    CN139_sign_in(6) <= VN383_sign_out(2);
    CN139_data_in(7) <= VN426_data_out(2);
    CN139_sign_in(7) <= VN426_sign_out(2);
    CN139_data_in(8) <= VN500_data_out(2);
    CN139_sign_in(8) <= VN500_sign_out(2);
    CN139_data_in(9) <= VN531_data_out(2);
    CN139_sign_in(9) <= VN531_sign_out(2);
    CN139_data_in(10) <= VN601_data_out(2);
    CN139_sign_in(10) <= VN601_sign_out(2);
    CN139_data_in(11) <= VN657_data_out(2);
    CN139_sign_in(11) <= VN657_sign_out(2);
    CN139_data_in(12) <= VN695_data_out(2);
    CN139_sign_in(12) <= VN695_sign_out(2);
    CN139_data_in(13) <= VN884_data_out(2);
    CN139_sign_in(13) <= VN884_sign_out(2);
    CN139_data_in(14) <= VN937_data_out(2);
    CN139_sign_in(14) <= VN937_sign_out(2);
    CN139_data_in(15) <= VN999_data_out(2);
    CN139_sign_in(15) <= VN999_sign_out(2);
    CN139_data_in(16) <= VN1022_data_out(2);
    CN139_sign_in(16) <= VN1022_sign_out(2);
    CN139_data_in(17) <= VN1072_data_out(2);
    CN139_sign_in(17) <= VN1072_sign_out(2);
    CN139_data_in(18) <= VN1126_data_out(2);
    CN139_sign_in(18) <= VN1126_sign_out(2);
    CN139_data_in(19) <= VN1186_data_out(2);
    CN139_sign_in(19) <= VN1186_sign_out(2);
    CN139_data_in(20) <= VN1253_data_out(2);
    CN139_sign_in(20) <= VN1253_sign_out(2);
    CN139_data_in(21) <= VN1317_data_out(2);
    CN139_sign_in(21) <= VN1317_sign_out(2);
    CN139_data_in(22) <= VN1338_data_out(2);
    CN139_sign_in(22) <= VN1338_sign_out(2);
    CN139_data_in(23) <= VN1386_data_out(2);
    CN139_sign_in(23) <= VN1386_sign_out(2);
    CN139_data_in(24) <= VN1396_data_out(2);
    CN139_sign_in(24) <= VN1396_sign_out(2);
    CN139_data_in(25) <= VN1445_data_out(2);
    CN139_sign_in(25) <= VN1445_sign_out(2);
    CN139_data_in(26) <= VN1582_data_out(2);
    CN139_sign_in(26) <= VN1582_sign_out(2);
    CN139_data_in(27) <= VN1633_data_out(2);
    CN139_sign_in(27) <= VN1633_sign_out(2);
    CN139_data_in(28) <= VN1746_data_out(2);
    CN139_sign_in(28) <= VN1746_sign_out(2);
    CN139_data_in(29) <= VN1779_data_out(2);
    CN139_sign_in(29) <= VN1779_sign_out(2);
    CN139_data_in(30) <= VN1815_data_out(2);
    CN139_sign_in(30) <= VN1815_sign_out(2);
    CN139_data_in(31) <= VN1881_data_out(2);
    CN139_sign_in(31) <= VN1881_sign_out(2);
    CN140_data_in(0) <= VN41_data_out(2);
    CN140_sign_in(0) <= VN41_sign_out(2);
    CN140_data_in(1) <= VN80_data_out(2);
    CN140_sign_in(1) <= VN80_sign_out(2);
    CN140_data_in(2) <= VN170_data_out(2);
    CN140_sign_in(2) <= VN170_sign_out(2);
    CN140_data_in(3) <= VN191_data_out(2);
    CN140_sign_in(3) <= VN191_sign_out(2);
    CN140_data_in(4) <= VN277_data_out(2);
    CN140_sign_in(4) <= VN277_sign_out(2);
    CN140_data_in(5) <= VN293_data_out(2);
    CN140_sign_in(5) <= VN293_sign_out(2);
    CN140_data_in(6) <= VN346_data_out(2);
    CN140_sign_in(6) <= VN346_sign_out(2);
    CN140_data_in(7) <= VN435_data_out(2);
    CN140_sign_in(7) <= VN435_sign_out(2);
    CN140_data_in(8) <= VN467_data_out(2);
    CN140_sign_in(8) <= VN467_sign_out(2);
    CN140_data_in(9) <= VN519_data_out(2);
    CN140_sign_in(9) <= VN519_sign_out(2);
    CN140_data_in(10) <= VN614_data_out(2);
    CN140_sign_in(10) <= VN614_sign_out(2);
    CN140_data_in(11) <= VN648_data_out(2);
    CN140_sign_in(11) <= VN648_sign_out(2);
    CN140_data_in(12) <= VN681_data_out(2);
    CN140_sign_in(12) <= VN681_sign_out(2);
    CN140_data_in(13) <= VN739_data_out(2);
    CN140_sign_in(13) <= VN739_sign_out(2);
    CN140_data_in(14) <= VN806_data_out(2);
    CN140_sign_in(14) <= VN806_sign_out(2);
    CN140_data_in(15) <= VN871_data_out(2);
    CN140_sign_in(15) <= VN871_sign_out(2);
    CN140_data_in(16) <= VN902_data_out(2);
    CN140_sign_in(16) <= VN902_sign_out(2);
    CN140_data_in(17) <= VN992_data_out(2);
    CN140_sign_in(17) <= VN992_sign_out(2);
    CN140_data_in(18) <= VN1101_data_out(2);
    CN140_sign_in(18) <= VN1101_sign_out(2);
    CN140_data_in(19) <= VN1154_data_out(2);
    CN140_sign_in(19) <= VN1154_sign_out(2);
    CN140_data_in(20) <= VN1182_data_out(2);
    CN140_sign_in(20) <= VN1182_sign_out(2);
    CN140_data_in(21) <= VN1261_data_out(2);
    CN140_sign_in(21) <= VN1261_sign_out(2);
    CN140_data_in(22) <= VN1278_data_out(2);
    CN140_sign_in(22) <= VN1278_sign_out(2);
    CN140_data_in(23) <= VN1287_data_out(2);
    CN140_sign_in(23) <= VN1287_sign_out(2);
    CN140_data_in(24) <= VN1467_data_out(2);
    CN140_sign_in(24) <= VN1467_sign_out(2);
    CN140_data_in(25) <= VN1504_data_out(2);
    CN140_sign_in(25) <= VN1504_sign_out(2);
    CN140_data_in(26) <= VN1533_data_out(2);
    CN140_sign_in(26) <= VN1533_sign_out(2);
    CN140_data_in(27) <= VN1544_data_out(2);
    CN140_sign_in(27) <= VN1544_sign_out(2);
    CN140_data_in(28) <= VN1580_data_out(2);
    CN140_sign_in(28) <= VN1580_sign_out(2);
    CN140_data_in(29) <= VN1611_data_out(2);
    CN140_sign_in(29) <= VN1611_sign_out(2);
    CN140_data_in(30) <= VN1708_data_out(2);
    CN140_sign_in(30) <= VN1708_sign_out(2);
    CN140_data_in(31) <= VN1757_data_out(2);
    CN140_sign_in(31) <= VN1757_sign_out(2);
    CN141_data_in(0) <= VN123_data_out(2);
    CN141_sign_in(0) <= VN123_sign_out(2);
    CN141_data_in(1) <= VN173_data_out(2);
    CN141_sign_in(1) <= VN173_sign_out(2);
    CN141_data_in(2) <= VN269_data_out(2);
    CN141_sign_in(2) <= VN269_sign_out(2);
    CN141_data_in(3) <= VN332_data_out(2);
    CN141_sign_in(3) <= VN332_sign_out(2);
    CN141_data_in(4) <= VN347_data_out(2);
    CN141_sign_in(4) <= VN347_sign_out(2);
    CN141_data_in(5) <= VN407_data_out(2);
    CN141_sign_in(5) <= VN407_sign_out(2);
    CN141_data_in(6) <= VN480_data_out(2);
    CN141_sign_in(6) <= VN480_sign_out(2);
    CN141_data_in(7) <= VN508_data_out(2);
    CN141_sign_in(7) <= VN508_sign_out(2);
    CN141_data_in(8) <= VN618_data_out(2);
    CN141_sign_in(8) <= VN618_sign_out(2);
    CN141_data_in(9) <= VN698_data_out(2);
    CN141_sign_in(9) <= VN698_sign_out(2);
    CN141_data_in(10) <= VN760_data_out(2);
    CN141_sign_in(10) <= VN760_sign_out(2);
    CN141_data_in(11) <= VN809_data_out(2);
    CN141_sign_in(11) <= VN809_sign_out(2);
    CN141_data_in(12) <= VN834_data_out(2);
    CN141_sign_in(12) <= VN834_sign_out(2);
    CN141_data_in(13) <= VN911_data_out(2);
    CN141_sign_in(13) <= VN911_sign_out(2);
    CN141_data_in(14) <= VN996_data_out(2);
    CN141_sign_in(14) <= VN996_sign_out(2);
    CN141_data_in(15) <= VN1040_data_out(2);
    CN141_sign_in(15) <= VN1040_sign_out(2);
    CN141_data_in(16) <= VN1085_data_out(2);
    CN141_sign_in(16) <= VN1085_sign_out(2);
    CN141_data_in(17) <= VN1142_data_out(2);
    CN141_sign_in(17) <= VN1142_sign_out(2);
    CN141_data_in(18) <= VN1187_data_out(2);
    CN141_sign_in(18) <= VN1187_sign_out(2);
    CN141_data_in(19) <= VN1332_data_out(2);
    CN141_sign_in(19) <= VN1332_sign_out(2);
    CN141_data_in(20) <= VN1364_data_out(2);
    CN141_sign_in(20) <= VN1364_sign_out(2);
    CN141_data_in(21) <= VN1459_data_out(2);
    CN141_sign_in(21) <= VN1459_sign_out(2);
    CN141_data_in(22) <= VN1474_data_out(2);
    CN141_sign_in(22) <= VN1474_sign_out(2);
    CN141_data_in(23) <= VN1546_data_out(2);
    CN141_sign_in(23) <= VN1546_sign_out(2);
    CN141_data_in(24) <= VN1741_data_out(2);
    CN141_sign_in(24) <= VN1741_sign_out(2);
    CN141_data_in(25) <= VN1788_data_out(2);
    CN141_sign_in(25) <= VN1788_sign_out(2);
    CN141_data_in(26) <= VN1810_data_out(2);
    CN141_sign_in(26) <= VN1810_sign_out(2);
    CN141_data_in(27) <= VN1814_data_out(2);
    CN141_sign_in(27) <= VN1814_sign_out(2);
    CN141_data_in(28) <= VN1848_data_out(2);
    CN141_sign_in(28) <= VN1848_sign_out(2);
    CN141_data_in(29) <= VN1872_data_out(2);
    CN141_sign_in(29) <= VN1872_sign_out(2);
    CN141_data_in(30) <= VN1879_data_out(2);
    CN141_sign_in(30) <= VN1879_sign_out(2);
    CN141_data_in(31) <= VN1910_data_out(2);
    CN141_sign_in(31) <= VN1910_sign_out(2);
    CN142_data_in(0) <= VN40_data_out(2);
    CN142_sign_in(0) <= VN40_sign_out(2);
    CN142_data_in(1) <= VN96_data_out(2);
    CN142_sign_in(1) <= VN96_sign_out(2);
    CN142_data_in(2) <= VN118_data_out(2);
    CN142_sign_in(2) <= VN118_sign_out(2);
    CN142_data_in(3) <= VN256_data_out(2);
    CN142_sign_in(3) <= VN256_sign_out(2);
    CN142_data_in(4) <= VN382_data_out(2);
    CN142_sign_in(4) <= VN382_sign_out(2);
    CN142_data_in(5) <= VN422_data_out(2);
    CN142_sign_in(5) <= VN422_sign_out(2);
    CN142_data_in(6) <= VN522_data_out(2);
    CN142_sign_in(6) <= VN522_sign_out(2);
    CN142_data_in(7) <= VN567_data_out(2);
    CN142_sign_in(7) <= VN567_sign_out(2);
    CN142_data_in(8) <= VN623_data_out(2);
    CN142_sign_in(8) <= VN623_sign_out(2);
    CN142_data_in(9) <= VN907_data_out(2);
    CN142_sign_in(9) <= VN907_sign_out(2);
    CN142_data_in(10) <= VN986_data_out(2);
    CN142_sign_in(10) <= VN986_sign_out(2);
    CN142_data_in(11) <= VN1054_data_out(2);
    CN142_sign_in(11) <= VN1054_sign_out(2);
    CN142_data_in(12) <= VN1129_data_out(2);
    CN142_sign_in(12) <= VN1129_sign_out(2);
    CN142_data_in(13) <= VN1262_data_out(2);
    CN142_sign_in(13) <= VN1262_sign_out(2);
    CN142_data_in(14) <= VN1315_data_out(2);
    CN142_sign_in(14) <= VN1315_sign_out(2);
    CN142_data_in(15) <= VN1348_data_out(2);
    CN142_sign_in(15) <= VN1348_sign_out(2);
    CN142_data_in(16) <= VN1408_data_out(2);
    CN142_sign_in(16) <= VN1408_sign_out(2);
    CN142_data_in(17) <= VN1623_data_out(2);
    CN142_sign_in(17) <= VN1623_sign_out(2);
    CN142_data_in(18) <= VN1658_data_out(2);
    CN142_sign_in(18) <= VN1658_sign_out(2);
    CN142_data_in(19) <= VN1747_data_out(2);
    CN142_sign_in(19) <= VN1747_sign_out(2);
    CN142_data_in(20) <= VN1797_data_out(2);
    CN142_sign_in(20) <= VN1797_sign_out(2);
    CN142_data_in(21) <= VN1818_data_out(2);
    CN142_sign_in(21) <= VN1818_sign_out(2);
    CN142_data_in(22) <= VN1827_data_out(2);
    CN142_sign_in(22) <= VN1827_sign_out(2);
    CN142_data_in(23) <= VN1873_data_out(2);
    CN142_sign_in(23) <= VN1873_sign_out(2);
    CN142_data_in(24) <= VN1899_data_out(2);
    CN142_sign_in(24) <= VN1899_sign_out(2);
    CN142_data_in(25) <= VN1902_data_out(2);
    CN142_sign_in(25) <= VN1902_sign_out(2);
    CN142_data_in(26) <= VN1918_data_out(2);
    CN142_sign_in(26) <= VN1918_sign_out(2);
    CN142_data_in(27) <= VN1955_data_out(2);
    CN142_sign_in(27) <= VN1955_sign_out(2);
    CN142_data_in(28) <= VN1973_data_out(2);
    CN142_sign_in(28) <= VN1973_sign_out(2);
    CN142_data_in(29) <= VN1989_data_out(2);
    CN142_sign_in(29) <= VN1989_sign_out(2);
    CN142_data_in(30) <= VN1998_data_out(2);
    CN142_sign_in(30) <= VN1998_sign_out(2);
    CN142_data_in(31) <= VN2003_data_out(2);
    CN142_sign_in(31) <= VN2003_sign_out(2);
    CN143_data_in(0) <= VN39_data_out(2);
    CN143_sign_in(0) <= VN39_sign_out(2);
    CN143_data_in(1) <= VN83_data_out(2);
    CN143_sign_in(1) <= VN83_sign_out(2);
    CN143_data_in(2) <= VN158_data_out(2);
    CN143_sign_in(2) <= VN158_sign_out(2);
    CN143_data_in(3) <= VN192_data_out(2);
    CN143_sign_in(3) <= VN192_sign_out(2);
    CN143_data_in(4) <= VN273_data_out(2);
    CN143_sign_in(4) <= VN273_sign_out(2);
    CN143_data_in(5) <= VN287_data_out(2);
    CN143_sign_in(5) <= VN287_sign_out(2);
    CN143_data_in(6) <= VN373_data_out(2);
    CN143_sign_in(6) <= VN373_sign_out(2);
    CN143_data_in(7) <= VN394_data_out(2);
    CN143_sign_in(7) <= VN394_sign_out(2);
    CN143_data_in(8) <= VN495_data_out(2);
    CN143_sign_in(8) <= VN495_sign_out(2);
    CN143_data_in(9) <= VN543_data_out(2);
    CN143_sign_in(9) <= VN543_sign_out(2);
    CN143_data_in(10) <= VN589_data_out(2);
    CN143_sign_in(10) <= VN589_sign_out(2);
    CN143_data_in(11) <= VN661_data_out(2);
    CN143_sign_in(11) <= VN661_sign_out(2);
    CN143_data_in(12) <= VN671_data_out(2);
    CN143_sign_in(12) <= VN671_sign_out(2);
    CN143_data_in(13) <= VN771_data_out(2);
    CN143_sign_in(13) <= VN771_sign_out(2);
    CN143_data_in(14) <= VN862_data_out(2);
    CN143_sign_in(14) <= VN862_sign_out(2);
    CN143_data_in(15) <= VN912_data_out(2);
    CN143_sign_in(15) <= VN912_sign_out(2);
    CN143_data_in(16) <= VN964_data_out(2);
    CN143_sign_in(16) <= VN964_sign_out(2);
    CN143_data_in(17) <= VN1008_data_out(2);
    CN143_sign_in(17) <= VN1008_sign_out(2);
    CN143_data_in(18) <= VN1075_data_out(2);
    CN143_sign_in(18) <= VN1075_sign_out(2);
    CN143_data_in(19) <= VN1145_data_out(2);
    CN143_sign_in(19) <= VN1145_sign_out(2);
    CN143_data_in(20) <= VN1199_data_out(2);
    CN143_sign_in(20) <= VN1199_sign_out(2);
    CN143_data_in(21) <= VN1252_data_out(2);
    CN143_sign_in(21) <= VN1252_sign_out(2);
    CN143_data_in(22) <= VN1299_data_out(2);
    CN143_sign_in(22) <= VN1299_sign_out(2);
    CN143_data_in(23) <= VN1360_data_out(2);
    CN143_sign_in(23) <= VN1360_sign_out(2);
    CN143_data_in(24) <= VN1391_data_out(2);
    CN143_sign_in(24) <= VN1391_sign_out(2);
    CN143_data_in(25) <= VN1436_data_out(2);
    CN143_sign_in(25) <= VN1436_sign_out(2);
    CN143_data_in(26) <= VN1455_data_out(2);
    CN143_sign_in(26) <= VN1455_sign_out(2);
    CN143_data_in(27) <= VN1592_data_out(2);
    CN143_sign_in(27) <= VN1592_sign_out(2);
    CN143_data_in(28) <= VN1615_data_out(2);
    CN143_sign_in(28) <= VN1615_sign_out(2);
    CN143_data_in(29) <= VN1679_data_out(2);
    CN143_sign_in(29) <= VN1679_sign_out(2);
    CN143_data_in(30) <= VN1688_data_out(2);
    CN143_sign_in(30) <= VN1688_sign_out(2);
    CN143_data_in(31) <= VN1758_data_out(2);
    CN143_sign_in(31) <= VN1758_sign_out(2);
    CN144_data_in(0) <= VN38_data_out(2);
    CN144_sign_in(0) <= VN38_sign_out(2);
    CN144_data_in(1) <= VN98_data_out(2);
    CN144_sign_in(1) <= VN98_sign_out(2);
    CN144_data_in(2) <= VN166_data_out(2);
    CN144_sign_in(2) <= VN166_sign_out(2);
    CN144_data_in(3) <= VN219_data_out(2);
    CN144_sign_in(3) <= VN219_sign_out(2);
    CN144_data_in(4) <= VN249_data_out(2);
    CN144_sign_in(4) <= VN249_sign_out(2);
    CN144_data_in(5) <= VN324_data_out(2);
    CN144_sign_in(5) <= VN324_sign_out(2);
    CN144_data_in(6) <= VN333_data_out(2);
    CN144_sign_in(6) <= VN333_sign_out(2);
    CN144_data_in(7) <= VN429_data_out(2);
    CN144_sign_in(7) <= VN429_sign_out(2);
    CN144_data_in(8) <= VN462_data_out(2);
    CN144_sign_in(8) <= VN462_sign_out(2);
    CN144_data_in(9) <= VN553_data_out(2);
    CN144_sign_in(9) <= VN553_sign_out(2);
    CN144_data_in(10) <= VN602_data_out(2);
    CN144_sign_in(10) <= VN602_sign_out(2);
    CN144_data_in(11) <= VN663_data_out(2);
    CN144_sign_in(11) <= VN663_sign_out(2);
    CN144_data_in(12) <= VN720_data_out(2);
    CN144_sign_in(12) <= VN720_sign_out(2);
    CN144_data_in(13) <= VN741_data_out(2);
    CN144_sign_in(13) <= VN741_sign_out(2);
    CN144_data_in(14) <= VN793_data_out(2);
    CN144_sign_in(14) <= VN793_sign_out(2);
    CN144_data_in(15) <= VN876_data_out(2);
    CN144_sign_in(15) <= VN876_sign_out(2);
    CN144_data_in(16) <= VN901_data_out(2);
    CN144_sign_in(16) <= VN901_sign_out(2);
    CN144_data_in(17) <= VN946_data_out(2);
    CN144_sign_in(17) <= VN946_sign_out(2);
    CN144_data_in(18) <= VN1034_data_out(2);
    CN144_sign_in(18) <= VN1034_sign_out(2);
    CN144_data_in(19) <= VN1102_data_out(2);
    CN144_sign_in(19) <= VN1102_sign_out(2);
    CN144_data_in(20) <= VN1206_data_out(2);
    CN144_sign_in(20) <= VN1206_sign_out(2);
    CN144_data_in(21) <= VN1301_data_out(2);
    CN144_sign_in(21) <= VN1301_sign_out(2);
    CN144_data_in(22) <= VN1330_data_out(2);
    CN144_sign_in(22) <= VN1330_sign_out(2);
    CN144_data_in(23) <= VN1370_data_out(2);
    CN144_sign_in(23) <= VN1370_sign_out(2);
    CN144_data_in(24) <= VN1400_data_out(2);
    CN144_sign_in(24) <= VN1400_sign_out(2);
    CN144_data_in(25) <= VN1511_data_out(2);
    CN144_sign_in(25) <= VN1511_sign_out(2);
    CN144_data_in(26) <= VN1520_data_out(2);
    CN144_sign_in(26) <= VN1520_sign_out(2);
    CN144_data_in(27) <= VN1566_data_out(2);
    CN144_sign_in(27) <= VN1566_sign_out(2);
    CN144_data_in(28) <= VN1583_data_out(2);
    CN144_sign_in(28) <= VN1583_sign_out(2);
    CN144_data_in(29) <= VN1643_data_out(2);
    CN144_sign_in(29) <= VN1643_sign_out(2);
    CN144_data_in(30) <= VN1785_data_out(2);
    CN144_sign_in(30) <= VN1785_sign_out(2);
    CN144_data_in(31) <= VN1835_data_out(2);
    CN144_sign_in(31) <= VN1835_sign_out(2);
    CN145_data_in(0) <= VN37_data_out(2);
    CN145_sign_in(0) <= VN37_sign_out(2);
    CN145_data_in(1) <= VN61_data_out(2);
    CN145_sign_in(1) <= VN61_sign_out(2);
    CN145_data_in(2) <= VN130_data_out(2);
    CN145_sign_in(2) <= VN130_sign_out(2);
    CN145_data_in(3) <= VN181_data_out(2);
    CN145_sign_in(3) <= VN181_sign_out(2);
    CN145_data_in(4) <= VN247_data_out(2);
    CN145_sign_in(4) <= VN247_sign_out(2);
    CN145_data_in(5) <= VN331_data_out(2);
    CN145_sign_in(5) <= VN331_sign_out(2);
    CN145_data_in(6) <= VN336_data_out(2);
    CN145_sign_in(6) <= VN336_sign_out(2);
    CN145_data_in(7) <= VN396_data_out(2);
    CN145_sign_in(7) <= VN396_sign_out(2);
    CN145_data_in(8) <= VN463_data_out(2);
    CN145_sign_in(8) <= VN463_sign_out(2);
    CN145_data_in(9) <= VN548_data_out(2);
    CN145_sign_in(9) <= VN548_sign_out(2);
    CN145_data_in(10) <= VN599_data_out(2);
    CN145_sign_in(10) <= VN599_sign_out(2);
    CN145_data_in(11) <= VN631_data_out(2);
    CN145_sign_in(11) <= VN631_sign_out(2);
    CN145_data_in(12) <= VN672_data_out(2);
    CN145_sign_in(12) <= VN672_sign_out(2);
    CN145_data_in(13) <= VN732_data_out(2);
    CN145_sign_in(13) <= VN732_sign_out(2);
    CN145_data_in(14) <= VN819_data_out(2);
    CN145_sign_in(14) <= VN819_sign_out(2);
    CN145_data_in(15) <= VN868_data_out(2);
    CN145_sign_in(15) <= VN868_sign_out(2);
    CN145_data_in(16) <= VN925_data_out(2);
    CN145_sign_in(16) <= VN925_sign_out(2);
    CN145_data_in(17) <= VN960_data_out(2);
    CN145_sign_in(17) <= VN960_sign_out(2);
    CN145_data_in(18) <= VN1024_data_out(2);
    CN145_sign_in(18) <= VN1024_sign_out(2);
    CN145_data_in(19) <= VN1071_data_out(2);
    CN145_sign_in(19) <= VN1071_sign_out(2);
    CN145_data_in(20) <= VN1117_data_out(2);
    CN145_sign_in(20) <= VN1117_sign_out(2);
    CN145_data_in(21) <= VN1165_data_out(2);
    CN145_sign_in(21) <= VN1165_sign_out(2);
    CN145_data_in(22) <= VN1191_data_out(2);
    CN145_sign_in(22) <= VN1191_sign_out(2);
    CN145_data_in(23) <= VN1227_data_out(2);
    CN145_sign_in(23) <= VN1227_sign_out(2);
    CN145_data_in(24) <= VN1288_data_out(2);
    CN145_sign_in(24) <= VN1288_sign_out(2);
    CN145_data_in(25) <= VN1342_data_out(2);
    CN145_sign_in(25) <= VN1342_sign_out(2);
    CN145_data_in(26) <= VN1409_data_out(2);
    CN145_sign_in(26) <= VN1409_sign_out(2);
    CN145_data_in(27) <= VN1442_data_out(2);
    CN145_sign_in(27) <= VN1442_sign_out(2);
    CN145_data_in(28) <= VN1460_data_out(2);
    CN145_sign_in(28) <= VN1460_sign_out(2);
    CN145_data_in(29) <= VN1492_data_out(2);
    CN145_sign_in(29) <= VN1492_sign_out(2);
    CN145_data_in(30) <= VN1669_data_out(2);
    CN145_sign_in(30) <= VN1669_sign_out(2);
    CN145_data_in(31) <= VN1759_data_out(2);
    CN145_sign_in(31) <= VN1759_sign_out(2);
    CN146_data_in(0) <= VN36_data_out(2);
    CN146_sign_in(0) <= VN36_sign_out(2);
    CN146_data_in(1) <= VN71_data_out(2);
    CN146_sign_in(1) <= VN71_sign_out(2);
    CN146_data_in(2) <= VN128_data_out(2);
    CN146_sign_in(2) <= VN128_sign_out(2);
    CN146_data_in(3) <= VN261_data_out(2);
    CN146_sign_in(3) <= VN261_sign_out(2);
    CN146_data_in(4) <= VN299_data_out(2);
    CN146_sign_in(4) <= VN299_sign_out(2);
    CN146_data_in(5) <= VN494_data_out(2);
    CN146_sign_in(5) <= VN494_sign_out(2);
    CN146_data_in(6) <= VN562_data_out(2);
    CN146_sign_in(6) <= VN562_sign_out(2);
    CN146_data_in(7) <= VN716_data_out(2);
    CN146_sign_in(7) <= VN716_sign_out(2);
    CN146_data_in(8) <= VN775_data_out(2);
    CN146_sign_in(8) <= VN775_sign_out(2);
    CN146_data_in(9) <= VN803_data_out(2);
    CN146_sign_in(9) <= VN803_sign_out(2);
    CN146_data_in(10) <= VN845_data_out(2);
    CN146_sign_in(10) <= VN845_sign_out(2);
    CN146_data_in(11) <= VN971_data_out(2);
    CN146_sign_in(11) <= VN971_sign_out(2);
    CN146_data_in(12) <= VN1011_data_out(2);
    CN146_sign_in(12) <= VN1011_sign_out(2);
    CN146_data_in(13) <= VN1266_data_out(2);
    CN146_sign_in(13) <= VN1266_sign_out(2);
    CN146_data_in(14) <= VN1316_data_out(2);
    CN146_sign_in(14) <= VN1316_sign_out(2);
    CN146_data_in(15) <= VN1457_data_out(2);
    CN146_sign_in(15) <= VN1457_sign_out(2);
    CN146_data_in(16) <= VN1496_data_out(2);
    CN146_sign_in(16) <= VN1496_sign_out(2);
    CN146_data_in(17) <= VN1535_data_out(2);
    CN146_sign_in(17) <= VN1535_sign_out(2);
    CN146_data_in(18) <= VN1545_data_out(2);
    CN146_sign_in(18) <= VN1545_sign_out(2);
    CN146_data_in(19) <= VN1646_data_out(2);
    CN146_sign_in(19) <= VN1646_sign_out(2);
    CN146_data_in(20) <= VN1654_data_out(2);
    CN146_sign_in(20) <= VN1654_sign_out(2);
    CN146_data_in(21) <= VN1689_data_out(2);
    CN146_sign_in(21) <= VN1689_sign_out(2);
    CN146_data_in(22) <= VN1854_data_out(2);
    CN146_sign_in(22) <= VN1854_sign_out(2);
    CN146_data_in(23) <= VN1890_data_out(2);
    CN146_sign_in(23) <= VN1890_sign_out(2);
    CN146_data_in(24) <= VN1946_data_out(2);
    CN146_sign_in(24) <= VN1946_sign_out(2);
    CN146_data_in(25) <= VN1948_data_out(2);
    CN146_sign_in(25) <= VN1948_sign_out(2);
    CN146_data_in(26) <= VN1972_data_out(2);
    CN146_sign_in(26) <= VN1972_sign_out(2);
    CN146_data_in(27) <= VN1980_data_out(2);
    CN146_sign_in(27) <= VN1980_sign_out(2);
    CN146_data_in(28) <= VN1991_data_out(2);
    CN146_sign_in(28) <= VN1991_sign_out(2);
    CN146_data_in(29) <= VN1997_data_out(2);
    CN146_sign_in(29) <= VN1997_sign_out(2);
    CN146_data_in(30) <= VN2032_data_out(2);
    CN146_sign_in(30) <= VN2032_sign_out(2);
    CN146_data_in(31) <= VN2039_data_out(2);
    CN146_sign_in(31) <= VN2039_sign_out(2);
    CN147_data_in(0) <= VN35_data_out(2);
    CN147_sign_in(0) <= VN35_sign_out(2);
    CN147_data_in(1) <= VN66_data_out(2);
    CN147_sign_in(1) <= VN66_sign_out(2);
    CN147_data_in(2) <= VN164_data_out(2);
    CN147_sign_in(2) <= VN164_sign_out(2);
    CN147_data_in(3) <= VN187_data_out(2);
    CN147_sign_in(3) <= VN187_sign_out(2);
    CN147_data_in(4) <= VN253_data_out(2);
    CN147_sign_in(4) <= VN253_sign_out(2);
    CN147_data_in(5) <= VN297_data_out(2);
    CN147_sign_in(5) <= VN297_sign_out(2);
    CN147_data_in(6) <= VN335_data_out(2);
    CN147_sign_in(6) <= VN335_sign_out(2);
    CN147_data_in(7) <= VN406_data_out(2);
    CN147_sign_in(7) <= VN406_sign_out(2);
    CN147_data_in(8) <= VN485_data_out(2);
    CN147_sign_in(8) <= VN485_sign_out(2);
    CN147_data_in(9) <= VN542_data_out(2);
    CN147_sign_in(9) <= VN542_sign_out(2);
    CN147_data_in(10) <= VN583_data_out(2);
    CN147_sign_in(10) <= VN583_sign_out(2);
    CN147_data_in(11) <= VN625_data_out(2);
    CN147_sign_in(11) <= VN625_sign_out(2);
    CN147_data_in(12) <= VN684_data_out(2);
    CN147_sign_in(12) <= VN684_sign_out(2);
    CN147_data_in(13) <= VN722_data_out(2);
    CN147_sign_in(13) <= VN722_sign_out(2);
    CN147_data_in(14) <= VN737_data_out(2);
    CN147_sign_in(14) <= VN737_sign_out(2);
    CN147_data_in(15) <= VN828_data_out(2);
    CN147_sign_in(15) <= VN828_sign_out(2);
    CN147_data_in(16) <= VN855_data_out(2);
    CN147_sign_in(16) <= VN855_sign_out(2);
    CN147_data_in(17) <= VN915_data_out(2);
    CN147_sign_in(17) <= VN915_sign_out(2);
    CN147_data_in(18) <= VN1026_data_out(2);
    CN147_sign_in(18) <= VN1026_sign_out(2);
    CN147_data_in(19) <= VN1081_data_out(2);
    CN147_sign_in(19) <= VN1081_sign_out(2);
    CN147_data_in(20) <= VN1118_data_out(2);
    CN147_sign_in(20) <= VN1118_sign_out(2);
    CN147_data_in(21) <= VN1215_data_out(2);
    CN147_sign_in(21) <= VN1215_sign_out(2);
    CN147_data_in(22) <= VN1268_data_out(2);
    CN147_sign_in(22) <= VN1268_sign_out(2);
    CN147_data_in(23) <= VN1285_data_out(2);
    CN147_sign_in(23) <= VN1285_sign_out(2);
    CN147_data_in(24) <= VN1373_data_out(2);
    CN147_sign_in(24) <= VN1373_sign_out(2);
    CN147_data_in(25) <= VN1489_data_out(2);
    CN147_sign_in(25) <= VN1489_sign_out(2);
    CN147_data_in(26) <= VN1567_data_out(2);
    CN147_sign_in(26) <= VN1567_sign_out(2);
    CN147_data_in(27) <= VN1600_data_out(2);
    CN147_sign_in(27) <= VN1600_sign_out(2);
    CN147_data_in(28) <= VN1739_data_out(2);
    CN147_sign_in(28) <= VN1739_sign_out(2);
    CN147_data_in(29) <= VN1752_data_out(2);
    CN147_sign_in(29) <= VN1752_sign_out(2);
    CN147_data_in(30) <= VN1807_data_out(2);
    CN147_sign_in(30) <= VN1807_sign_out(2);
    CN147_data_in(31) <= VN1836_data_out(2);
    CN147_sign_in(31) <= VN1836_sign_out(2);
    CN148_data_in(0) <= VN34_data_out(2);
    CN148_sign_in(0) <= VN34_sign_out(2);
    CN148_data_in(1) <= VN72_data_out(2);
    CN148_sign_in(1) <= VN72_sign_out(2);
    CN148_data_in(2) <= VN143_data_out(2);
    CN148_sign_in(2) <= VN143_sign_out(2);
    CN148_data_in(3) <= VN207_data_out(2);
    CN148_sign_in(3) <= VN207_sign_out(2);
    CN148_data_in(4) <= VN231_data_out(2);
    CN148_sign_in(4) <= VN231_sign_out(2);
    CN148_data_in(5) <= VN329_data_out(2);
    CN148_sign_in(5) <= VN329_sign_out(2);
    CN148_data_in(6) <= VN390_data_out(2);
    CN148_sign_in(6) <= VN390_sign_out(2);
    CN148_data_in(7) <= VN424_data_out(2);
    CN148_sign_in(7) <= VN424_sign_out(2);
    CN148_data_in(8) <= VN504_data_out(2);
    CN148_sign_in(8) <= VN504_sign_out(2);
    CN148_data_in(9) <= VN510_data_out(2);
    CN148_sign_in(9) <= VN510_sign_out(2);
    CN148_data_in(10) <= VN584_data_out(2);
    CN148_sign_in(10) <= VN584_sign_out(2);
    CN148_data_in(11) <= VN632_data_out(2);
    CN148_sign_in(11) <= VN632_sign_out(2);
    CN148_data_in(12) <= VN690_data_out(2);
    CN148_sign_in(12) <= VN690_sign_out(2);
    CN148_data_in(13) <= VN768_data_out(2);
    CN148_sign_in(13) <= VN768_sign_out(2);
    CN148_data_in(14) <= VN820_data_out(2);
    CN148_sign_in(14) <= VN820_sign_out(2);
    CN148_data_in(15) <= VN849_data_out(2);
    CN148_sign_in(15) <= VN849_sign_out(2);
    CN148_data_in(16) <= VN917_data_out(2);
    CN148_sign_in(16) <= VN917_sign_out(2);
    CN148_data_in(17) <= VN988_data_out(2);
    CN148_sign_in(17) <= VN988_sign_out(2);
    CN148_data_in(18) <= VN1046_data_out(2);
    CN148_sign_in(18) <= VN1046_sign_out(2);
    CN148_data_in(19) <= VN1104_data_out(2);
    CN148_sign_in(19) <= VN1104_sign_out(2);
    CN148_data_in(20) <= VN1198_data_out(2);
    CN148_sign_in(20) <= VN1198_sign_out(2);
    CN148_data_in(21) <= VN1238_data_out(2);
    CN148_sign_in(21) <= VN1238_sign_out(2);
    CN148_data_in(22) <= VN1308_data_out(2);
    CN148_sign_in(22) <= VN1308_sign_out(2);
    CN148_data_in(23) <= VN1331_data_out(2);
    CN148_sign_in(23) <= VN1331_sign_out(2);
    CN148_data_in(24) <= VN1335_data_out(2);
    CN148_sign_in(24) <= VN1335_sign_out(2);
    CN148_data_in(25) <= VN1424_data_out(2);
    CN148_sign_in(25) <= VN1424_sign_out(2);
    CN148_data_in(26) <= VN1435_data_out(2);
    CN148_sign_in(26) <= VN1435_sign_out(2);
    CN148_data_in(27) <= VN1510_data_out(2);
    CN148_sign_in(27) <= VN1510_sign_out(2);
    CN148_data_in(28) <= VN1589_data_out(2);
    CN148_sign_in(28) <= VN1589_sign_out(2);
    CN148_data_in(29) <= VN1640_data_out(2);
    CN148_sign_in(29) <= VN1640_sign_out(2);
    CN148_data_in(30) <= VN1803_data_out(2);
    CN148_sign_in(30) <= VN1803_sign_out(2);
    CN148_data_in(31) <= VN1837_data_out(2);
    CN148_sign_in(31) <= VN1837_sign_out(2);
    CN149_data_in(0) <= VN33_data_out(2);
    CN149_sign_in(0) <= VN33_sign_out(2);
    CN149_data_in(1) <= VN60_data_out(2);
    CN149_sign_in(1) <= VN60_sign_out(2);
    CN149_data_in(2) <= VN146_data_out(2);
    CN149_sign_in(2) <= VN146_sign_out(2);
    CN149_data_in(3) <= VN221_data_out(2);
    CN149_sign_in(3) <= VN221_sign_out(2);
    CN149_data_in(4) <= VN241_data_out(2);
    CN149_sign_in(4) <= VN241_sign_out(2);
    CN149_data_in(5) <= VN309_data_out(2);
    CN149_sign_in(5) <= VN309_sign_out(2);
    CN149_data_in(6) <= VN370_data_out(2);
    CN149_sign_in(6) <= VN370_sign_out(2);
    CN149_data_in(7) <= VN446_data_out(2);
    CN149_sign_in(7) <= VN446_sign_out(2);
    CN149_data_in(8) <= VN452_data_out(2);
    CN149_sign_in(8) <= VN452_sign_out(2);
    CN149_data_in(9) <= VN516_data_out(2);
    CN149_sign_in(9) <= VN516_sign_out(2);
    CN149_data_in(10) <= VN561_data_out(2);
    CN149_sign_in(10) <= VN561_sign_out(2);
    CN149_data_in(11) <= VN662_data_out(2);
    CN149_sign_in(11) <= VN662_sign_out(2);
    CN149_data_in(12) <= VN675_data_out(2);
    CN149_sign_in(12) <= VN675_sign_out(2);
    CN149_data_in(13) <= VN765_data_out(2);
    CN149_sign_in(13) <= VN765_sign_out(2);
    CN149_data_in(14) <= VN807_data_out(2);
    CN149_sign_in(14) <= VN807_sign_out(2);
    CN149_data_in(15) <= VN853_data_out(2);
    CN149_sign_in(15) <= VN853_sign_out(2);
    CN149_data_in(16) <= VN941_data_out(2);
    CN149_sign_in(16) <= VN941_sign_out(2);
    CN149_data_in(17) <= VN974_data_out(2);
    CN149_sign_in(17) <= VN974_sign_out(2);
    CN149_data_in(18) <= VN1056_data_out(2);
    CN149_sign_in(18) <= VN1056_sign_out(2);
    CN149_data_in(19) <= VN1096_data_out(2);
    CN149_sign_in(19) <= VN1096_sign_out(2);
    CN149_data_in(20) <= VN1131_data_out(2);
    CN149_sign_in(20) <= VN1131_sign_out(2);
    CN149_data_in(21) <= VN1210_data_out(2);
    CN149_sign_in(21) <= VN1210_sign_out(2);
    CN149_data_in(22) <= VN1275_data_out(2);
    CN149_sign_in(22) <= VN1275_sign_out(2);
    CN149_data_in(23) <= VN1296_data_out(2);
    CN149_sign_in(23) <= VN1296_sign_out(2);
    CN149_data_in(24) <= VN1354_data_out(2);
    CN149_sign_in(24) <= VN1354_sign_out(2);
    CN149_data_in(25) <= VN1403_data_out(2);
    CN149_sign_in(25) <= VN1403_sign_out(2);
    CN149_data_in(26) <= VN1454_data_out(2);
    CN149_sign_in(26) <= VN1454_sign_out(2);
    CN149_data_in(27) <= VN1462_data_out(2);
    CN149_sign_in(27) <= VN1462_sign_out(2);
    CN149_data_in(28) <= VN1473_data_out(2);
    CN149_sign_in(28) <= VN1473_sign_out(2);
    CN149_data_in(29) <= VN1624_data_out(2);
    CN149_sign_in(29) <= VN1624_sign_out(2);
    CN149_data_in(30) <= VN1726_data_out(2);
    CN149_sign_in(30) <= VN1726_sign_out(2);
    CN149_data_in(31) <= VN1838_data_out(2);
    CN149_sign_in(31) <= VN1838_sign_out(2);
    CN150_data_in(0) <= VN32_data_out(2);
    CN150_sign_in(0) <= VN32_sign_out(2);
    CN150_data_in(1) <= VN86_data_out(2);
    CN150_sign_in(1) <= VN86_sign_out(2);
    CN150_data_in(2) <= VN131_data_out(2);
    CN150_sign_in(2) <= VN131_sign_out(2);
    CN150_data_in(3) <= VN217_data_out(2);
    CN150_sign_in(3) <= VN217_sign_out(2);
    CN150_data_in(4) <= VN312_data_out(2);
    CN150_sign_in(4) <= VN312_sign_out(2);
    CN150_data_in(5) <= VN378_data_out(2);
    CN150_sign_in(5) <= VN378_sign_out(2);
    CN150_data_in(6) <= VN392_data_out(2);
    CN150_sign_in(6) <= VN392_sign_out(2);
    CN150_data_in(7) <= VN505_data_out(2);
    CN150_sign_in(7) <= VN505_sign_out(2);
    CN150_data_in(8) <= VN557_data_out(2);
    CN150_sign_in(8) <= VN557_sign_out(2);
    CN150_data_in(9) <= VN622_data_out(2);
    CN150_sign_in(9) <= VN622_sign_out(2);
    CN150_data_in(10) <= VN826_data_out(2);
    CN150_sign_in(10) <= VN826_sign_out(2);
    CN150_data_in(11) <= VN842_data_out(2);
    CN150_sign_in(11) <= VN842_sign_out(2);
    CN150_data_in(12) <= VN923_data_out(2);
    CN150_sign_in(12) <= VN923_sign_out(2);
    CN150_data_in(13) <= VN991_data_out(2);
    CN150_sign_in(13) <= VN991_sign_out(2);
    CN150_data_in(14) <= VN1051_data_out(2);
    CN150_sign_in(14) <= VN1051_sign_out(2);
    CN150_data_in(15) <= VN1086_data_out(2);
    CN150_sign_in(15) <= VN1086_sign_out(2);
    CN150_data_in(16) <= VN1138_data_out(2);
    CN150_sign_in(16) <= VN1138_sign_out(2);
    CN150_data_in(17) <= VN1216_data_out(2);
    CN150_sign_in(17) <= VN1216_sign_out(2);
    CN150_data_in(18) <= VN1231_data_out(2);
    CN150_sign_in(18) <= VN1231_sign_out(2);
    CN150_data_in(19) <= VN1276_data_out(2);
    CN150_sign_in(19) <= VN1276_sign_out(2);
    CN150_data_in(20) <= VN1318_data_out(2);
    CN150_sign_in(20) <= VN1318_sign_out(2);
    CN150_data_in(21) <= VN1362_data_out(2);
    CN150_sign_in(21) <= VN1362_sign_out(2);
    CN150_data_in(22) <= VN1388_data_out(2);
    CN150_sign_in(22) <= VN1388_sign_out(2);
    CN150_data_in(23) <= VN1602_data_out(2);
    CN150_sign_in(23) <= VN1602_sign_out(2);
    CN150_data_in(24) <= VN1749_data_out(2);
    CN150_sign_in(24) <= VN1749_sign_out(2);
    CN150_data_in(25) <= VN1805_data_out(2);
    CN150_sign_in(25) <= VN1805_sign_out(2);
    CN150_data_in(26) <= VN1847_data_out(2);
    CN150_sign_in(26) <= VN1847_sign_out(2);
    CN150_data_in(27) <= VN1858_data_out(2);
    CN150_sign_in(27) <= VN1858_sign_out(2);
    CN150_data_in(28) <= VN1859_data_out(2);
    CN150_sign_in(28) <= VN1859_sign_out(2);
    CN150_data_in(29) <= VN1911_data_out(2);
    CN150_sign_in(29) <= VN1911_sign_out(2);
    CN150_data_in(30) <= VN1925_data_out(2);
    CN150_sign_in(30) <= VN1925_sign_out(2);
    CN150_data_in(31) <= VN1930_data_out(2);
    CN150_sign_in(31) <= VN1930_sign_out(2);
    CN151_data_in(0) <= VN31_data_out(2);
    CN151_sign_in(0) <= VN31_sign_out(2);
    CN151_data_in(1) <= VN92_data_out(2);
    CN151_sign_in(1) <= VN92_sign_out(2);
    CN151_data_in(2) <= VN165_data_out(2);
    CN151_sign_in(2) <= VN165_sign_out(2);
    CN151_data_in(3) <= VN184_data_out(2);
    CN151_sign_in(3) <= VN184_sign_out(2);
    CN151_data_in(4) <= VN238_data_out(2);
    CN151_sign_in(4) <= VN238_sign_out(2);
    CN151_data_in(5) <= VN342_data_out(2);
    CN151_sign_in(5) <= VN342_sign_out(2);
    CN151_data_in(6) <= VN451_data_out(2);
    CN151_sign_in(6) <= VN451_sign_out(2);
    CN151_data_in(7) <= VN570_data_out(2);
    CN151_sign_in(7) <= VN570_sign_out(2);
    CN151_data_in(8) <= VN650_data_out(2);
    CN151_sign_in(8) <= VN650_sign_out(2);
    CN151_data_in(9) <= VN702_data_out(2);
    CN151_sign_in(9) <= VN702_sign_out(2);
    CN151_data_in(10) <= VN800_data_out(2);
    CN151_sign_in(10) <= VN800_sign_out(2);
    CN151_data_in(11) <= VN933_data_out(2);
    CN151_sign_in(11) <= VN933_sign_out(2);
    CN151_data_in(12) <= VN952_data_out(2);
    CN151_sign_in(12) <= VN952_sign_out(2);
    CN151_data_in(13) <= VN1057_data_out(2);
    CN151_sign_in(13) <= VN1057_sign_out(2);
    CN151_data_in(14) <= VN1110_data_out(2);
    CN151_sign_in(14) <= VN1110_sign_out(2);
    CN151_data_in(15) <= VN1192_data_out(2);
    CN151_sign_in(15) <= VN1192_sign_out(2);
    CN151_data_in(16) <= VN1239_data_out(2);
    CN151_sign_in(16) <= VN1239_sign_out(2);
    CN151_data_in(17) <= VN1547_data_out(2);
    CN151_sign_in(17) <= VN1547_sign_out(2);
    CN151_data_in(18) <= VN1562_data_out(2);
    CN151_sign_in(18) <= VN1562_sign_out(2);
    CN151_data_in(19) <= VN1619_data_out(2);
    CN151_sign_in(19) <= VN1619_sign_out(2);
    CN151_data_in(20) <= VN1667_data_out(2);
    CN151_sign_in(20) <= VN1667_sign_out(2);
    CN151_data_in(21) <= VN1714_data_out(2);
    CN151_sign_in(21) <= VN1714_sign_out(2);
    CN151_data_in(22) <= VN1822_data_out(2);
    CN151_sign_in(22) <= VN1822_sign_out(2);
    CN151_data_in(23) <= VN1864_data_out(2);
    CN151_sign_in(23) <= VN1864_sign_out(2);
    CN151_data_in(24) <= VN1867_data_out(2);
    CN151_sign_in(24) <= VN1867_sign_out(2);
    CN151_data_in(25) <= VN1912_data_out(2);
    CN151_sign_in(25) <= VN1912_sign_out(2);
    CN151_data_in(26) <= VN1950_data_out(2);
    CN151_sign_in(26) <= VN1950_sign_out(2);
    CN151_data_in(27) <= VN2021_data_out(2);
    CN151_sign_in(27) <= VN2021_sign_out(2);
    CN151_data_in(28) <= VN2029_data_out(2);
    CN151_sign_in(28) <= VN2029_sign_out(2);
    CN151_data_in(29) <= VN2031_data_out(2);
    CN151_sign_in(29) <= VN2031_sign_out(2);
    CN151_data_in(30) <= VN2034_data_out(2);
    CN151_sign_in(30) <= VN2034_sign_out(2);
    CN151_data_in(31) <= VN2041_data_out(2);
    CN151_sign_in(31) <= VN2041_sign_out(2);
    CN152_data_in(0) <= VN30_data_out(2);
    CN152_sign_in(0) <= VN30_sign_out(2);
    CN152_data_in(1) <= VN76_data_out(2);
    CN152_sign_in(1) <= VN76_sign_out(2);
    CN152_data_in(2) <= VN127_data_out(2);
    CN152_sign_in(2) <= VN127_sign_out(2);
    CN152_data_in(3) <= VN202_data_out(2);
    CN152_sign_in(3) <= VN202_sign_out(2);
    CN152_data_in(4) <= VN228_data_out(2);
    CN152_sign_in(4) <= VN228_sign_out(2);
    CN152_data_in(5) <= VN330_data_out(2);
    CN152_sign_in(5) <= VN330_sign_out(2);
    CN152_data_in(6) <= VN340_data_out(2);
    CN152_sign_in(6) <= VN340_sign_out(2);
    CN152_data_in(7) <= VN415_data_out(2);
    CN152_sign_in(7) <= VN415_sign_out(2);
    CN152_data_in(8) <= VN502_data_out(2);
    CN152_sign_in(8) <= VN502_sign_out(2);
    CN152_data_in(9) <= VN525_data_out(2);
    CN152_sign_in(9) <= VN525_sign_out(2);
    CN152_data_in(10) <= VN575_data_out(2);
    CN152_sign_in(10) <= VN575_sign_out(2);
    CN152_data_in(11) <= VN628_data_out(2);
    CN152_sign_in(11) <= VN628_sign_out(2);
    CN152_data_in(12) <= VN682_data_out(2);
    CN152_sign_in(12) <= VN682_sign_out(2);
    CN152_data_in(13) <= VN748_data_out(2);
    CN152_sign_in(13) <= VN748_sign_out(2);
    CN152_data_in(14) <= VN798_data_out(2);
    CN152_sign_in(14) <= VN798_sign_out(2);
    CN152_data_in(15) <= VN861_data_out(2);
    CN152_sign_in(15) <= VN861_sign_out(2);
    CN152_data_in(16) <= VN942_data_out(2);
    CN152_sign_in(16) <= VN942_sign_out(2);
    CN152_data_in(17) <= VN962_data_out(2);
    CN152_sign_in(17) <= VN962_sign_out(2);
    CN152_data_in(18) <= VN1045_data_out(2);
    CN152_sign_in(18) <= VN1045_sign_out(2);
    CN152_data_in(19) <= VN1079_data_out(2);
    CN152_sign_in(19) <= VN1079_sign_out(2);
    CN152_data_in(20) <= VN1123_data_out(2);
    CN152_sign_in(20) <= VN1123_sign_out(2);
    CN152_data_in(21) <= VN1205_data_out(2);
    CN152_sign_in(21) <= VN1205_sign_out(2);
    CN152_data_in(22) <= VN1267_data_out(2);
    CN152_sign_in(22) <= VN1267_sign_out(2);
    CN152_data_in(23) <= VN1300_data_out(2);
    CN152_sign_in(23) <= VN1300_sign_out(2);
    CN152_data_in(24) <= VN1363_data_out(2);
    CN152_sign_in(24) <= VN1363_sign_out(2);
    CN152_data_in(25) <= VN1390_data_out(2);
    CN152_sign_in(25) <= VN1390_sign_out(2);
    CN152_data_in(26) <= VN1458_data_out(2);
    CN152_sign_in(26) <= VN1458_sign_out(2);
    CN152_data_in(27) <= VN1543_data_out(2);
    CN152_sign_in(27) <= VN1543_sign_out(2);
    CN152_data_in(28) <= VN1711_data_out(2);
    CN152_sign_in(28) <= VN1711_sign_out(2);
    CN152_data_in(29) <= VN1742_data_out(2);
    CN152_sign_in(29) <= VN1742_sign_out(2);
    CN152_data_in(30) <= VN1802_data_out(2);
    CN152_sign_in(30) <= VN1802_sign_out(2);
    CN152_data_in(31) <= VN1839_data_out(2);
    CN152_sign_in(31) <= VN1839_sign_out(2);
    CN153_data_in(0) <= VN29_data_out(2);
    CN153_sign_in(0) <= VN29_sign_out(2);
    CN153_data_in(1) <= VN78_data_out(2);
    CN153_sign_in(1) <= VN78_sign_out(2);
    CN153_data_in(2) <= VN155_data_out(2);
    CN153_sign_in(2) <= VN155_sign_out(2);
    CN153_data_in(3) <= VN203_data_out(2);
    CN153_sign_in(3) <= VN203_sign_out(2);
    CN153_data_in(4) <= VN262_data_out(2);
    CN153_sign_in(4) <= VN262_sign_out(2);
    CN153_data_in(5) <= VN296_data_out(2);
    CN153_sign_in(5) <= VN296_sign_out(2);
    CN153_data_in(6) <= VN376_data_out(2);
    CN153_sign_in(6) <= VN376_sign_out(2);
    CN153_data_in(7) <= VN433_data_out(2);
    CN153_sign_in(7) <= VN433_sign_out(2);
    CN153_data_in(8) <= VN509_data_out(2);
    CN153_sign_in(8) <= VN509_sign_out(2);
    CN153_data_in(9) <= VN616_data_out(2);
    CN153_sign_in(9) <= VN616_sign_out(2);
    CN153_data_in(10) <= VN652_data_out(2);
    CN153_sign_in(10) <= VN652_sign_out(2);
    CN153_data_in(11) <= VN694_data_out(2);
    CN153_sign_in(11) <= VN694_sign_out(2);
    CN153_data_in(12) <= VN758_data_out(2);
    CN153_sign_in(12) <= VN758_sign_out(2);
    CN153_data_in(13) <= VN812_data_out(2);
    CN153_sign_in(13) <= VN812_sign_out(2);
    CN153_data_in(14) <= VN872_data_out(2);
    CN153_sign_in(14) <= VN872_sign_out(2);
    CN153_data_in(15) <= VN916_data_out(2);
    CN153_sign_in(15) <= VN916_sign_out(2);
    CN153_data_in(16) <= VN957_data_out(2);
    CN153_sign_in(16) <= VN957_sign_out(2);
    CN153_data_in(17) <= VN1077_data_out(2);
    CN153_sign_in(17) <= VN1077_sign_out(2);
    CN153_data_in(18) <= VN1149_data_out(2);
    CN153_sign_in(18) <= VN1149_sign_out(2);
    CN153_data_in(19) <= VN1178_data_out(2);
    CN153_sign_in(19) <= VN1178_sign_out(2);
    CN153_data_in(20) <= VN1226_data_out(2);
    CN153_sign_in(20) <= VN1226_sign_out(2);
    CN153_data_in(21) <= VN1314_data_out(2);
    CN153_sign_in(21) <= VN1314_sign_out(2);
    CN153_data_in(22) <= VN1353_data_out(2);
    CN153_sign_in(22) <= VN1353_sign_out(2);
    CN153_data_in(23) <= VN1398_data_out(2);
    CN153_sign_in(23) <= VN1398_sign_out(2);
    CN153_data_in(24) <= VN1437_data_out(2);
    CN153_sign_in(24) <= VN1437_sign_out(2);
    CN153_data_in(25) <= VN1484_data_out(2);
    CN153_sign_in(25) <= VN1484_sign_out(2);
    CN153_data_in(26) <= VN1553_data_out(2);
    CN153_sign_in(26) <= VN1553_sign_out(2);
    CN153_data_in(27) <= VN1587_data_out(2);
    CN153_sign_in(27) <= VN1587_sign_out(2);
    CN153_data_in(28) <= VN1651_data_out(2);
    CN153_sign_in(28) <= VN1651_sign_out(2);
    CN153_data_in(29) <= VN1699_data_out(2);
    CN153_sign_in(29) <= VN1699_sign_out(2);
    CN153_data_in(30) <= VN1729_data_out(2);
    CN153_sign_in(30) <= VN1729_sign_out(2);
    CN153_data_in(31) <= VN1840_data_out(2);
    CN153_sign_in(31) <= VN1840_sign_out(2);
    CN154_data_in(0) <= VN28_data_out(2);
    CN154_sign_in(0) <= VN28_sign_out(2);
    CN154_data_in(1) <= VN139_data_out(2);
    CN154_sign_in(1) <= VN139_sign_out(2);
    CN154_data_in(2) <= VN183_data_out(2);
    CN154_sign_in(2) <= VN183_sign_out(2);
    CN154_data_in(3) <= VN246_data_out(2);
    CN154_sign_in(3) <= VN246_sign_out(2);
    CN154_data_in(4) <= VN322_data_out(2);
    CN154_sign_in(4) <= VN322_sign_out(2);
    CN154_data_in(5) <= VN490_data_out(2);
    CN154_sign_in(5) <= VN490_sign_out(2);
    CN154_data_in(6) <= VN574_data_out(2);
    CN154_sign_in(6) <= VN574_sign_out(2);
    CN154_data_in(7) <= VN703_data_out(2);
    CN154_sign_in(7) <= VN703_sign_out(2);
    CN154_data_in(8) <= VN751_data_out(2);
    CN154_sign_in(8) <= VN751_sign_out(2);
    CN154_data_in(9) <= VN805_data_out(2);
    CN154_sign_in(9) <= VN805_sign_out(2);
    CN154_data_in(10) <= VN883_data_out(2);
    CN154_sign_in(10) <= VN883_sign_out(2);
    CN154_data_in(11) <= VN930_data_out(2);
    CN154_sign_in(11) <= VN930_sign_out(2);
    CN154_data_in(12) <= VN963_data_out(2);
    CN154_sign_in(12) <= VN963_sign_out(2);
    CN154_data_in(13) <= VN1020_data_out(2);
    CN154_sign_in(13) <= VN1020_sign_out(2);
    CN154_data_in(14) <= VN1166_data_out(2);
    CN154_sign_in(14) <= VN1166_sign_out(2);
    CN154_data_in(15) <= VN1254_data_out(2);
    CN154_sign_in(15) <= VN1254_sign_out(2);
    CN154_data_in(16) <= VN1376_data_out(2);
    CN154_sign_in(16) <= VN1376_sign_out(2);
    CN154_data_in(17) <= VN1420_data_out(2);
    CN154_sign_in(17) <= VN1420_sign_out(2);
    CN154_data_in(18) <= VN1434_data_out(2);
    CN154_sign_in(18) <= VN1434_sign_out(2);
    CN154_data_in(19) <= VN1584_data_out(2);
    CN154_sign_in(19) <= VN1584_sign_out(2);
    CN154_data_in(20) <= VN1642_data_out(2);
    CN154_sign_in(20) <= VN1642_sign_out(2);
    CN154_data_in(21) <= VN1685_data_out(2);
    CN154_sign_in(21) <= VN1685_sign_out(2);
    CN154_data_in(22) <= VN1706_data_out(2);
    CN154_sign_in(22) <= VN1706_sign_out(2);
    CN154_data_in(23) <= VN1855_data_out(2);
    CN154_sign_in(23) <= VN1855_sign_out(2);
    CN154_data_in(24) <= VN1868_data_out(2);
    CN154_sign_in(24) <= VN1868_sign_out(2);
    CN154_data_in(25) <= VN1891_data_out(2);
    CN154_sign_in(25) <= VN1891_sign_out(2);
    CN154_data_in(26) <= VN1942_data_out(2);
    CN154_sign_in(26) <= VN1942_sign_out(2);
    CN154_data_in(27) <= VN1999_data_out(2);
    CN154_sign_in(27) <= VN1999_sign_out(2);
    CN154_data_in(28) <= VN2013_data_out(2);
    CN154_sign_in(28) <= VN2013_sign_out(2);
    CN154_data_in(29) <= VN2015_data_out(2);
    CN154_sign_in(29) <= VN2015_sign_out(2);
    CN154_data_in(30) <= VN2045_data_out(2);
    CN154_sign_in(30) <= VN2045_sign_out(2);
    CN154_data_in(31) <= VN2046_data_out(2);
    CN154_sign_in(31) <= VN2046_sign_out(2);
    CN155_data_in(0) <= VN27_data_out(2);
    CN155_sign_in(0) <= VN27_sign_out(2);
    CN155_data_in(1) <= VN84_data_out(2);
    CN155_sign_in(1) <= VN84_sign_out(2);
    CN155_data_in(2) <= VN167_data_out(2);
    CN155_sign_in(2) <= VN167_sign_out(2);
    CN155_data_in(3) <= VN174_data_out(2);
    CN155_sign_in(3) <= VN174_sign_out(2);
    CN155_data_in(4) <= VN257_data_out(2);
    CN155_sign_in(4) <= VN257_sign_out(2);
    CN155_data_in(5) <= VN306_data_out(2);
    CN155_sign_in(5) <= VN306_sign_out(2);
    CN155_data_in(6) <= VN357_data_out(2);
    CN155_sign_in(6) <= VN357_sign_out(2);
    CN155_data_in(7) <= VN447_data_out(2);
    CN155_sign_in(7) <= VN447_sign_out(2);
    CN155_data_in(8) <= VN458_data_out(2);
    CN155_sign_in(8) <= VN458_sign_out(2);
    CN155_data_in(9) <= VN526_data_out(2);
    CN155_sign_in(9) <= VN526_sign_out(2);
    CN155_data_in(10) <= VN569_data_out(2);
    CN155_sign_in(10) <= VN569_sign_out(2);
    CN155_data_in(11) <= VN660_data_out(2);
    CN155_sign_in(11) <= VN660_sign_out(2);
    CN155_data_in(12) <= VN676_data_out(2);
    CN155_sign_in(12) <= VN676_sign_out(2);
    CN155_data_in(13) <= VN755_data_out(2);
    CN155_sign_in(13) <= VN755_sign_out(2);
    CN155_data_in(14) <= VN782_data_out(2);
    CN155_sign_in(14) <= VN782_sign_out(2);
    CN155_data_in(15) <= VN856_data_out(2);
    CN155_sign_in(15) <= VN856_sign_out(2);
    CN155_data_in(16) <= VN903_data_out(2);
    CN155_sign_in(16) <= VN903_sign_out(2);
    CN155_data_in(17) <= VN951_data_out(2);
    CN155_sign_in(17) <= VN951_sign_out(2);
    CN155_data_in(18) <= VN1005_data_out(2);
    CN155_sign_in(18) <= VN1005_sign_out(2);
    CN155_data_in(19) <= VN1083_data_out(2);
    CN155_sign_in(19) <= VN1083_sign_out(2);
    CN155_data_in(20) <= VN1141_data_out(2);
    CN155_sign_in(20) <= VN1141_sign_out(2);
    CN155_data_in(21) <= VN1180_data_out(2);
    CN155_sign_in(21) <= VN1180_sign_out(2);
    CN155_data_in(22) <= VN1234_data_out(2);
    CN155_sign_in(22) <= VN1234_sign_out(2);
    CN155_data_in(23) <= VN1290_data_out(2);
    CN155_sign_in(23) <= VN1290_sign_out(2);
    CN155_data_in(24) <= VN1329_data_out(2);
    CN155_sign_in(24) <= VN1329_sign_out(2);
    CN155_data_in(25) <= VN1382_data_out(2);
    CN155_sign_in(25) <= VN1382_sign_out(2);
    CN155_data_in(26) <= VN1421_data_out(2);
    CN155_sign_in(26) <= VN1421_sign_out(2);
    CN155_data_in(27) <= VN1456_data_out(2);
    CN155_sign_in(27) <= VN1456_sign_out(2);
    CN155_data_in(28) <= VN1595_data_out(2);
    CN155_sign_in(28) <= VN1595_sign_out(2);
    CN155_data_in(29) <= VN1657_data_out(2);
    CN155_sign_in(29) <= VN1657_sign_out(2);
    CN155_data_in(30) <= VN1702_data_out(2);
    CN155_sign_in(30) <= VN1702_sign_out(2);
    CN155_data_in(31) <= VN1760_data_out(2);
    CN155_sign_in(31) <= VN1760_sign_out(2);
    CN156_data_in(0) <= VN26_data_out(2);
    CN156_sign_in(0) <= VN26_sign_out(2);
    CN156_data_in(1) <= VN95_data_out(2);
    CN156_sign_in(1) <= VN95_sign_out(2);
    CN156_data_in(2) <= VN157_data_out(2);
    CN156_sign_in(2) <= VN157_sign_out(2);
    CN156_data_in(3) <= VN343_data_out(2);
    CN156_sign_in(3) <= VN343_sign_out(2);
    CN156_data_in(4) <= VN437_data_out(2);
    CN156_sign_in(4) <= VN437_sign_out(2);
    CN156_data_in(5) <= VN456_data_out(2);
    CN156_sign_in(5) <= VN456_sign_out(2);
    CN156_data_in(6) <= VN558_data_out(2);
    CN156_sign_in(6) <= VN558_sign_out(2);
    CN156_data_in(7) <= VN605_data_out(2);
    CN156_sign_in(7) <= VN605_sign_out(2);
    CN156_data_in(8) <= VN745_data_out(2);
    CN156_sign_in(8) <= VN745_sign_out(2);
    CN156_data_in(9) <= VN844_data_out(2);
    CN156_sign_in(9) <= VN844_sign_out(2);
    CN156_data_in(10) <= VN936_data_out(2);
    CN156_sign_in(10) <= VN936_sign_out(2);
    CN156_data_in(11) <= VN977_data_out(2);
    CN156_sign_in(11) <= VN977_sign_out(2);
    CN156_data_in(12) <= VN1003_data_out(2);
    CN156_sign_in(12) <= VN1003_sign_out(2);
    CN156_data_in(13) <= VN1006_data_out(2);
    CN156_sign_in(13) <= VN1006_sign_out(2);
    CN156_data_in(14) <= VN1150_data_out(2);
    CN156_sign_in(14) <= VN1150_sign_out(2);
    CN156_data_in(15) <= VN1255_data_out(2);
    CN156_sign_in(15) <= VN1255_sign_out(2);
    CN156_data_in(16) <= VN1303_data_out(2);
    CN156_sign_in(16) <= VN1303_sign_out(2);
    CN156_data_in(17) <= VN1366_data_out(2);
    CN156_sign_in(17) <= VN1366_sign_out(2);
    CN156_data_in(18) <= VN1397_data_out(2);
    CN156_sign_in(18) <= VN1397_sign_out(2);
    CN156_data_in(19) <= VN1508_data_out(2);
    CN156_sign_in(19) <= VN1508_sign_out(2);
    CN156_data_in(20) <= VN1644_data_out(2);
    CN156_sign_in(20) <= VN1644_sign_out(2);
    CN156_data_in(21) <= VN1661_data_out(2);
    CN156_sign_in(21) <= VN1661_sign_out(2);
    CN156_data_in(22) <= VN1728_data_out(2);
    CN156_sign_in(22) <= VN1728_sign_out(2);
    CN156_data_in(23) <= VN1789_data_out(2);
    CN156_sign_in(23) <= VN1789_sign_out(2);
    CN156_data_in(24) <= VN1913_data_out(2);
    CN156_sign_in(24) <= VN1913_sign_out(2);
    CN156_data_in(25) <= VN1921_data_out(2);
    CN156_sign_in(25) <= VN1921_sign_out(2);
    CN156_data_in(26) <= VN1936_data_out(2);
    CN156_sign_in(26) <= VN1936_sign_out(2);
    CN156_data_in(27) <= VN1971_data_out(2);
    CN156_sign_in(27) <= VN1971_sign_out(2);
    CN156_data_in(28) <= VN1975_data_out(2);
    CN156_sign_in(28) <= VN1975_sign_out(2);
    CN156_data_in(29) <= VN1984_data_out(2);
    CN156_sign_in(29) <= VN1984_sign_out(2);
    CN156_data_in(30) <= VN2019_data_out(2);
    CN156_sign_in(30) <= VN2019_sign_out(2);
    CN156_data_in(31) <= VN2022_data_out(2);
    CN156_sign_in(31) <= VN2022_sign_out(2);
    CN157_data_in(0) <= VN25_data_out(2);
    CN157_sign_in(0) <= VN25_sign_out(2);
    CN157_data_in(1) <= VN102_data_out(2);
    CN157_sign_in(1) <= VN102_sign_out(2);
    CN157_data_in(2) <= VN144_data_out(2);
    CN157_sign_in(2) <= VN144_sign_out(2);
    CN157_data_in(3) <= VN194_data_out(2);
    CN157_sign_in(3) <= VN194_sign_out(2);
    CN157_data_in(4) <= VN323_data_out(2);
    CN157_sign_in(4) <= VN323_sign_out(2);
    CN157_data_in(5) <= VN377_data_out(2);
    CN157_sign_in(5) <= VN377_sign_out(2);
    CN157_data_in(6) <= VN431_data_out(2);
    CN157_sign_in(6) <= VN431_sign_out(2);
    CN157_data_in(7) <= VN488_data_out(2);
    CN157_sign_in(7) <= VN488_sign_out(2);
    CN157_data_in(8) <= VN515_data_out(2);
    CN157_sign_in(8) <= VN515_sign_out(2);
    CN157_data_in(9) <= VN612_data_out(2);
    CN157_sign_in(9) <= VN612_sign_out(2);
    CN157_data_in(10) <= VN645_data_out(2);
    CN157_sign_in(10) <= VN645_sign_out(2);
    CN157_data_in(11) <= VN717_data_out(2);
    CN157_sign_in(11) <= VN717_sign_out(2);
    CN157_data_in(12) <= VN725_data_out(2);
    CN157_sign_in(12) <= VN725_sign_out(2);
    CN157_data_in(13) <= VN785_data_out(2);
    CN157_sign_in(13) <= VN785_sign_out(2);
    CN157_data_in(14) <= VN830_data_out(2);
    CN157_sign_in(14) <= VN830_sign_out(2);
    CN157_data_in(15) <= VN886_data_out(2);
    CN157_sign_in(15) <= VN886_sign_out(2);
    CN157_data_in(16) <= VN905_data_out(2);
    CN157_sign_in(16) <= VN905_sign_out(2);
    CN157_data_in(17) <= VN983_data_out(2);
    CN157_sign_in(17) <= VN983_sign_out(2);
    CN157_data_in(18) <= VN1029_data_out(2);
    CN157_sign_in(18) <= VN1029_sign_out(2);
    CN157_data_in(19) <= VN1069_data_out(2);
    CN157_sign_in(19) <= VN1069_sign_out(2);
    CN157_data_in(20) <= VN1122_data_out(2);
    CN157_sign_in(20) <= VN1122_sign_out(2);
    CN157_data_in(21) <= VN1190_data_out(2);
    CN157_sign_in(21) <= VN1190_sign_out(2);
    CN157_data_in(22) <= VN1269_data_out(2);
    CN157_sign_in(22) <= VN1269_sign_out(2);
    CN157_data_in(23) <= VN1297_data_out(2);
    CN157_sign_in(23) <= VN1297_sign_out(2);
    CN157_data_in(24) <= VN1368_data_out(2);
    CN157_sign_in(24) <= VN1368_sign_out(2);
    CN157_data_in(25) <= VN1384_data_out(2);
    CN157_sign_in(25) <= VN1384_sign_out(2);
    CN157_data_in(26) <= VN1392_data_out(2);
    CN157_sign_in(26) <= VN1392_sign_out(2);
    CN157_data_in(27) <= VN1477_data_out(2);
    CN157_sign_in(27) <= VN1477_sign_out(2);
    CN157_data_in(28) <= VN1612_data_out(2);
    CN157_sign_in(28) <= VN1612_sign_out(2);
    CN157_data_in(29) <= VN1687_data_out(2);
    CN157_sign_in(29) <= VN1687_sign_out(2);
    CN157_data_in(30) <= VN1696_data_out(2);
    CN157_sign_in(30) <= VN1696_sign_out(2);
    CN157_data_in(31) <= VN1761_data_out(2);
    CN157_sign_in(31) <= VN1761_sign_out(2);
    CN158_data_in(0) <= VN24_data_out(2);
    CN158_sign_in(0) <= VN24_sign_out(2);
    CN158_data_in(1) <= VN77_data_out(2);
    CN158_sign_in(1) <= VN77_sign_out(2);
    CN158_data_in(2) <= VN163_data_out(2);
    CN158_sign_in(2) <= VN163_sign_out(2);
    CN158_data_in(3) <= VN224_data_out(2);
    CN158_sign_in(3) <= VN224_sign_out(2);
    CN158_data_in(4) <= VN230_data_out(2);
    CN158_sign_in(4) <= VN230_sign_out(2);
    CN158_data_in(5) <= VN310_data_out(2);
    CN158_sign_in(5) <= VN310_sign_out(2);
    CN158_data_in(6) <= VN339_data_out(2);
    CN158_sign_in(6) <= VN339_sign_out(2);
    CN158_data_in(7) <= VN412_data_out(2);
    CN158_sign_in(7) <= VN412_sign_out(2);
    CN158_data_in(8) <= VN470_data_out(2);
    CN158_sign_in(8) <= VN470_sign_out(2);
    CN158_data_in(9) <= VN544_data_out(2);
    CN158_sign_in(9) <= VN544_sign_out(2);
    CN158_data_in(10) <= VN580_data_out(2);
    CN158_sign_in(10) <= VN580_sign_out(2);
    CN158_data_in(11) <= VN646_data_out(2);
    CN158_sign_in(11) <= VN646_sign_out(2);
    CN158_data_in(12) <= VN697_data_out(2);
    CN158_sign_in(12) <= VN697_sign_out(2);
    CN158_data_in(13) <= VN764_data_out(2);
    CN158_sign_in(13) <= VN764_sign_out(2);
    CN158_data_in(14) <= VN789_data_out(2);
    CN158_sign_in(14) <= VN789_sign_out(2);
    CN158_data_in(15) <= VN847_data_out(2);
    CN158_sign_in(15) <= VN847_sign_out(2);
    CN158_data_in(16) <= VN918_data_out(2);
    CN158_sign_in(16) <= VN918_sign_out(2);
    CN158_data_in(17) <= VN966_data_out(2);
    CN158_sign_in(17) <= VN966_sign_out(2);
    CN158_data_in(18) <= VN1012_data_out(2);
    CN158_sign_in(18) <= VN1012_sign_out(2);
    CN158_data_in(19) <= VN1063_data_out(2);
    CN158_sign_in(19) <= VN1063_sign_out(2);
    CN158_data_in(20) <= VN1137_data_out(2);
    CN158_sign_in(20) <= VN1137_sign_out(2);
    CN158_data_in(21) <= VN1208_data_out(2);
    CN158_sign_in(21) <= VN1208_sign_out(2);
    CN158_data_in(22) <= VN1218_data_out(2);
    CN158_sign_in(22) <= VN1218_sign_out(2);
    CN158_data_in(23) <= VN1265_data_out(2);
    CN158_sign_in(23) <= VN1265_sign_out(2);
    CN158_data_in(24) <= VN1326_data_out(2);
    CN158_sign_in(24) <= VN1326_sign_out(2);
    CN158_data_in(25) <= VN1337_data_out(2);
    CN158_sign_in(25) <= VN1337_sign_out(2);
    CN158_data_in(26) <= VN1407_data_out(2);
    CN158_sign_in(26) <= VN1407_sign_out(2);
    CN158_data_in(27) <= VN1475_data_out(2);
    CN158_sign_in(27) <= VN1475_sign_out(2);
    CN158_data_in(28) <= VN1578_data_out(2);
    CN158_sign_in(28) <= VN1578_sign_out(2);
    CN158_data_in(29) <= VN1621_data_out(2);
    CN158_sign_in(29) <= VN1621_sign_out(2);
    CN158_data_in(30) <= VN1660_data_out(2);
    CN158_sign_in(30) <= VN1660_sign_out(2);
    CN158_data_in(31) <= VN1762_data_out(2);
    CN158_sign_in(31) <= VN1762_sign_out(2);
    CN159_data_in(0) <= VN23_data_out(2);
    CN159_sign_in(0) <= VN23_sign_out(2);
    CN159_data_in(1) <= VN91_data_out(2);
    CN159_sign_in(1) <= VN91_sign_out(2);
    CN159_data_in(2) <= VN136_data_out(2);
    CN159_sign_in(2) <= VN136_sign_out(2);
    CN159_data_in(3) <= VN271_data_out(2);
    CN159_sign_in(3) <= VN271_sign_out(2);
    CN159_data_in(4) <= VN367_data_out(2);
    CN159_sign_in(4) <= VN367_sign_out(2);
    CN159_data_in(5) <= VN420_data_out(2);
    CN159_sign_in(5) <= VN420_sign_out(2);
    CN159_data_in(6) <= VN473_data_out(2);
    CN159_sign_in(6) <= VN473_sign_out(2);
    CN159_data_in(7) <= VN521_data_out(2);
    CN159_sign_in(7) <= VN521_sign_out(2);
    CN159_data_in(8) <= VN578_data_out(2);
    CN159_sign_in(8) <= VN578_sign_out(2);
    CN159_data_in(9) <= VN624_data_out(2);
    CN159_sign_in(9) <= VN624_sign_out(2);
    CN159_data_in(10) <= VN866_data_out(2);
    CN159_sign_in(10) <= VN866_sign_out(2);
    CN159_data_in(11) <= VN968_data_out(2);
    CN159_sign_in(11) <= VN968_sign_out(2);
    CN159_data_in(12) <= VN1023_data_out(2);
    CN159_sign_in(12) <= VN1023_sign_out(2);
    CN159_data_in(13) <= VN1067_data_out(2);
    CN159_sign_in(13) <= VN1067_sign_out(2);
    CN159_data_in(14) <= VN1113_data_out(2);
    CN159_sign_in(14) <= VN1113_sign_out(2);
    CN159_data_in(15) <= VN1229_data_out(2);
    CN159_sign_in(15) <= VN1229_sign_out(2);
    CN159_data_in(16) <= VN1374_data_out(2);
    CN159_sign_in(16) <= VN1374_sign_out(2);
    CN159_data_in(17) <= VN1481_data_out(2);
    CN159_sign_in(17) <= VN1481_sign_out(2);
    CN159_data_in(18) <= VN1512_data_out(2);
    CN159_sign_in(18) <= VN1512_sign_out(2);
    CN159_data_in(19) <= VN1616_data_out(2);
    CN159_sign_in(19) <= VN1616_sign_out(2);
    CN159_data_in(20) <= VN1735_data_out(2);
    CN159_sign_in(20) <= VN1735_sign_out(2);
    CN159_data_in(21) <= VN1755_data_out(2);
    CN159_sign_in(21) <= VN1755_sign_out(2);
    CN159_data_in(22) <= VN1775_data_out(2);
    CN159_sign_in(22) <= VN1775_sign_out(2);
    CN159_data_in(23) <= VN1900_data_out(2);
    CN159_sign_in(23) <= VN1900_sign_out(2);
    CN159_data_in(24) <= VN1951_data_out(2);
    CN159_sign_in(24) <= VN1951_sign_out(2);
    CN159_data_in(25) <= VN1956_data_out(2);
    CN159_sign_in(25) <= VN1956_sign_out(2);
    CN159_data_in(26) <= VN1958_data_out(2);
    CN159_sign_in(26) <= VN1958_sign_out(2);
    CN159_data_in(27) <= VN1967_data_out(2);
    CN159_sign_in(27) <= VN1967_sign_out(2);
    CN159_data_in(28) <= VN1969_data_out(2);
    CN159_sign_in(28) <= VN1969_sign_out(2);
    CN159_data_in(29) <= VN1974_data_out(2);
    CN159_sign_in(29) <= VN1974_sign_out(2);
    CN159_data_in(30) <= VN1985_data_out(2);
    CN159_sign_in(30) <= VN1985_sign_out(2);
    CN159_data_in(31) <= VN1987_data_out(2);
    CN159_sign_in(31) <= VN1987_sign_out(2);
    CN160_data_in(0) <= VN22_data_out(2);
    CN160_sign_in(0) <= VN22_sign_out(2);
    CN160_data_in(1) <= VN62_data_out(2);
    CN160_sign_in(1) <= VN62_sign_out(2);
    CN160_data_in(2) <= VN133_data_out(2);
    CN160_sign_in(2) <= VN133_sign_out(2);
    CN160_data_in(3) <= VN189_data_out(2);
    CN160_sign_in(3) <= VN189_sign_out(2);
    CN160_data_in(4) <= VN233_data_out(2);
    CN160_sign_in(4) <= VN233_sign_out(2);
    CN160_data_in(5) <= VN302_data_out(2);
    CN160_sign_in(5) <= VN302_sign_out(2);
    CN160_data_in(6) <= VN351_data_out(2);
    CN160_sign_in(6) <= VN351_sign_out(2);
    CN160_data_in(7) <= VN442_data_out(2);
    CN160_sign_in(7) <= VN442_sign_out(2);
    CN160_data_in(8) <= VN459_data_out(2);
    CN160_sign_in(8) <= VN459_sign_out(2);
    CN160_data_in(9) <= VN546_data_out(2);
    CN160_sign_in(9) <= VN546_sign_out(2);
    CN160_data_in(10) <= VN610_data_out(2);
    CN160_sign_in(10) <= VN610_sign_out(2);
    CN160_data_in(11) <= VN617_data_out(2);
    CN160_sign_in(11) <= VN617_sign_out(2);
    CN160_data_in(12) <= VN677_data_out(2);
    CN160_sign_in(12) <= VN677_sign_out(2);
    CN160_data_in(13) <= VN731_data_out(2);
    CN160_sign_in(13) <= VN731_sign_out(2);
    CN160_data_in(14) <= VN813_data_out(2);
    CN160_sign_in(14) <= VN813_sign_out(2);
    CN160_data_in(15) <= VN874_data_out(2);
    CN160_sign_in(15) <= VN874_sign_out(2);
    CN160_data_in(16) <= VN931_data_out(2);
    CN160_sign_in(16) <= VN931_sign_out(2);
    CN160_data_in(17) <= VN994_data_out(2);
    CN160_sign_in(17) <= VN994_sign_out(2);
    CN160_data_in(18) <= VN1030_data_out(2);
    CN160_sign_in(18) <= VN1030_sign_out(2);
    CN160_data_in(19) <= VN1109_data_out(2);
    CN160_sign_in(19) <= VN1109_sign_out(2);
    CN160_data_in(20) <= VN1144_data_out(2);
    CN160_sign_in(20) <= VN1144_sign_out(2);
    CN160_data_in(21) <= VN1175_data_out(2);
    CN160_sign_in(21) <= VN1175_sign_out(2);
    CN160_data_in(22) <= VN1249_data_out(2);
    CN160_sign_in(22) <= VN1249_sign_out(2);
    CN160_data_in(23) <= VN1443_data_out(2);
    CN160_sign_in(23) <= VN1443_sign_out(2);
    CN160_data_in(24) <= VN1527_data_out(2);
    CN160_sign_in(24) <= VN1527_sign_out(2);
    CN160_data_in(25) <= VN1534_data_out(2);
    CN160_sign_in(25) <= VN1534_sign_out(2);
    CN160_data_in(26) <= VN1552_data_out(2);
    CN160_sign_in(26) <= VN1552_sign_out(2);
    CN160_data_in(27) <= VN1565_data_out(2);
    CN160_sign_in(27) <= VN1565_sign_out(2);
    CN160_data_in(28) <= VN1576_data_out(2);
    CN160_sign_in(28) <= VN1576_sign_out(2);
    CN160_data_in(29) <= VN1622_data_out(2);
    CN160_sign_in(29) <= VN1622_sign_out(2);
    CN160_data_in(30) <= VN1683_data_out(2);
    CN160_sign_in(30) <= VN1683_sign_out(2);
    CN160_data_in(31) <= VN1763_data_out(2);
    CN160_sign_in(31) <= VN1763_sign_out(2);
    CN161_data_in(0) <= VN21_data_out(2);
    CN161_sign_in(0) <= VN21_sign_out(2);
    CN161_data_in(1) <= VN97_data_out(2);
    CN161_sign_in(1) <= VN97_sign_out(2);
    CN161_data_in(2) <= VN149_data_out(2);
    CN161_sign_in(2) <= VN149_sign_out(2);
    CN161_data_in(3) <= VN171_data_out(2);
    CN161_sign_in(3) <= VN171_sign_out(2);
    CN161_data_in(4) <= VN250_data_out(2);
    CN161_sign_in(4) <= VN250_sign_out(2);
    CN161_data_in(5) <= VN300_data_out(2);
    CN161_sign_in(5) <= VN300_sign_out(2);
    CN161_data_in(6) <= VN379_data_out(2);
    CN161_sign_in(6) <= VN379_sign_out(2);
    CN161_data_in(7) <= VN440_data_out(2);
    CN161_sign_in(7) <= VN440_sign_out(2);
    CN161_data_in(8) <= VN489_data_out(2);
    CN161_sign_in(8) <= VN489_sign_out(2);
    CN161_data_in(9) <= VN559_data_out(2);
    CN161_sign_in(9) <= VN559_sign_out(2);
    CN161_data_in(10) <= VN630_data_out(2);
    CN161_sign_in(10) <= VN630_sign_out(2);
    CN161_data_in(11) <= VN674_data_out(2);
    CN161_sign_in(11) <= VN674_sign_out(2);
    CN161_data_in(12) <= VN759_data_out(2);
    CN161_sign_in(12) <= VN759_sign_out(2);
    CN161_data_in(13) <= VN797_data_out(2);
    CN161_sign_in(13) <= VN797_sign_out(2);
    CN161_data_in(14) <= VN869_data_out(2);
    CN161_sign_in(14) <= VN869_sign_out(2);
    CN161_data_in(15) <= VN898_data_out(2);
    CN161_sign_in(15) <= VN898_sign_out(2);
    CN161_data_in(16) <= VN975_data_out(2);
    CN161_sign_in(16) <= VN975_sign_out(2);
    CN161_data_in(17) <= VN1207_data_out(2);
    CN161_sign_in(17) <= VN1207_sign_out(2);
    CN161_data_in(18) <= VN1250_data_out(2);
    CN161_sign_in(18) <= VN1250_sign_out(2);
    CN161_data_in(19) <= VN1411_data_out(2);
    CN161_sign_in(19) <= VN1411_sign_out(2);
    CN161_data_in(20) <= VN1452_data_out(2);
    CN161_sign_in(20) <= VN1452_sign_out(2);
    CN161_data_in(21) <= VN1531_data_out(2);
    CN161_sign_in(21) <= VN1531_sign_out(2);
    CN161_data_in(22) <= VN1570_data_out(2);
    CN161_sign_in(22) <= VN1570_sign_out(2);
    CN161_data_in(23) <= VN1650_data_out(2);
    CN161_sign_in(23) <= VN1650_sign_out(2);
    CN161_data_in(24) <= VN1743_data_out(2);
    CN161_sign_in(24) <= VN1743_sign_out(2);
    CN161_data_in(25) <= VN1745_data_out(2);
    CN161_sign_in(25) <= VN1745_sign_out(2);
    CN161_data_in(26) <= VN1784_data_out(2);
    CN161_sign_in(26) <= VN1784_sign_out(2);
    CN161_data_in(27) <= VN1790_data_out(2);
    CN161_sign_in(27) <= VN1790_sign_out(2);
    CN161_data_in(28) <= VN1823_data_out(2);
    CN161_sign_in(28) <= VN1823_sign_out(2);
    CN161_data_in(29) <= VN1830_data_out(2);
    CN161_sign_in(29) <= VN1830_sign_out(2);
    CN161_data_in(30) <= VN1861_data_out(2);
    CN161_sign_in(30) <= VN1861_sign_out(2);
    CN161_data_in(31) <= VN1882_data_out(2);
    CN161_sign_in(31) <= VN1882_sign_out(2);
    CN162_data_in(0) <= VN20_data_out(2);
    CN162_sign_in(0) <= VN20_sign_out(2);
    CN162_data_in(1) <= VN64_data_out(2);
    CN162_sign_in(1) <= VN64_sign_out(2);
    CN162_data_in(2) <= VN141_data_out(2);
    CN162_sign_in(2) <= VN141_sign_out(2);
    CN162_data_in(3) <= VN179_data_out(2);
    CN162_sign_in(3) <= VN179_sign_out(2);
    CN162_data_in(4) <= VN259_data_out(2);
    CN162_sign_in(4) <= VN259_sign_out(2);
    CN162_data_in(5) <= VN315_data_out(2);
    CN162_sign_in(5) <= VN315_sign_out(2);
    CN162_data_in(6) <= VN369_data_out(2);
    CN162_sign_in(6) <= VN369_sign_out(2);
    CN162_data_in(7) <= VN418_data_out(2);
    CN162_sign_in(7) <= VN418_sign_out(2);
    CN162_data_in(8) <= VN455_data_out(2);
    CN162_sign_in(8) <= VN455_sign_out(2);
    CN162_data_in(9) <= VN556_data_out(2);
    CN162_sign_in(9) <= VN556_sign_out(2);
    CN162_data_in(10) <= VN594_data_out(2);
    CN162_sign_in(10) <= VN594_sign_out(2);
    CN162_data_in(11) <= VN635_data_out(2);
    CN162_sign_in(11) <= VN635_sign_out(2);
    CN162_data_in(12) <= VN692_data_out(2);
    CN162_sign_in(12) <= VN692_sign_out(2);
    CN162_data_in(13) <= VN747_data_out(2);
    CN162_sign_in(13) <= VN747_sign_out(2);
    CN162_data_in(14) <= VN808_data_out(2);
    CN162_sign_in(14) <= VN808_sign_out(2);
    CN162_data_in(15) <= VN875_data_out(2);
    CN162_sign_in(15) <= VN875_sign_out(2);
    CN162_data_in(16) <= VN899_data_out(2);
    CN162_sign_in(16) <= VN899_sign_out(2);
    CN162_data_in(17) <= VN987_data_out(2);
    CN162_sign_in(17) <= VN987_sign_out(2);
    CN162_data_in(18) <= VN1019_data_out(2);
    CN162_sign_in(18) <= VN1019_sign_out(2);
    CN162_data_in(19) <= VN1076_data_out(2);
    CN162_sign_in(19) <= VN1076_sign_out(2);
    CN162_data_in(20) <= VN1124_data_out(2);
    CN162_sign_in(20) <= VN1124_sign_out(2);
    CN162_data_in(21) <= VN1228_data_out(2);
    CN162_sign_in(21) <= VN1228_sign_out(2);
    CN162_data_in(22) <= VN1323_data_out(2);
    CN162_sign_in(22) <= VN1323_sign_out(2);
    CN162_data_in(23) <= VN1367_data_out(2);
    CN162_sign_in(23) <= VN1367_sign_out(2);
    CN162_data_in(24) <= VN1405_data_out(2);
    CN162_sign_in(24) <= VN1405_sign_out(2);
    CN162_data_in(25) <= VN1446_data_out(2);
    CN162_sign_in(25) <= VN1446_sign_out(2);
    CN162_data_in(26) <= VN1575_data_out(2);
    CN162_sign_in(26) <= VN1575_sign_out(2);
    CN162_data_in(27) <= VN1632_data_out(2);
    CN162_sign_in(27) <= VN1632_sign_out(2);
    CN162_data_in(28) <= VN1664_data_out(2);
    CN162_sign_in(28) <= VN1664_sign_out(2);
    CN162_data_in(29) <= VN1725_data_out(2);
    CN162_sign_in(29) <= VN1725_sign_out(2);
    CN162_data_in(30) <= VN1919_data_out(2);
    CN162_sign_in(30) <= VN1919_sign_out(2);
    CN162_data_in(31) <= VN1923_data_out(2);
    CN162_sign_in(31) <= VN1923_sign_out(2);
    CN163_data_in(0) <= VN19_data_out(2);
    CN163_sign_in(0) <= VN19_sign_out(2);
    CN163_data_in(1) <= VN79_data_out(2);
    CN163_sign_in(1) <= VN79_sign_out(2);
    CN163_data_in(2) <= VN115_data_out(2);
    CN163_sign_in(2) <= VN115_sign_out(2);
    CN163_data_in(3) <= VN254_data_out(2);
    CN163_sign_in(3) <= VN254_sign_out(2);
    CN163_data_in(4) <= VN355_data_out(2);
    CN163_sign_in(4) <= VN355_sign_out(2);
    CN163_data_in(5) <= VN399_data_out(2);
    CN163_sign_in(5) <= VN399_sign_out(2);
    CN163_data_in(6) <= VN481_data_out(2);
    CN163_sign_in(6) <= VN481_sign_out(2);
    CN163_data_in(7) <= VN517_data_out(2);
    CN163_sign_in(7) <= VN517_sign_out(2);
    CN163_data_in(8) <= VN581_data_out(2);
    CN163_sign_in(8) <= VN581_sign_out(2);
    CN163_data_in(9) <= VN668_data_out(2);
    CN163_sign_in(9) <= VN668_sign_out(2);
    CN163_data_in(10) <= VN734_data_out(2);
    CN163_sign_in(10) <= VN734_sign_out(2);
    CN163_data_in(11) <= VN865_data_out(2);
    CN163_sign_in(11) <= VN865_sign_out(2);
    CN163_data_in(12) <= VN995_data_out(2);
    CN163_sign_in(12) <= VN995_sign_out(2);
    CN163_data_in(13) <= VN1047_data_out(2);
    CN163_sign_in(13) <= VN1047_sign_out(2);
    CN163_data_in(14) <= VN1087_data_out(2);
    CN163_sign_in(14) <= VN1087_sign_out(2);
    CN163_data_in(15) <= VN1121_data_out(2);
    CN163_sign_in(15) <= VN1121_sign_out(2);
    CN163_data_in(16) <= VN1381_data_out(2);
    CN163_sign_in(16) <= VN1381_sign_out(2);
    CN163_data_in(17) <= VN1550_data_out(2);
    CN163_sign_in(17) <= VN1550_sign_out(2);
    CN163_data_in(18) <= VN1569_data_out(2);
    CN163_sign_in(18) <= VN1569_sign_out(2);
    CN163_data_in(19) <= VN1637_data_out(2);
    CN163_sign_in(19) <= VN1637_sign_out(2);
    CN163_data_in(20) <= VN1663_data_out(2);
    CN163_sign_in(20) <= VN1663_sign_out(2);
    CN163_data_in(21) <= VN1698_data_out(2);
    CN163_sign_in(21) <= VN1698_sign_out(2);
    CN163_data_in(22) <= VN1801_data_out(2);
    CN163_sign_in(22) <= VN1801_sign_out(2);
    CN163_data_in(23) <= VN1874_data_out(2);
    CN163_sign_in(23) <= VN1874_sign_out(2);
    CN163_data_in(24) <= VN1896_data_out(2);
    CN163_sign_in(24) <= VN1896_sign_out(2);
    CN163_data_in(25) <= VN1907_data_out(2);
    CN163_sign_in(25) <= VN1907_sign_out(2);
    CN163_data_in(26) <= VN1915_data_out(2);
    CN163_sign_in(26) <= VN1915_sign_out(2);
    CN163_data_in(27) <= VN1960_data_out(2);
    CN163_sign_in(27) <= VN1960_sign_out(2);
    CN163_data_in(28) <= VN1976_data_out(2);
    CN163_sign_in(28) <= VN1976_sign_out(2);
    CN163_data_in(29) <= VN1979_data_out(2);
    CN163_sign_in(29) <= VN1979_sign_out(2);
    CN163_data_in(30) <= VN2006_data_out(2);
    CN163_sign_in(30) <= VN2006_sign_out(2);
    CN163_data_in(31) <= VN2011_data_out(2);
    CN163_sign_in(31) <= VN2011_sign_out(2);
    CN164_data_in(0) <= VN18_data_out(2);
    CN164_sign_in(0) <= VN18_sign_out(2);
    CN164_data_in(1) <= VN75_data_out(2);
    CN164_sign_in(1) <= VN75_sign_out(2);
    CN164_data_in(2) <= VN125_data_out(2);
    CN164_sign_in(2) <= VN125_sign_out(2);
    CN164_data_in(3) <= VN197_data_out(2);
    CN164_sign_in(3) <= VN197_sign_out(2);
    CN164_data_in(4) <= VN260_data_out(2);
    CN164_sign_in(4) <= VN260_sign_out(2);
    CN164_data_in(5) <= VN375_data_out(2);
    CN164_sign_in(5) <= VN375_sign_out(2);
    CN164_data_in(6) <= VN401_data_out(2);
    CN164_sign_in(6) <= VN401_sign_out(2);
    CN164_data_in(7) <= VN539_data_out(2);
    CN164_sign_in(7) <= VN539_sign_out(2);
    CN164_data_in(8) <= VN611_data_out(2);
    CN164_sign_in(8) <= VN611_sign_out(2);
    CN164_data_in(9) <= VN634_data_out(2);
    CN164_sign_in(9) <= VN634_sign_out(2);
    CN164_data_in(10) <= VN714_data_out(2);
    CN164_sign_in(10) <= VN714_sign_out(2);
    CN164_data_in(11) <= VN749_data_out(2);
    CN164_sign_in(11) <= VN749_sign_out(2);
    CN164_data_in(12) <= VN792_data_out(2);
    CN164_sign_in(12) <= VN792_sign_out(2);
    CN164_data_in(13) <= VN833_data_out(2);
    CN164_sign_in(13) <= VN833_sign_out(2);
    CN164_data_in(14) <= VN924_data_out(2);
    CN164_sign_in(14) <= VN924_sign_out(2);
    CN164_data_in(15) <= VN967_data_out(2);
    CN164_sign_in(15) <= VN967_sign_out(2);
    CN164_data_in(16) <= VN1025_data_out(2);
    CN164_sign_in(16) <= VN1025_sign_out(2);
    CN164_data_in(17) <= VN1095_data_out(2);
    CN164_sign_in(17) <= VN1095_sign_out(2);
    CN164_data_in(18) <= VN1139_data_out(2);
    CN164_sign_in(18) <= VN1139_sign_out(2);
    CN164_data_in(19) <= VN1237_data_out(2);
    CN164_sign_in(19) <= VN1237_sign_out(2);
    CN164_data_in(20) <= VN1289_data_out(2);
    CN164_sign_in(20) <= VN1289_sign_out(2);
    CN164_data_in(21) <= VN1394_data_out(2);
    CN164_sign_in(21) <= VN1394_sign_out(2);
    CN164_data_in(22) <= VN1494_data_out(2);
    CN164_sign_in(22) <= VN1494_sign_out(2);
    CN164_data_in(23) <= VN1516_data_out(2);
    CN164_sign_in(23) <= VN1516_sign_out(2);
    CN164_data_in(24) <= VN1557_data_out(2);
    CN164_sign_in(24) <= VN1557_sign_out(2);
    CN164_data_in(25) <= VN1563_data_out(2);
    CN164_sign_in(25) <= VN1563_sign_out(2);
    CN164_data_in(26) <= VN1690_data_out(2);
    CN164_sign_in(26) <= VN1690_sign_out(2);
    CN164_data_in(27) <= VN1732_data_out(2);
    CN164_sign_in(27) <= VN1732_sign_out(2);
    CN164_data_in(28) <= VN1826_data_out(2);
    CN164_sign_in(28) <= VN1826_sign_out(2);
    CN164_data_in(29) <= VN1897_data_out(2);
    CN164_sign_in(29) <= VN1897_sign_out(2);
    CN164_data_in(30) <= VN1914_data_out(2);
    CN164_sign_in(30) <= VN1914_sign_out(2);
    CN164_data_in(31) <= VN1916_data_out(2);
    CN164_sign_in(31) <= VN1916_sign_out(2);
    CN165_data_in(0) <= VN17_data_out(2);
    CN165_sign_in(0) <= VN17_sign_out(2);
    CN165_data_in(1) <= VN93_data_out(2);
    CN165_sign_in(1) <= VN93_sign_out(2);
    CN165_data_in(2) <= VN119_data_out(2);
    CN165_sign_in(2) <= VN119_sign_out(2);
    CN165_data_in(3) <= VN177_data_out(2);
    CN165_sign_in(3) <= VN177_sign_out(2);
    CN165_data_in(4) <= VN294_data_out(2);
    CN165_sign_in(4) <= VN294_sign_out(2);
    CN165_data_in(5) <= VN348_data_out(2);
    CN165_sign_in(5) <= VN348_sign_out(2);
    CN165_data_in(6) <= VN443_data_out(2);
    CN165_sign_in(6) <= VN443_sign_out(2);
    CN165_data_in(7) <= VN491_data_out(2);
    CN165_sign_in(7) <= VN491_sign_out(2);
    CN165_data_in(8) <= VN540_data_out(2);
    CN165_sign_in(8) <= VN540_sign_out(2);
    CN165_data_in(9) <= VN629_data_out(2);
    CN165_sign_in(9) <= VN629_sign_out(2);
    CN165_data_in(10) <= VN691_data_out(2);
    CN165_sign_in(10) <= VN691_sign_out(2);
    CN165_data_in(11) <= VN769_data_out(2);
    CN165_sign_in(11) <= VN769_sign_out(2);
    CN165_data_in(12) <= VN781_data_out(2);
    CN165_sign_in(12) <= VN781_sign_out(2);
    CN165_data_in(13) <= VN839_data_out(2);
    CN165_sign_in(13) <= VN839_sign_out(2);
    CN165_data_in(14) <= VN940_data_out(2);
    CN165_sign_in(14) <= VN940_sign_out(2);
    CN165_data_in(15) <= VN982_data_out(2);
    CN165_sign_in(15) <= VN982_sign_out(2);
    CN165_data_in(16) <= VN1049_data_out(2);
    CN165_sign_in(16) <= VN1049_sign_out(2);
    CN165_data_in(17) <= VN1070_data_out(2);
    CN165_sign_in(17) <= VN1070_sign_out(2);
    CN165_data_in(18) <= VN1162_data_out(2);
    CN165_sign_in(18) <= VN1162_sign_out(2);
    CN165_data_in(19) <= VN1219_data_out(2);
    CN165_sign_in(19) <= VN1219_sign_out(2);
    CN165_data_in(20) <= VN1416_data_out(2);
    CN165_sign_in(20) <= VN1416_sign_out(2);
    CN165_data_in(21) <= VN1440_data_out(2);
    CN165_sign_in(21) <= VN1440_sign_out(2);
    CN165_data_in(22) <= VN1519_data_out(2);
    CN165_sign_in(22) <= VN1519_sign_out(2);
    CN165_data_in(23) <= VN1601_data_out(2);
    CN165_sign_in(23) <= VN1601_sign_out(2);
    CN165_data_in(24) <= VN1701_data_out(2);
    CN165_sign_in(24) <= VN1701_sign_out(2);
    CN165_data_in(25) <= VN1780_data_out(2);
    CN165_sign_in(25) <= VN1780_sign_out(2);
    CN165_data_in(26) <= VN1806_data_out(2);
    CN165_sign_in(26) <= VN1806_sign_out(2);
    CN165_data_in(27) <= VN1811_data_out(2);
    CN165_sign_in(27) <= VN1811_sign_out(2);
    CN165_data_in(28) <= VN1906_data_out(2);
    CN165_sign_in(28) <= VN1906_sign_out(2);
    CN165_data_in(29) <= VN1917_data_out(2);
    CN165_sign_in(29) <= VN1917_sign_out(2);
    CN165_data_in(30) <= VN2018_data_out(2);
    CN165_sign_in(30) <= VN2018_sign_out(2);
    CN165_data_in(31) <= VN2026_data_out(2);
    CN165_sign_in(31) <= VN2026_sign_out(2);
    CN166_data_in(0) <= VN16_data_out(2);
    CN166_sign_in(0) <= VN16_sign_out(2);
    CN166_data_in(1) <= VN57_data_out(2);
    CN166_sign_in(1) <= VN57_sign_out(2);
    CN166_data_in(2) <= VN122_data_out(2);
    CN166_sign_in(2) <= VN122_sign_out(2);
    CN166_data_in(3) <= VN210_data_out(2);
    CN166_sign_in(3) <= VN210_sign_out(2);
    CN166_data_in(4) <= VN288_data_out(2);
    CN166_sign_in(4) <= VN288_sign_out(2);
    CN166_data_in(5) <= VN345_data_out(2);
    CN166_sign_in(5) <= VN345_sign_out(2);
    CN166_data_in(6) <= VN419_data_out(2);
    CN166_sign_in(6) <= VN419_sign_out(2);
    CN166_data_in(7) <= VN483_data_out(2);
    CN166_sign_in(7) <= VN483_sign_out(2);
    CN166_data_in(8) <= VN667_data_out(2);
    CN166_sign_in(8) <= VN667_sign_out(2);
    CN166_data_in(9) <= VN683_data_out(2);
    CN166_sign_in(9) <= VN683_sign_out(2);
    CN166_data_in(10) <= VN723_data_out(2);
    CN166_sign_in(10) <= VN723_sign_out(2);
    CN166_data_in(11) <= VN777_data_out(2);
    CN166_sign_in(11) <= VN777_sign_out(2);
    CN166_data_in(12) <= VN822_data_out(2);
    CN166_sign_in(12) <= VN822_sign_out(2);
    CN166_data_in(13) <= VN878_data_out(2);
    CN166_sign_in(13) <= VN878_sign_out(2);
    CN166_data_in(14) <= VN888_data_out(2);
    CN166_sign_in(14) <= VN888_sign_out(2);
    CN166_data_in(15) <= VN953_data_out(2);
    CN166_sign_in(15) <= VN953_sign_out(2);
    CN166_data_in(16) <= VN1007_data_out(2);
    CN166_sign_in(16) <= VN1007_sign_out(2);
    CN166_data_in(17) <= VN1111_data_out(2);
    CN166_sign_in(17) <= VN1111_sign_out(2);
    CN166_data_in(18) <= VN1163_data_out(2);
    CN166_sign_in(18) <= VN1163_sign_out(2);
    CN166_data_in(19) <= VN1309_data_out(2);
    CN166_sign_in(19) <= VN1309_sign_out(2);
    CN166_data_in(20) <= VN1356_data_out(2);
    CN166_sign_in(20) <= VN1356_sign_out(2);
    CN166_data_in(21) <= VN1415_data_out(2);
    CN166_sign_in(21) <= VN1415_sign_out(2);
    CN166_data_in(22) <= VN1471_data_out(2);
    CN166_sign_in(22) <= VN1471_sign_out(2);
    CN166_data_in(23) <= VN1515_data_out(2);
    CN166_sign_in(23) <= VN1515_sign_out(2);
    CN166_data_in(24) <= VN1525_data_out(2);
    CN166_sign_in(24) <= VN1525_sign_out(2);
    CN166_data_in(25) <= VN1579_data_out(2);
    CN166_sign_in(25) <= VN1579_sign_out(2);
    CN166_data_in(26) <= VN1673_data_out(2);
    CN166_sign_in(26) <= VN1673_sign_out(2);
    CN166_data_in(27) <= VN1709_data_out(2);
    CN166_sign_in(27) <= VN1709_sign_out(2);
    CN166_data_in(28) <= VN1808_data_out(2);
    CN166_sign_in(28) <= VN1808_sign_out(2);
    CN166_data_in(29) <= VN1862_data_out(2);
    CN166_sign_in(29) <= VN1862_sign_out(2);
    CN166_data_in(30) <= VN1863_data_out(2);
    CN166_sign_in(30) <= VN1863_sign_out(2);
    CN166_data_in(31) <= VN1883_data_out(2);
    CN166_sign_in(31) <= VN1883_sign_out(2);
    CN167_data_in(0) <= VN15_data_out(2);
    CN167_sign_in(0) <= VN15_sign_out(2);
    CN167_data_in(1) <= VN58_data_out(2);
    CN167_sign_in(1) <= VN58_sign_out(2);
    CN167_data_in(2) <= VN112_data_out(2);
    CN167_sign_in(2) <= VN112_sign_out(2);
    CN167_data_in(3) <= VN213_data_out(2);
    CN167_sign_in(3) <= VN213_sign_out(2);
    CN167_data_in(4) <= VN225_data_out(2);
    CN167_sign_in(4) <= VN225_sign_out(2);
    CN167_data_in(5) <= VN292_data_out(2);
    CN167_sign_in(5) <= VN292_sign_out(2);
    CN167_data_in(6) <= VN360_data_out(2);
    CN167_sign_in(6) <= VN360_sign_out(2);
    CN167_data_in(7) <= VN471_data_out(2);
    CN167_sign_in(7) <= VN471_sign_out(2);
    CN167_data_in(8) <= VN588_data_out(2);
    CN167_sign_in(8) <= VN588_sign_out(2);
    CN167_data_in(9) <= VN701_data_out(2);
    CN167_sign_in(9) <= VN701_sign_out(2);
    CN167_data_in(10) <= VN773_data_out(2);
    CN167_sign_in(10) <= VN773_sign_out(2);
    CN167_data_in(11) <= VN784_data_out(2);
    CN167_sign_in(11) <= VN784_sign_out(2);
    CN167_data_in(12) <= VN880_data_out(2);
    CN167_sign_in(12) <= VN880_sign_out(2);
    CN167_data_in(13) <= VN990_data_out(2);
    CN167_sign_in(13) <= VN990_sign_out(2);
    CN167_data_in(14) <= VN1004_data_out(2);
    CN167_sign_in(14) <= VN1004_sign_out(2);
    CN167_data_in(15) <= VN1167_data_out(2);
    CN167_sign_in(15) <= VN1167_sign_out(2);
    CN167_data_in(16) <= VN1214_data_out(2);
    CN167_sign_in(16) <= VN1214_sign_out(2);
    CN167_data_in(17) <= VN1240_data_out(2);
    CN167_sign_in(17) <= VN1240_sign_out(2);
    CN167_data_in(18) <= VN1369_data_out(2);
    CN167_sign_in(18) <= VN1369_sign_out(2);
    CN167_data_in(19) <= VN1393_data_out(2);
    CN167_sign_in(19) <= VN1393_sign_out(2);
    CN167_data_in(20) <= VN1502_data_out(2);
    CN167_sign_in(20) <= VN1502_sign_out(2);
    CN167_data_in(21) <= VN1574_data_out(2);
    CN167_sign_in(21) <= VN1574_sign_out(2);
    CN167_data_in(22) <= VN1630_data_out(2);
    CN167_sign_in(22) <= VN1630_sign_out(2);
    CN167_data_in(23) <= VN1665_data_out(2);
    CN167_sign_in(23) <= VN1665_sign_out(2);
    CN167_data_in(24) <= VN1791_data_out(2);
    CN167_sign_in(24) <= VN1791_sign_out(2);
    CN167_data_in(25) <= VN1895_data_out(2);
    CN167_sign_in(25) <= VN1895_sign_out(2);
    CN167_data_in(26) <= VN1927_data_out(2);
    CN167_sign_in(26) <= VN1927_sign_out(2);
    CN167_data_in(27) <= VN1990_data_out(2);
    CN167_sign_in(27) <= VN1990_sign_out(2);
    CN167_data_in(28) <= VN2030_data_out(2);
    CN167_sign_in(28) <= VN2030_sign_out(2);
    CN167_data_in(29) <= VN2035_data_out(2);
    CN167_sign_in(29) <= VN2035_sign_out(2);
    CN167_data_in(30) <= VN2037_data_out(2);
    CN167_sign_in(30) <= VN2037_sign_out(2);
    CN167_data_in(31) <= VN2043_data_out(2);
    CN167_sign_in(31) <= VN2043_sign_out(2);
    CN168_data_in(0) <= VN14_data_out(2);
    CN168_sign_in(0) <= VN14_sign_out(2);
    CN168_data_in(1) <= VN150_data_out(2);
    CN168_sign_in(1) <= VN150_sign_out(2);
    CN168_data_in(2) <= VN199_data_out(2);
    CN168_sign_in(2) <= VN199_sign_out(2);
    CN168_data_in(3) <= VN264_data_out(2);
    CN168_sign_in(3) <= VN264_sign_out(2);
    CN168_data_in(4) <= VN283_data_out(2);
    CN168_sign_in(4) <= VN283_sign_out(2);
    CN168_data_in(5) <= VN353_data_out(2);
    CN168_sign_in(5) <= VN353_sign_out(2);
    CN168_data_in(6) <= VN409_data_out(2);
    CN168_sign_in(6) <= VN409_sign_out(2);
    CN168_data_in(7) <= VN487_data_out(2);
    CN168_sign_in(7) <= VN487_sign_out(2);
    CN168_data_in(8) <= VN524_data_out(2);
    CN168_sign_in(8) <= VN524_sign_out(2);
    CN168_data_in(9) <= VN613_data_out(2);
    CN168_sign_in(9) <= VN613_sign_out(2);
    CN168_data_in(10) <= VN641_data_out(2);
    CN168_sign_in(10) <= VN641_sign_out(2);
    CN168_data_in(11) <= VN705_data_out(2);
    CN168_sign_in(11) <= VN705_sign_out(2);
    CN168_data_in(12) <= VN724_data_out(2);
    CN168_sign_in(12) <= VN724_sign_out(2);
    CN168_data_in(13) <= VN801_data_out(2);
    CN168_sign_in(13) <= VN801_sign_out(2);
    CN168_data_in(14) <= VN851_data_out(2);
    CN168_sign_in(14) <= VN851_sign_out(2);
    CN168_data_in(15) <= VN943_data_out(2);
    CN168_sign_in(15) <= VN943_sign_out(2);
    CN168_data_in(16) <= VN955_data_out(2);
    CN168_sign_in(16) <= VN955_sign_out(2);
    CN168_data_in(17) <= VN1021_data_out(2);
    CN168_sign_in(17) <= VN1021_sign_out(2);
    CN168_data_in(18) <= VN1061_data_out(2);
    CN168_sign_in(18) <= VN1061_sign_out(2);
    CN168_data_in(19) <= VN1130_data_out(2);
    CN168_sign_in(19) <= VN1130_sign_out(2);
    CN168_data_in(20) <= VN1196_data_out(2);
    CN168_sign_in(20) <= VN1196_sign_out(2);
    CN168_data_in(21) <= VN1235_data_out(2);
    CN168_sign_in(21) <= VN1235_sign_out(2);
    CN168_data_in(22) <= VN1277_data_out(2);
    CN168_sign_in(22) <= VN1277_sign_out(2);
    CN168_data_in(23) <= VN1325_data_out(2);
    CN168_sign_in(23) <= VN1325_sign_out(2);
    CN168_data_in(24) <= VN1365_data_out(2);
    CN168_sign_in(24) <= VN1365_sign_out(2);
    CN168_data_in(25) <= VN1603_data_out(2);
    CN168_sign_in(25) <= VN1603_sign_out(2);
    CN168_data_in(26) <= VN1641_data_out(2);
    CN168_sign_in(26) <= VN1641_sign_out(2);
    CN168_data_in(27) <= VN1649_data_out(2);
    CN168_sign_in(27) <= VN1649_sign_out(2);
    CN168_data_in(28) <= VN1734_data_out(2);
    CN168_sign_in(28) <= VN1734_sign_out(2);
    CN168_data_in(29) <= VN1786_data_out(2);
    CN168_sign_in(29) <= VN1786_sign_out(2);
    CN168_data_in(30) <= VN1996_data_out(2);
    CN168_sign_in(30) <= VN1996_sign_out(2);
    CN168_data_in(31) <= VN2000_data_out(2);
    CN168_sign_in(31) <= VN2000_sign_out(2);
    CN169_data_in(0) <= VN13_data_out(2);
    CN169_sign_in(0) <= VN13_sign_out(2);
    CN169_data_in(1) <= VN85_data_out(2);
    CN169_sign_in(1) <= VN85_sign_out(2);
    CN169_data_in(2) <= VN132_data_out(2);
    CN169_sign_in(2) <= VN132_sign_out(2);
    CN169_data_in(3) <= VN178_data_out(2);
    CN169_sign_in(3) <= VN178_sign_out(2);
    CN169_data_in(4) <= VN266_data_out(2);
    CN169_sign_in(4) <= VN266_sign_out(2);
    CN169_data_in(5) <= VN316_data_out(2);
    CN169_sign_in(5) <= VN316_sign_out(2);
    CN169_data_in(6) <= VN387_data_out(2);
    CN169_sign_in(6) <= VN387_sign_out(2);
    CN169_data_in(7) <= VN395_data_out(2);
    CN169_sign_in(7) <= VN395_sign_out(2);
    CN169_data_in(8) <= VN529_data_out(2);
    CN169_sign_in(8) <= VN529_sign_out(2);
    CN169_data_in(9) <= VN604_data_out(2);
    CN169_sign_in(9) <= VN604_sign_out(2);
    CN169_data_in(10) <= VN639_data_out(2);
    CN169_sign_in(10) <= VN639_sign_out(2);
    CN169_data_in(11) <= VN810_data_out(2);
    CN169_sign_in(11) <= VN810_sign_out(2);
    CN169_data_in(12) <= VN831_data_out(2);
    CN169_sign_in(12) <= VN831_sign_out(2);
    CN169_data_in(13) <= VN938_data_out(2);
    CN169_sign_in(13) <= VN938_sign_out(2);
    CN169_data_in(14) <= VN969_data_out(2);
    CN169_sign_in(14) <= VN969_sign_out(2);
    CN169_data_in(15) <= VN1042_data_out(2);
    CN169_sign_in(15) <= VN1042_sign_out(2);
    CN169_data_in(16) <= VN1148_data_out(2);
    CN169_sign_in(16) <= VN1148_sign_out(2);
    CN169_data_in(17) <= VN1203_data_out(2);
    CN169_sign_in(17) <= VN1203_sign_out(2);
    CN169_data_in(18) <= VN1273_data_out(2);
    CN169_sign_in(18) <= VN1273_sign_out(2);
    CN169_data_in(19) <= VN1311_data_out(2);
    CN169_sign_in(19) <= VN1311_sign_out(2);
    CN169_data_in(20) <= VN1453_data_out(2);
    CN169_sign_in(20) <= VN1453_sign_out(2);
    CN169_data_in(21) <= VN1469_data_out(2);
    CN169_sign_in(21) <= VN1469_sign_out(2);
    CN169_data_in(22) <= VN1479_data_out(2);
    CN169_sign_in(22) <= VN1479_sign_out(2);
    CN169_data_in(23) <= VN1488_data_out(2);
    CN169_sign_in(23) <= VN1488_sign_out(2);
    CN169_data_in(24) <= VN1498_data_out(2);
    CN169_sign_in(24) <= VN1498_sign_out(2);
    CN169_data_in(25) <= VN1539_data_out(2);
    CN169_sign_in(25) <= VN1539_sign_out(2);
    CN169_data_in(26) <= VN1713_data_out(2);
    CN169_sign_in(26) <= VN1713_sign_out(2);
    CN169_data_in(27) <= VN1751_data_out(2);
    CN169_sign_in(27) <= VN1751_sign_out(2);
    CN169_data_in(28) <= VN1819_data_out(2);
    CN169_sign_in(28) <= VN1819_sign_out(2);
    CN169_data_in(29) <= VN1961_data_out(2);
    CN169_sign_in(29) <= VN1961_sign_out(2);
    CN169_data_in(30) <= VN1962_data_out(2);
    CN169_sign_in(30) <= VN1962_sign_out(2);
    CN169_data_in(31) <= VN1977_data_out(2);
    CN169_sign_in(31) <= VN1977_sign_out(2);
    CN170_data_in(0) <= VN12_data_out(2);
    CN170_sign_in(0) <= VN12_sign_out(2);
    CN170_data_in(1) <= VN101_data_out(2);
    CN170_sign_in(1) <= VN101_sign_out(2);
    CN170_data_in(2) <= VN145_data_out(2);
    CN170_sign_in(2) <= VN145_sign_out(2);
    CN170_data_in(3) <= VN236_data_out(2);
    CN170_sign_in(3) <= VN236_sign_out(2);
    CN170_data_in(4) <= VN337_data_out(2);
    CN170_sign_in(4) <= VN337_sign_out(2);
    CN170_data_in(5) <= VN421_data_out(2);
    CN170_sign_in(5) <= VN421_sign_out(2);
    CN170_data_in(6) <= VN461_data_out(2);
    CN170_sign_in(6) <= VN461_sign_out(2);
    CN170_data_in(7) <= VN592_data_out(2);
    CN170_sign_in(7) <= VN592_sign_out(2);
    CN170_data_in(8) <= VN620_data_out(2);
    CN170_sign_in(8) <= VN620_sign_out(2);
    CN170_data_in(9) <= VN843_data_out(2);
    CN170_sign_in(9) <= VN843_sign_out(2);
    CN170_data_in(10) <= VN965_data_out(2);
    CN170_sign_in(10) <= VN965_sign_out(2);
    CN170_data_in(11) <= VN1043_data_out(2);
    CN170_sign_in(11) <= VN1043_sign_out(2);
    CN170_data_in(12) <= VN1088_data_out(2);
    CN170_sign_in(12) <= VN1088_sign_out(2);
    CN170_data_in(13) <= VN1153_data_out(2);
    CN170_sign_in(13) <= VN1153_sign_out(2);
    CN170_data_in(14) <= VN1171_data_out(2);
    CN170_sign_in(14) <= VN1171_sign_out(2);
    CN170_data_in(15) <= VN1328_data_out(2);
    CN170_sign_in(15) <= VN1328_sign_out(2);
    CN170_data_in(16) <= VN1350_data_out(2);
    CN170_sign_in(16) <= VN1350_sign_out(2);
    CN170_data_in(17) <= VN1417_data_out(2);
    CN170_sign_in(17) <= VN1417_sign_out(2);
    CN170_data_in(18) <= VN1497_data_out(2);
    CN170_sign_in(18) <= VN1497_sign_out(2);
    CN170_data_in(19) <= VN1524_data_out(2);
    CN170_sign_in(19) <= VN1524_sign_out(2);
    CN170_data_in(20) <= VN1588_data_out(2);
    CN170_sign_in(20) <= VN1588_sign_out(2);
    CN170_data_in(21) <= VN1626_data_out(2);
    CN170_sign_in(21) <= VN1626_sign_out(2);
    CN170_data_in(22) <= VN1681_data_out(2);
    CN170_sign_in(22) <= VN1681_sign_out(2);
    CN170_data_in(23) <= VN1800_data_out(2);
    CN170_sign_in(23) <= VN1800_sign_out(2);
    CN170_data_in(24) <= VN1804_data_out(2);
    CN170_sign_in(24) <= VN1804_sign_out(2);
    CN170_data_in(25) <= VN1898_data_out(2);
    CN170_sign_in(25) <= VN1898_sign_out(2);
    CN170_data_in(26) <= VN1924_data_out(2);
    CN170_sign_in(26) <= VN1924_sign_out(2);
    CN170_data_in(27) <= VN1959_data_out(2);
    CN170_sign_in(27) <= VN1959_sign_out(2);
    CN170_data_in(28) <= VN1986_data_out(2);
    CN170_sign_in(28) <= VN1986_sign_out(2);
    CN170_data_in(29) <= VN1993_data_out(2);
    CN170_sign_in(29) <= VN1993_sign_out(2);
    CN170_data_in(30) <= VN2020_data_out(2);
    CN170_sign_in(30) <= VN2020_sign_out(2);
    CN170_data_in(31) <= VN2025_data_out(2);
    CN170_sign_in(31) <= VN2025_sign_out(2);
    CN171_data_in(0) <= VN105_data_out(2);
    CN171_sign_in(0) <= VN105_sign_out(2);
    CN171_data_in(1) <= VN156_data_out(2);
    CN171_sign_in(1) <= VN156_sign_out(2);
    CN171_data_in(2) <= VN222_data_out(2);
    CN171_sign_in(2) <= VN222_sign_out(2);
    CN171_data_in(3) <= VN311_data_out(2);
    CN171_sign_in(3) <= VN311_sign_out(2);
    CN171_data_in(4) <= VN411_data_out(2);
    CN171_sign_in(4) <= VN411_sign_out(2);
    CN171_data_in(5) <= VN476_data_out(2);
    CN171_sign_in(5) <= VN476_sign_out(2);
    CN171_data_in(6) <= VN528_data_out(2);
    CN171_sign_in(6) <= VN528_sign_out(2);
    CN171_data_in(7) <= VN609_data_out(2);
    CN171_sign_in(7) <= VN609_sign_out(2);
    CN171_data_in(8) <= VN699_data_out(2);
    CN171_sign_in(8) <= VN699_sign_out(2);
    CN171_data_in(9) <= VN743_data_out(2);
    CN171_sign_in(9) <= VN743_sign_out(2);
    CN171_data_in(10) <= VN811_data_out(2);
    CN171_sign_in(10) <= VN811_sign_out(2);
    CN171_data_in(11) <= VN852_data_out(2);
    CN171_sign_in(11) <= VN852_sign_out(2);
    CN171_data_in(12) <= VN928_data_out(2);
    CN171_sign_in(12) <= VN928_sign_out(2);
    CN171_data_in(13) <= VN985_data_out(2);
    CN171_sign_in(13) <= VN985_sign_out(2);
    CN171_data_in(14) <= VN1084_data_out(2);
    CN171_sign_in(14) <= VN1084_sign_out(2);
    CN171_data_in(15) <= VN1245_data_out(2);
    CN171_sign_in(15) <= VN1245_sign_out(2);
    CN171_data_in(16) <= VN1279_data_out(2);
    CN171_sign_in(16) <= VN1279_sign_out(2);
    CN171_data_in(17) <= VN1294_data_out(2);
    CN171_sign_in(17) <= VN1294_sign_out(2);
    CN171_data_in(18) <= VN1351_data_out(2);
    CN171_sign_in(18) <= VN1351_sign_out(2);
    CN171_data_in(19) <= VN1430_data_out(2);
    CN171_sign_in(19) <= VN1430_sign_out(2);
    CN171_data_in(20) <= VN1514_data_out(2);
    CN171_sign_in(20) <= VN1514_sign_out(2);
    CN171_data_in(21) <= VN1518_data_out(2);
    CN171_sign_in(21) <= VN1518_sign_out(2);
    CN171_data_in(22) <= VN1593_data_out(2);
    CN171_sign_in(22) <= VN1593_sign_out(2);
    CN171_data_in(23) <= VN1692_data_out(2);
    CN171_sign_in(23) <= VN1692_sign_out(2);
    CN171_data_in(24) <= VN1730_data_out(2);
    CN171_sign_in(24) <= VN1730_sign_out(2);
    CN171_data_in(25) <= VN1798_data_out(2);
    CN171_sign_in(25) <= VN1798_sign_out(2);
    CN171_data_in(26) <= VN1857_data_out(2);
    CN171_sign_in(26) <= VN1857_sign_out(2);
    CN171_data_in(27) <= VN1889_data_out(2);
    CN171_sign_in(27) <= VN1889_sign_out(2);
    CN171_data_in(28) <= VN1892_data_out(2);
    CN171_sign_in(28) <= VN1892_sign_out(2);
    CN171_data_in(29) <= VN1922_data_out(2);
    CN171_sign_in(29) <= VN1922_sign_out(2);
    CN171_data_in(30) <= VN1933_data_out(2);
    CN171_sign_in(30) <= VN1933_sign_out(2);
    CN171_data_in(31) <= VN1937_data_out(2);
    CN171_sign_in(31) <= VN1937_sign_out(2);
    CN172_data_in(0) <= VN11_data_out(2);
    CN172_sign_in(0) <= VN11_sign_out(2);
    CN172_data_in(1) <= VN110_data_out(2);
    CN172_sign_in(1) <= VN110_sign_out(2);
    CN172_data_in(2) <= VN126_data_out(2);
    CN172_sign_in(2) <= VN126_sign_out(2);
    CN172_data_in(3) <= VN229_data_out(2);
    CN172_sign_in(3) <= VN229_sign_out(2);
    CN172_data_in(4) <= VN400_data_out(2);
    CN172_sign_in(4) <= VN400_sign_out(2);
    CN172_data_in(5) <= VN468_data_out(2);
    CN172_sign_in(5) <= VN468_sign_out(2);
    CN172_data_in(6) <= VN523_data_out(2);
    CN172_sign_in(6) <= VN523_sign_out(2);
    CN172_data_in(7) <= VN585_data_out(2);
    CN172_sign_in(7) <= VN585_sign_out(2);
    CN172_data_in(8) <= VN655_data_out(2);
    CN172_sign_in(8) <= VN655_sign_out(2);
    CN172_data_in(9) <= VN727_data_out(2);
    CN172_sign_in(9) <= VN727_sign_out(2);
    CN172_data_in(10) <= VN879_data_out(2);
    CN172_sign_in(10) <= VN879_sign_out(2);
    CN172_data_in(11) <= VN894_data_out(2);
    CN172_sign_in(11) <= VN894_sign_out(2);
    CN172_data_in(12) <= VN948_data_out(2);
    CN172_sign_in(12) <= VN948_sign_out(2);
    CN172_data_in(13) <= VN1013_data_out(2);
    CN172_sign_in(13) <= VN1013_sign_out(2);
    CN172_data_in(14) <= VN1089_data_out(2);
    CN172_sign_in(14) <= VN1089_sign_out(2);
    CN172_data_in(15) <= VN1152_data_out(2);
    CN172_sign_in(15) <= VN1152_sign_out(2);
    CN172_data_in(16) <= VN1201_data_out(2);
    CN172_sign_in(16) <= VN1201_sign_out(2);
    CN172_data_in(17) <= VN1243_data_out(2);
    CN172_sign_in(17) <= VN1243_sign_out(2);
    CN172_data_in(18) <= VN1383_data_out(2);
    CN172_sign_in(18) <= VN1383_sign_out(2);
    CN172_data_in(19) <= VN1414_data_out(2);
    CN172_sign_in(19) <= VN1414_sign_out(2);
    CN172_data_in(20) <= VN1591_data_out(2);
    CN172_sign_in(20) <= VN1591_sign_out(2);
    CN172_data_in(21) <= VN1613_data_out(2);
    CN172_sign_in(21) <= VN1613_sign_out(2);
    CN172_data_in(22) <= VN1754_data_out(2);
    CN172_sign_in(22) <= VN1754_sign_out(2);
    CN172_data_in(23) <= VN1795_data_out(2);
    CN172_sign_in(23) <= VN1795_sign_out(2);
    CN172_data_in(24) <= VN1866_data_out(2);
    CN172_sign_in(24) <= VN1866_sign_out(2);
    CN172_data_in(25) <= VN1875_data_out(2);
    CN172_sign_in(25) <= VN1875_sign_out(2);
    CN172_data_in(26) <= VN1908_data_out(2);
    CN172_sign_in(26) <= VN1908_sign_out(2);
    CN172_data_in(27) <= VN1957_data_out(2);
    CN172_sign_in(27) <= VN1957_sign_out(2);
    CN172_data_in(28) <= VN1983_data_out(2);
    CN172_sign_in(28) <= VN1983_sign_out(2);
    CN172_data_in(29) <= VN2009_data_out(2);
    CN172_sign_in(29) <= VN2009_sign_out(2);
    CN172_data_in(30) <= VN2027_data_out(2);
    CN172_sign_in(30) <= VN2027_sign_out(2);
    CN172_data_in(31) <= VN2033_data_out(2);
    CN172_sign_in(31) <= VN2033_sign_out(2);
    CN173_data_in(0) <= VN10_data_out(2);
    CN173_sign_in(0) <= VN10_sign_out(2);
    CN173_data_in(1) <= VN104_data_out(2);
    CN173_sign_in(1) <= VN104_sign_out(2);
    CN173_data_in(2) <= VN114_data_out(2);
    CN173_sign_in(2) <= VN114_sign_out(2);
    CN173_data_in(3) <= VN180_data_out(2);
    CN173_sign_in(3) <= VN180_sign_out(2);
    CN173_data_in(4) <= VN237_data_out(2);
    CN173_sign_in(4) <= VN237_sign_out(2);
    CN173_data_in(5) <= VN295_data_out(2);
    CN173_sign_in(5) <= VN295_sign_out(2);
    CN173_data_in(6) <= VN384_data_out(2);
    CN173_sign_in(6) <= VN384_sign_out(2);
    CN173_data_in(7) <= VN417_data_out(2);
    CN173_sign_in(7) <= VN417_sign_out(2);
    CN173_data_in(8) <= VN499_data_out(2);
    CN173_sign_in(8) <= VN499_sign_out(2);
    CN173_data_in(9) <= VN642_data_out(2);
    CN173_sign_in(9) <= VN642_sign_out(2);
    CN173_data_in(10) <= VN688_data_out(2);
    CN173_sign_in(10) <= VN688_sign_out(2);
    CN173_data_in(11) <= VN729_data_out(2);
    CN173_sign_in(11) <= VN729_sign_out(2);
    CN173_data_in(12) <= VN825_data_out(2);
    CN173_sign_in(12) <= VN825_sign_out(2);
    CN173_data_in(13) <= VN838_data_out(2);
    CN173_sign_in(13) <= VN838_sign_out(2);
    CN173_data_in(14) <= VN892_data_out(2);
    CN173_sign_in(14) <= VN892_sign_out(2);
    CN173_data_in(15) <= VN949_data_out(2);
    CN173_sign_in(15) <= VN949_sign_out(2);
    CN173_data_in(16) <= VN1060_data_out(2);
    CN173_sign_in(16) <= VN1060_sign_out(2);
    CN173_data_in(17) <= VN1146_data_out(2);
    CN173_sign_in(17) <= VN1146_sign_out(2);
    CN173_data_in(18) <= VN1183_data_out(2);
    CN173_sign_in(18) <= VN1183_sign_out(2);
    CN173_data_in(19) <= VN1298_data_out(2);
    CN173_sign_in(19) <= VN1298_sign_out(2);
    CN173_data_in(20) <= VN1375_data_out(2);
    CN173_sign_in(20) <= VN1375_sign_out(2);
    CN173_data_in(21) <= VN1470_data_out(2);
    CN173_sign_in(21) <= VN1470_sign_out(2);
    CN173_data_in(22) <= VN1522_data_out(2);
    CN173_sign_in(22) <= VN1522_sign_out(2);
    CN173_data_in(23) <= VN1594_data_out(2);
    CN173_sign_in(23) <= VN1594_sign_out(2);
    CN173_data_in(24) <= VN1682_data_out(2);
    CN173_sign_in(24) <= VN1682_sign_out(2);
    CN173_data_in(25) <= VN1716_data_out(2);
    CN173_sign_in(25) <= VN1716_sign_out(2);
    CN173_data_in(26) <= VN1727_data_out(2);
    CN173_sign_in(26) <= VN1727_sign_out(2);
    CN173_data_in(27) <= VN1820_data_out(2);
    CN173_sign_in(27) <= VN1820_sign_out(2);
    CN173_data_in(28) <= VN1829_data_out(2);
    CN173_sign_in(28) <= VN1829_sign_out(2);
    CN173_data_in(29) <= VN1853_data_out(2);
    CN173_sign_in(29) <= VN1853_sign_out(2);
    CN173_data_in(30) <= VN1934_data_out(2);
    CN173_sign_in(30) <= VN1934_sign_out(2);
    CN173_data_in(31) <= VN1944_data_out(2);
    CN173_sign_in(31) <= VN1944_sign_out(2);
    CN174_data_in(0) <= VN9_data_out(2);
    CN174_sign_in(0) <= VN9_sign_out(2);
    CN174_data_in(1) <= VN99_data_out(2);
    CN174_sign_in(1) <= VN99_sign_out(2);
    CN174_data_in(2) <= VN159_data_out(2);
    CN174_sign_in(2) <= VN159_sign_out(2);
    CN174_data_in(3) <= VN265_data_out(2);
    CN174_sign_in(3) <= VN265_sign_out(2);
    CN174_data_in(4) <= VN361_data_out(2);
    CN174_sign_in(4) <= VN361_sign_out(2);
    CN174_data_in(5) <= VN453_data_out(2);
    CN174_sign_in(5) <= VN453_sign_out(2);
    CN174_data_in(6) <= VN514_data_out(2);
    CN174_sign_in(6) <= VN514_sign_out(2);
    CN174_data_in(7) <= VN597_data_out(2);
    CN174_sign_in(7) <= VN597_sign_out(2);
    CN174_data_in(8) <= VN753_data_out(2);
    CN174_sign_in(8) <= VN753_sign_out(2);
    CN174_data_in(9) <= VN984_data_out(2);
    CN174_sign_in(9) <= VN984_sign_out(2);
    CN174_data_in(10) <= VN1033_data_out(2);
    CN174_sign_in(10) <= VN1033_sign_out(2);
    CN174_data_in(11) <= VN1100_data_out(2);
    CN174_sign_in(11) <= VN1100_sign_out(2);
    CN174_data_in(12) <= VN1128_data_out(2);
    CN174_sign_in(12) <= VN1128_sign_out(2);
    CN174_data_in(13) <= VN1168_data_out(2);
    CN174_sign_in(13) <= VN1168_sign_out(2);
    CN174_data_in(14) <= VN1257_data_out(2);
    CN174_sign_in(14) <= VN1257_sign_out(2);
    CN174_data_in(15) <= VN1302_data_out(2);
    CN174_sign_in(15) <= VN1302_sign_out(2);
    CN174_data_in(16) <= VN1336_data_out(2);
    CN174_sign_in(16) <= VN1336_sign_out(2);
    CN174_data_in(17) <= VN1425_data_out(2);
    CN174_sign_in(17) <= VN1425_sign_out(2);
    CN174_data_in(18) <= VN1614_data_out(2);
    CN174_sign_in(18) <= VN1614_sign_out(2);
    CN174_data_in(19) <= VN1671_data_out(2);
    CN174_sign_in(19) <= VN1671_sign_out(2);
    CN174_data_in(20) <= VN1736_data_out(2);
    CN174_sign_in(20) <= VN1736_sign_out(2);
    CN174_data_in(21) <= VN1770_data_out(2);
    CN174_sign_in(21) <= VN1770_sign_out(2);
    CN174_data_in(22) <= VN1799_data_out(2);
    CN174_sign_in(22) <= VN1799_sign_out(2);
    CN174_data_in(23) <= VN1849_data_out(2);
    CN174_sign_in(23) <= VN1849_sign_out(2);
    CN174_data_in(24) <= VN1877_data_out(2);
    CN174_sign_in(24) <= VN1877_sign_out(2);
    CN174_data_in(25) <= VN1887_data_out(2);
    CN174_sign_in(25) <= VN1887_sign_out(2);
    CN174_data_in(26) <= VN1904_data_out(2);
    CN174_sign_in(26) <= VN1904_sign_out(2);
    CN174_data_in(27) <= VN1966_data_out(2);
    CN174_sign_in(27) <= VN1966_sign_out(2);
    CN174_data_in(28) <= VN1970_data_out(2);
    CN174_sign_in(28) <= VN1970_sign_out(2);
    CN174_data_in(29) <= VN1988_data_out(2);
    CN174_sign_in(29) <= VN1988_sign_out(2);
    CN174_data_in(30) <= VN1992_data_out(2);
    CN174_sign_in(30) <= VN1992_sign_out(2);
    CN174_data_in(31) <= VN1995_data_out(2);
    CN174_sign_in(31) <= VN1995_sign_out(2);
    CN175_data_in(0) <= VN8_data_out(2);
    CN175_sign_in(0) <= VN8_sign_out(2);
    CN175_data_in(1) <= VN82_data_out(2);
    CN175_sign_in(1) <= VN82_sign_out(2);
    CN175_data_in(2) <= VN117_data_out(2);
    CN175_sign_in(2) <= VN117_sign_out(2);
    CN175_data_in(3) <= VN211_data_out(2);
    CN175_sign_in(3) <= VN211_sign_out(2);
    CN175_data_in(4) <= VN278_data_out(2);
    CN175_sign_in(4) <= VN278_sign_out(2);
    CN175_data_in(5) <= VN325_data_out(2);
    CN175_sign_in(5) <= VN325_sign_out(2);
    CN175_data_in(6) <= VN344_data_out(2);
    CN175_sign_in(6) <= VN344_sign_out(2);
    CN175_data_in(7) <= VN445_data_out(2);
    CN175_sign_in(7) <= VN445_sign_out(2);
    CN175_data_in(8) <= VN503_data_out(2);
    CN175_sign_in(8) <= VN503_sign_out(2);
    CN175_data_in(9) <= VN535_data_out(2);
    CN175_sign_in(9) <= VN535_sign_out(2);
    CN175_data_in(10) <= VN590_data_out(2);
    CN175_sign_in(10) <= VN590_sign_out(2);
    CN175_data_in(11) <= VN638_data_out(2);
    CN175_sign_in(11) <= VN638_sign_out(2);
    CN175_data_in(12) <= VN709_data_out(2);
    CN175_sign_in(12) <= VN709_sign_out(2);
    CN175_data_in(13) <= VN735_data_out(2);
    CN175_sign_in(13) <= VN735_sign_out(2);
    CN175_data_in(14) <= VN815_data_out(2);
    CN175_sign_in(14) <= VN815_sign_out(2);
    CN175_data_in(15) <= VN846_data_out(2);
    CN175_sign_in(15) <= VN846_sign_out(2);
    CN175_data_in(16) <= VN908_data_out(2);
    CN175_sign_in(16) <= VN908_sign_out(2);
    CN175_data_in(17) <= VN976_data_out(2);
    CN175_sign_in(17) <= VN976_sign_out(2);
    CN175_data_in(18) <= VN1106_data_out(2);
    CN175_sign_in(18) <= VN1106_sign_out(2);
    CN175_data_in(19) <= VN1135_data_out(2);
    CN175_sign_in(19) <= VN1135_sign_out(2);
    CN175_data_in(20) <= VN1164_data_out(2);
    CN175_sign_in(20) <= VN1164_sign_out(2);
    CN175_data_in(21) <= VN1172_data_out(2);
    CN175_sign_in(21) <= VN1172_sign_out(2);
    CN175_data_in(22) <= VN1260_data_out(2);
    CN175_sign_in(22) <= VN1260_sign_out(2);
    CN175_data_in(23) <= VN1293_data_out(2);
    CN175_sign_in(23) <= VN1293_sign_out(2);
    CN175_data_in(24) <= VN1340_data_out(2);
    CN175_sign_in(24) <= VN1340_sign_out(2);
    CN175_data_in(25) <= VN1395_data_out(2);
    CN175_sign_in(25) <= VN1395_sign_out(2);
    CN175_data_in(26) <= VN1438_data_out(2);
    CN175_sign_in(26) <= VN1438_sign_out(2);
    CN175_data_in(27) <= VN1495_data_out(2);
    CN175_sign_in(27) <= VN1495_sign_out(2);
    CN175_data_in(28) <= VN1505_data_out(2);
    CN175_sign_in(28) <= VN1505_sign_out(2);
    CN175_data_in(29) <= VN1606_data_out(2);
    CN175_sign_in(29) <= VN1606_sign_out(2);
    CN175_data_in(30) <= VN1627_data_out(2);
    CN175_sign_in(30) <= VN1627_sign_out(2);
    CN175_data_in(31) <= VN1764_data_out(2);
    CN175_sign_in(31) <= VN1764_sign_out(2);
    CN176_data_in(0) <= VN7_data_out(2);
    CN176_sign_in(0) <= VN7_sign_out(2);
    CN176_data_in(1) <= VN89_data_out(2);
    CN176_sign_in(1) <= VN89_sign_out(2);
    CN176_data_in(2) <= VN137_data_out(2);
    CN176_sign_in(2) <= VN137_sign_out(2);
    CN176_data_in(3) <= VN176_data_out(2);
    CN176_sign_in(3) <= VN176_sign_out(2);
    CN176_data_in(4) <= VN251_data_out(2);
    CN176_sign_in(4) <= VN251_sign_out(2);
    CN176_data_in(5) <= VN286_data_out(2);
    CN176_sign_in(5) <= VN286_sign_out(2);
    CN176_data_in(6) <= VN356_data_out(2);
    CN176_sign_in(6) <= VN356_sign_out(2);
    CN176_data_in(7) <= VN404_data_out(2);
    CN176_sign_in(7) <= VN404_sign_out(2);
    CN176_data_in(8) <= VN450_data_out(2);
    CN176_sign_in(8) <= VN450_sign_out(2);
    CN176_data_in(9) <= VN533_data_out(2);
    CN176_sign_in(9) <= VN533_sign_out(2);
    CN176_data_in(10) <= VN566_data_out(2);
    CN176_sign_in(10) <= VN566_sign_out(2);
    CN176_data_in(11) <= VN664_data_out(2);
    CN176_sign_in(11) <= VN664_sign_out(2);
    CN176_data_in(12) <= VN686_data_out(2);
    CN176_sign_in(12) <= VN686_sign_out(2);
    CN176_data_in(13) <= VN746_data_out(2);
    CN176_sign_in(13) <= VN746_sign_out(2);
    CN176_data_in(14) <= VN817_data_out(2);
    CN176_sign_in(14) <= VN817_sign_out(2);
    CN176_data_in(15) <= VN867_data_out(2);
    CN176_sign_in(15) <= VN867_sign_out(2);
    CN176_data_in(16) <= VN910_data_out(2);
    CN176_sign_in(16) <= VN910_sign_out(2);
    CN176_data_in(17) <= VN993_data_out(2);
    CN176_sign_in(17) <= VN993_sign_out(2);
    CN176_data_in(18) <= VN1032_data_out(2);
    CN176_sign_in(18) <= VN1032_sign_out(2);
    CN176_data_in(19) <= VN1091_data_out(2);
    CN176_sign_in(19) <= VN1091_sign_out(2);
    CN176_data_in(20) <= VN1158_data_out(2);
    CN176_sign_in(20) <= VN1158_sign_out(2);
    CN176_data_in(21) <= VN1169_data_out(2);
    CN176_sign_in(21) <= VN1169_sign_out(2);
    CN176_data_in(22) <= VN1202_data_out(2);
    CN176_sign_in(22) <= VN1202_sign_out(2);
    CN176_data_in(23) <= VN1246_data_out(2);
    CN176_sign_in(23) <= VN1246_sign_out(2);
    CN176_data_in(24) <= VN1313_data_out(2);
    CN176_sign_in(24) <= VN1313_sign_out(2);
    CN176_data_in(25) <= VN1389_data_out(2);
    CN176_sign_in(25) <= VN1389_sign_out(2);
    CN176_data_in(26) <= VN1464_data_out(2);
    CN176_sign_in(26) <= VN1464_sign_out(2);
    CN176_data_in(27) <= VN1536_data_out(2);
    CN176_sign_in(27) <= VN1536_sign_out(2);
    CN176_data_in(28) <= VN1549_data_out(2);
    CN176_sign_in(28) <= VN1549_sign_out(2);
    CN176_data_in(29) <= VN1625_data_out(2);
    CN176_sign_in(29) <= VN1625_sign_out(2);
    CN176_data_in(30) <= VN1691_data_out(2);
    CN176_sign_in(30) <= VN1691_sign_out(2);
    CN176_data_in(31) <= VN1765_data_out(2);
    CN176_sign_in(31) <= VN1765_sign_out(2);
    CN177_data_in(0) <= VN6_data_out(2);
    CN177_sign_in(0) <= VN6_sign_out(2);
    CN177_data_in(1) <= VN109_data_out(2);
    CN177_sign_in(1) <= VN109_sign_out(2);
    CN177_data_in(2) <= VN147_data_out(2);
    CN177_sign_in(2) <= VN147_sign_out(2);
    CN177_data_in(3) <= VN204_data_out(2);
    CN177_sign_in(3) <= VN204_sign_out(2);
    CN177_data_in(4) <= VN232_data_out(2);
    CN177_sign_in(4) <= VN232_sign_out(2);
    CN177_data_in(5) <= VN304_data_out(2);
    CN177_sign_in(5) <= VN304_sign_out(2);
    CN177_data_in(6) <= VN368_data_out(2);
    CN177_sign_in(6) <= VN368_sign_out(2);
    CN177_data_in(7) <= VN397_data_out(2);
    CN177_sign_in(7) <= VN397_sign_out(2);
    CN177_data_in(8) <= VN496_data_out(2);
    CN177_sign_in(8) <= VN496_sign_out(2);
    CN177_data_in(9) <= VN512_data_out(2);
    CN177_sign_in(9) <= VN512_sign_out(2);
    CN177_data_in(10) <= VN576_data_out(2);
    CN177_sign_in(10) <= VN576_sign_out(2);
    CN177_data_in(11) <= VN651_data_out(2);
    CN177_sign_in(11) <= VN651_sign_out(2);
    CN177_data_in(12) <= VN721_data_out(2);
    CN177_sign_in(12) <= VN721_sign_out(2);
    CN177_data_in(13) <= VN754_data_out(2);
    CN177_sign_in(13) <= VN754_sign_out(2);
    CN177_data_in(14) <= VN787_data_out(2);
    CN177_sign_in(14) <= VN787_sign_out(2);
    CN177_data_in(15) <= VN881_data_out(2);
    CN177_sign_in(15) <= VN881_sign_out(2);
    CN177_data_in(16) <= VN895_data_out(2);
    CN177_sign_in(16) <= VN895_sign_out(2);
    CN177_data_in(17) <= VN998_data_out(2);
    CN177_sign_in(17) <= VN998_sign_out(2);
    CN177_data_in(18) <= VN1027_data_out(2);
    CN177_sign_in(18) <= VN1027_sign_out(2);
    CN177_data_in(19) <= VN1059_data_out(2);
    CN177_sign_in(19) <= VN1059_sign_out(2);
    CN177_data_in(20) <= VN1093_data_out(2);
    CN177_sign_in(20) <= VN1093_sign_out(2);
    CN177_data_in(21) <= VN1156_data_out(2);
    CN177_sign_in(21) <= VN1156_sign_out(2);
    CN177_data_in(22) <= VN1320_data_out(2);
    CN177_sign_in(22) <= VN1320_sign_out(2);
    CN177_data_in(23) <= VN1339_data_out(2);
    CN177_sign_in(23) <= VN1339_sign_out(2);
    CN177_data_in(24) <= VN1472_data_out(2);
    CN177_sign_in(24) <= VN1472_sign_out(2);
    CN177_data_in(25) <= VN1517_data_out(2);
    CN177_sign_in(25) <= VN1517_sign_out(2);
    CN177_data_in(26) <= VN1523_data_out(2);
    CN177_sign_in(26) <= VN1523_sign_out(2);
    CN177_data_in(27) <= VN1538_data_out(2);
    CN177_sign_in(27) <= VN1538_sign_out(2);
    CN177_data_in(28) <= VN1597_data_out(2);
    CN177_sign_in(28) <= VN1597_sign_out(2);
    CN177_data_in(29) <= VN1639_data_out(2);
    CN177_sign_in(29) <= VN1639_sign_out(2);
    CN177_data_in(30) <= VN1697_data_out(2);
    CN177_sign_in(30) <= VN1697_sign_out(2);
    CN177_data_in(31) <= VN1766_data_out(2);
    CN177_sign_in(31) <= VN1766_sign_out(2);
    CN178_data_in(0) <= VN5_data_out(2);
    CN178_sign_in(0) <= VN5_sign_out(2);
    CN178_data_in(1) <= VN107_data_out(2);
    CN178_sign_in(1) <= VN107_sign_out(2);
    CN178_data_in(2) <= VN142_data_out(2);
    CN178_sign_in(2) <= VN142_sign_out(2);
    CN178_data_in(3) <= VN201_data_out(2);
    CN178_sign_in(3) <= VN201_sign_out(2);
    CN178_data_in(4) <= VN313_data_out(2);
    CN178_sign_in(4) <= VN313_sign_out(2);
    CN178_data_in(5) <= VN338_data_out(2);
    CN178_sign_in(5) <= VN338_sign_out(2);
    CN178_data_in(6) <= VN428_data_out(2);
    CN178_sign_in(6) <= VN428_sign_out(2);
    CN178_data_in(7) <= VN549_data_out(2);
    CN178_sign_in(7) <= VN549_sign_out(2);
    CN178_data_in(8) <= VN621_data_out(2);
    CN178_sign_in(8) <= VN621_sign_out(2);
    CN178_data_in(9) <= VN728_data_out(2);
    CN178_sign_in(9) <= VN728_sign_out(2);
    CN178_data_in(10) <= VN823_data_out(2);
    CN178_sign_in(10) <= VN823_sign_out(2);
    CN178_data_in(11) <= VN877_data_out(2);
    CN178_sign_in(11) <= VN877_sign_out(2);
    CN178_data_in(12) <= VN927_data_out(2);
    CN178_sign_in(12) <= VN927_sign_out(2);
    CN178_data_in(13) <= VN1010_data_out(2);
    CN178_sign_in(13) <= VN1010_sign_out(2);
    CN178_data_in(14) <= VN1065_data_out(2);
    CN178_sign_in(14) <= VN1065_sign_out(2);
    CN178_data_in(15) <= VN1133_data_out(2);
    CN178_sign_in(15) <= VN1133_sign_out(2);
    CN178_data_in(16) <= VN1193_data_out(2);
    CN178_sign_in(16) <= VN1193_sign_out(2);
    CN178_data_in(17) <= VN1242_data_out(2);
    CN178_sign_in(17) <= VN1242_sign_out(2);
    CN178_data_in(18) <= VN1282_data_out(2);
    CN178_sign_in(18) <= VN1282_sign_out(2);
    CN178_data_in(19) <= VN1304_data_out(2);
    CN178_sign_in(19) <= VN1304_sign_out(2);
    CN178_data_in(20) <= VN1503_data_out(2);
    CN178_sign_in(20) <= VN1503_sign_out(2);
    CN178_data_in(21) <= VN1599_data_out(2);
    CN178_sign_in(21) <= VN1599_sign_out(2);
    CN178_data_in(22) <= VN1609_data_out(2);
    CN178_sign_in(22) <= VN1609_sign_out(2);
    CN178_data_in(23) <= VN1676_data_out(2);
    CN178_sign_in(23) <= VN1676_sign_out(2);
    CN178_data_in(24) <= VN1704_data_out(2);
    CN178_sign_in(24) <= VN1704_sign_out(2);
    CN178_data_in(25) <= VN1796_data_out(2);
    CN178_sign_in(25) <= VN1796_sign_out(2);
    CN178_data_in(26) <= VN1813_data_out(2);
    CN178_sign_in(26) <= VN1813_sign_out(2);
    CN178_data_in(27) <= VN1871_data_out(2);
    CN178_sign_in(27) <= VN1871_sign_out(2);
    CN178_data_in(28) <= VN1888_data_out(2);
    CN178_sign_in(28) <= VN1888_sign_out(2);
    CN178_data_in(29) <= VN1920_data_out(2);
    CN178_sign_in(29) <= VN1920_sign_out(2);
    CN178_data_in(30) <= VN1963_data_out(2);
    CN178_sign_in(30) <= VN1963_sign_out(2);
    CN178_data_in(31) <= VN1978_data_out(2);
    CN178_sign_in(31) <= VN1978_sign_out(2);
    CN179_data_in(0) <= VN4_data_out(2);
    CN179_sign_in(0) <= VN4_sign_out(2);
    CN179_data_in(1) <= VN87_data_out(2);
    CN179_sign_in(1) <= VN87_sign_out(2);
    CN179_data_in(2) <= VN148_data_out(2);
    CN179_sign_in(2) <= VN148_sign_out(2);
    CN179_data_in(3) <= VN215_data_out(2);
    CN179_sign_in(3) <= VN215_sign_out(2);
    CN179_data_in(4) <= VN267_data_out(2);
    CN179_sign_in(4) <= VN267_sign_out(2);
    CN179_data_in(5) <= VN308_data_out(2);
    CN179_sign_in(5) <= VN308_sign_out(2);
    CN179_data_in(6) <= VN386_data_out(2);
    CN179_sign_in(6) <= VN386_sign_out(2);
    CN179_data_in(7) <= VN438_data_out(2);
    CN179_sign_in(7) <= VN438_sign_out(2);
    CN179_data_in(8) <= VN460_data_out(2);
    CN179_sign_in(8) <= VN460_sign_out(2);
    CN179_data_in(9) <= VN552_data_out(2);
    CN179_sign_in(9) <= VN552_sign_out(2);
    CN179_data_in(10) <= VN573_data_out(2);
    CN179_sign_in(10) <= VN573_sign_out(2);
    CN179_data_in(11) <= VN666_data_out(2);
    CN179_sign_in(11) <= VN666_sign_out(2);
    CN179_data_in(12) <= VN711_data_out(2);
    CN179_sign_in(12) <= VN711_sign_out(2);
    CN179_data_in(13) <= VN742_data_out(2);
    CN179_sign_in(13) <= VN742_sign_out(2);
    CN179_data_in(14) <= VN780_data_out(2);
    CN179_sign_in(14) <= VN780_sign_out(2);
    CN179_data_in(15) <= VN841_data_out(2);
    CN179_sign_in(15) <= VN841_sign_out(2);
    CN179_data_in(16) <= VN891_data_out(2);
    CN179_sign_in(16) <= VN891_sign_out(2);
    CN179_data_in(17) <= VN997_data_out(2);
    CN179_sign_in(17) <= VN997_sign_out(2);
    CN179_data_in(18) <= VN1017_data_out(2);
    CN179_sign_in(18) <= VN1017_sign_out(2);
    CN179_data_in(19) <= VN1098_data_out(2);
    CN179_sign_in(19) <= VN1098_sign_out(2);
    CN179_data_in(20) <= VN1114_data_out(2);
    CN179_sign_in(20) <= VN1114_sign_out(2);
    CN179_data_in(21) <= VN1179_data_out(2);
    CN179_sign_in(21) <= VN1179_sign_out(2);
    CN179_data_in(22) <= VN1270_data_out(2);
    CN179_sign_in(22) <= VN1270_sign_out(2);
    CN179_data_in(23) <= VN1306_data_out(2);
    CN179_sign_in(23) <= VN1306_sign_out(2);
    CN179_data_in(24) <= VN1372_data_out(2);
    CN179_sign_in(24) <= VN1372_sign_out(2);
    CN179_data_in(25) <= VN1428_data_out(2);
    CN179_sign_in(25) <= VN1428_sign_out(2);
    CN179_data_in(26) <= VN1483_data_out(2);
    CN179_sign_in(26) <= VN1483_sign_out(2);
    CN179_data_in(27) <= VN1610_data_out(2);
    CN179_sign_in(27) <= VN1610_sign_out(2);
    CN179_data_in(28) <= VN1670_data_out(2);
    CN179_sign_in(28) <= VN1670_sign_out(2);
    CN179_data_in(29) <= VN1717_data_out(2);
    CN179_sign_in(29) <= VN1717_sign_out(2);
    CN179_data_in(30) <= VN1771_data_out(2);
    CN179_sign_in(30) <= VN1771_sign_out(2);
    CN179_data_in(31) <= VN1841_data_out(2);
    CN179_sign_in(31) <= VN1841_sign_out(2);
    CN180_data_in(0) <= VN67_data_out(2);
    CN180_sign_in(0) <= VN67_sign_out(2);
    CN180_data_in(1) <= VN208_data_out(2);
    CN180_sign_in(1) <= VN208_sign_out(2);
    CN180_data_in(2) <= VN263_data_out(2);
    CN180_sign_in(2) <= VN263_sign_out(2);
    CN180_data_in(3) <= VN314_data_out(2);
    CN180_sign_in(3) <= VN314_sign_out(2);
    CN180_data_in(4) <= VN371_data_out(2);
    CN180_sign_in(4) <= VN371_sign_out(2);
    CN180_data_in(5) <= VN432_data_out(2);
    CN180_sign_in(5) <= VN432_sign_out(2);
    CN180_data_in(6) <= VN472_data_out(2);
    CN180_sign_in(6) <= VN472_sign_out(2);
    CN180_data_in(7) <= VN536_data_out(2);
    CN180_sign_in(7) <= VN536_sign_out(2);
    CN180_data_in(8) <= VN563_data_out(2);
    CN180_sign_in(8) <= VN563_sign_out(2);
    CN180_data_in(9) <= VN687_data_out(2);
    CN180_sign_in(9) <= VN687_sign_out(2);
    CN180_data_in(10) <= VN770_data_out(2);
    CN180_sign_in(10) <= VN770_sign_out(2);
    CN180_data_in(11) <= VN788_data_out(2);
    CN180_sign_in(11) <= VN788_sign_out(2);
    CN180_data_in(12) <= VN863_data_out(2);
    CN180_sign_in(12) <= VN863_sign_out(2);
    CN180_data_in(13) <= VN919_data_out(2);
    CN180_sign_in(13) <= VN919_sign_out(2);
    CN180_data_in(14) <= VN1038_data_out(2);
    CN180_sign_in(14) <= VN1038_sign_out(2);
    CN180_data_in(15) <= VN1116_data_out(2);
    CN180_sign_in(15) <= VN1116_sign_out(2);
    CN180_data_in(16) <= VN1204_data_out(2);
    CN180_sign_in(16) <= VN1204_sign_out(2);
    CN180_data_in(17) <= VN1221_data_out(2);
    CN180_sign_in(17) <= VN1221_sign_out(2);
    CN180_data_in(18) <= VN1379_data_out(2);
    CN180_sign_in(18) <= VN1379_sign_out(2);
    CN180_data_in(19) <= VN1419_data_out(2);
    CN180_sign_in(19) <= VN1419_sign_out(2);
    CN180_data_in(20) <= VN1468_data_out(2);
    CN180_sign_in(20) <= VN1468_sign_out(2);
    CN180_data_in(21) <= VN1507_data_out(2);
    CN180_sign_in(21) <= VN1507_sign_out(2);
    CN180_data_in(22) <= VN1529_data_out(2);
    CN180_sign_in(22) <= VN1529_sign_out(2);
    CN180_data_in(23) <= VN1604_data_out(2);
    CN180_sign_in(23) <= VN1604_sign_out(2);
    CN180_data_in(24) <= VN1638_data_out(2);
    CN180_sign_in(24) <= VN1638_sign_out(2);
    CN180_data_in(25) <= VN1695_data_out(2);
    CN180_sign_in(25) <= VN1695_sign_out(2);
    CN180_data_in(26) <= VN1738_data_out(2);
    CN180_sign_in(26) <= VN1738_sign_out(2);
    CN180_data_in(27) <= VN1885_data_out(2);
    CN180_sign_in(27) <= VN1885_sign_out(2);
    CN180_data_in(28) <= VN1901_data_out(2);
    CN180_sign_in(28) <= VN1901_sign_out(2);
    CN180_data_in(29) <= VN1935_data_out(2);
    CN180_sign_in(29) <= VN1935_sign_out(2);
    CN180_data_in(30) <= VN2016_data_out(2);
    CN180_sign_in(30) <= VN2016_sign_out(2);
    CN180_data_in(31) <= VN2024_data_out(2);
    CN180_sign_in(31) <= VN2024_sign_out(2);
    CN181_data_in(0) <= VN3_data_out(2);
    CN181_sign_in(0) <= VN3_sign_out(2);
    CN181_data_in(1) <= VN70_data_out(2);
    CN181_sign_in(1) <= VN70_sign_out(2);
    CN181_data_in(2) <= VN162_data_out(2);
    CN181_sign_in(2) <= VN162_sign_out(2);
    CN181_data_in(3) <= VN186_data_out(2);
    CN181_sign_in(3) <= VN186_sign_out(2);
    CN181_data_in(4) <= VN227_data_out(2);
    CN181_sign_in(4) <= VN227_sign_out(2);
    CN181_data_in(5) <= VN303_data_out(2);
    CN181_sign_in(5) <= VN303_sign_out(2);
    CN181_data_in(6) <= VN389_data_out(2);
    CN181_sign_in(6) <= VN389_sign_out(2);
    CN181_data_in(7) <= VN436_data_out(2);
    CN181_sign_in(7) <= VN436_sign_out(2);
    CN181_data_in(8) <= VN482_data_out(2);
    CN181_sign_in(8) <= VN482_sign_out(2);
    CN181_data_in(9) <= VN513_data_out(2);
    CN181_sign_in(9) <= VN513_sign_out(2);
    CN181_data_in(10) <= VN598_data_out(2);
    CN181_sign_in(10) <= VN598_sign_out(2);
    CN181_data_in(11) <= VN619_data_out(2);
    CN181_sign_in(11) <= VN619_sign_out(2);
    CN181_data_in(12) <= VN708_data_out(2);
    CN181_sign_in(12) <= VN708_sign_out(2);
    CN181_data_in(13) <= VN816_data_out(2);
    CN181_sign_in(13) <= VN816_sign_out(2);
    CN181_data_in(14) <= VN864_data_out(2);
    CN181_sign_in(14) <= VN864_sign_out(2);
    CN181_data_in(15) <= VN904_data_out(2);
    CN181_sign_in(15) <= VN904_sign_out(2);
    CN181_data_in(16) <= VN973_data_out(2);
    CN181_sign_in(16) <= VN973_sign_out(2);
    CN181_data_in(17) <= VN1036_data_out(2);
    CN181_sign_in(17) <= VN1036_sign_out(2);
    CN181_data_in(18) <= VN1066_data_out(2);
    CN181_sign_in(18) <= VN1066_sign_out(2);
    CN181_data_in(19) <= VN1159_data_out(2);
    CN181_sign_in(19) <= VN1159_sign_out(2);
    CN181_data_in(20) <= VN1195_data_out(2);
    CN181_sign_in(20) <= VN1195_sign_out(2);
    CN181_data_in(21) <= VN1223_data_out(2);
    CN181_sign_in(21) <= VN1223_sign_out(2);
    CN181_data_in(22) <= VN1225_data_out(2);
    CN181_sign_in(22) <= VN1225_sign_out(2);
    CN181_data_in(23) <= VN1312_data_out(2);
    CN181_sign_in(23) <= VN1312_sign_out(2);
    CN181_data_in(24) <= VN1346_data_out(2);
    CN181_sign_in(24) <= VN1346_sign_out(2);
    CN181_data_in(25) <= VN1385_data_out(2);
    CN181_sign_in(25) <= VN1385_sign_out(2);
    CN181_data_in(26) <= VN1476_data_out(2);
    CN181_sign_in(26) <= VN1476_sign_out(2);
    CN181_data_in(27) <= VN1541_data_out(2);
    CN181_sign_in(27) <= VN1541_sign_out(2);
    CN181_data_in(28) <= VN1631_data_out(2);
    CN181_sign_in(28) <= VN1631_sign_out(2);
    CN181_data_in(29) <= VN1710_data_out(2);
    CN181_sign_in(29) <= VN1710_sign_out(2);
    CN181_data_in(30) <= VN1733_data_out(2);
    CN181_sign_in(30) <= VN1733_sign_out(2);
    CN181_data_in(31) <= VN1842_data_out(2);
    CN181_sign_in(31) <= VN1842_sign_out(2);
    CN182_data_in(0) <= VN2_data_out(2);
    CN182_sign_in(0) <= VN2_sign_out(2);
    CN182_data_in(1) <= VN54_data_out(2);
    CN182_sign_in(1) <= VN54_sign_out(2);
    CN182_data_in(2) <= VN169_data_out(2);
    CN182_sign_in(2) <= VN169_sign_out(2);
    CN182_data_in(3) <= VN195_data_out(2);
    CN182_sign_in(3) <= VN195_sign_out(2);
    CN182_data_in(4) <= VN248_data_out(2);
    CN182_sign_in(4) <= VN248_sign_out(2);
    CN182_data_in(5) <= VN328_data_out(2);
    CN182_sign_in(5) <= VN328_sign_out(2);
    CN182_data_in(6) <= VN350_data_out(2);
    CN182_sign_in(6) <= VN350_sign_out(2);
    CN182_data_in(7) <= VN425_data_out(2);
    CN182_sign_in(7) <= VN425_sign_out(2);
    CN182_data_in(8) <= VN454_data_out(2);
    CN182_sign_in(8) <= VN454_sign_out(2);
    CN182_data_in(9) <= VN532_data_out(2);
    CN182_sign_in(9) <= VN532_sign_out(2);
    CN182_data_in(10) <= VN582_data_out(2);
    CN182_sign_in(10) <= VN582_sign_out(2);
    CN182_data_in(11) <= VN647_data_out(2);
    CN182_sign_in(11) <= VN647_sign_out(2);
    CN182_data_in(12) <= VN678_data_out(2);
    CN182_sign_in(12) <= VN678_sign_out(2);
    CN182_data_in(13) <= VN772_data_out(2);
    CN182_sign_in(13) <= VN772_sign_out(2);
    CN182_data_in(14) <= VN829_data_out(2);
    CN182_sign_in(14) <= VN829_sign_out(2);
    CN182_data_in(15) <= VN840_data_out(2);
    CN182_sign_in(15) <= VN840_sign_out(2);
    CN182_data_in(16) <= VN929_data_out(2);
    CN182_sign_in(16) <= VN929_sign_out(2);
    CN182_data_in(17) <= VN1015_data_out(2);
    CN182_sign_in(17) <= VN1015_sign_out(2);
    CN182_data_in(18) <= VN1092_data_out(2);
    CN182_sign_in(18) <= VN1092_sign_out(2);
    CN182_data_in(19) <= VN1134_data_out(2);
    CN182_sign_in(19) <= VN1134_sign_out(2);
    CN182_data_in(20) <= VN1184_data_out(2);
    CN182_sign_in(20) <= VN1184_sign_out(2);
    CN182_data_in(21) <= VN1272_data_out(2);
    CN182_sign_in(21) <= VN1272_sign_out(2);
    CN182_data_in(22) <= VN1324_data_out(2);
    CN182_sign_in(22) <= VN1324_sign_out(2);
    CN182_data_in(23) <= VN1334_data_out(2);
    CN182_sign_in(23) <= VN1334_sign_out(2);
    CN182_data_in(24) <= VN1344_data_out(2);
    CN182_sign_in(24) <= VN1344_sign_out(2);
    CN182_data_in(25) <= VN1448_data_out(2);
    CN182_sign_in(25) <= VN1448_sign_out(2);
    CN182_data_in(26) <= VN1486_data_out(2);
    CN182_sign_in(26) <= VN1486_sign_out(2);
    CN182_data_in(27) <= VN1647_data_out(2);
    CN182_sign_in(27) <= VN1647_sign_out(2);
    CN182_data_in(28) <= VN1656_data_out(2);
    CN182_sign_in(28) <= VN1656_sign_out(2);
    CN182_data_in(29) <= VN1700_data_out(2);
    CN182_sign_in(29) <= VN1700_sign_out(2);
    CN182_data_in(30) <= VN1772_data_out(2);
    CN182_sign_in(30) <= VN1772_sign_out(2);
    CN182_data_in(31) <= VN1843_data_out(2);
    CN182_sign_in(31) <= VN1843_sign_out(2);
    CN183_data_in(0) <= VN1_data_out(2);
    CN183_sign_in(0) <= VN1_sign_out(2);
    CN183_data_in(1) <= VN88_data_out(2);
    CN183_sign_in(1) <= VN88_sign_out(2);
    CN183_data_in(2) <= VN190_data_out(2);
    CN183_sign_in(2) <= VN190_sign_out(2);
    CN183_data_in(3) <= VN281_data_out(2);
    CN183_sign_in(3) <= VN281_sign_out(2);
    CN183_data_in(4) <= VN358_data_out(2);
    CN183_sign_in(4) <= VN358_sign_out(2);
    CN183_data_in(5) <= VN405_data_out(2);
    CN183_sign_in(5) <= VN405_sign_out(2);
    CN183_data_in(6) <= VN498_data_out(2);
    CN183_sign_in(6) <= VN498_sign_out(2);
    CN183_data_in(7) <= VN560_data_out(2);
    CN183_sign_in(7) <= VN560_sign_out(2);
    CN183_data_in(8) <= VN593_data_out(2);
    CN183_sign_in(8) <= VN593_sign_out(2);
    CN183_data_in(9) <= VN644_data_out(2);
    CN183_sign_in(9) <= VN644_sign_out(2);
    CN183_data_in(10) <= VN718_data_out(2);
    CN183_sign_in(10) <= VN718_sign_out(2);
    CN183_data_in(11) <= VN730_data_out(2);
    CN183_sign_in(11) <= VN730_sign_out(2);
    CN183_data_in(12) <= VN802_data_out(2);
    CN183_sign_in(12) <= VN802_sign_out(2);
    CN183_data_in(13) <= VN832_data_out(2);
    CN183_sign_in(13) <= VN832_sign_out(2);
    CN183_data_in(14) <= VN921_data_out(2);
    CN183_sign_in(14) <= VN921_sign_out(2);
    CN183_data_in(15) <= VN944_data_out(2);
    CN183_sign_in(15) <= VN944_sign_out(2);
    CN183_data_in(16) <= VN1052_data_out(2);
    CN183_sign_in(16) <= VN1052_sign_out(2);
    CN183_data_in(17) <= VN1105_data_out(2);
    CN183_sign_in(17) <= VN1105_sign_out(2);
    CN183_data_in(18) <= VN1155_data_out(2);
    CN183_sign_in(18) <= VN1155_sign_out(2);
    CN183_data_in(19) <= VN1200_data_out(2);
    CN183_sign_in(19) <= VN1200_sign_out(2);
    CN183_data_in(20) <= VN1258_data_out(2);
    CN183_sign_in(20) <= VN1258_sign_out(2);
    CN183_data_in(21) <= VN1280_data_out(2);
    CN183_sign_in(21) <= VN1280_sign_out(2);
    CN183_data_in(22) <= VN1402_data_out(2);
    CN183_sign_in(22) <= VN1402_sign_out(2);
    CN183_data_in(23) <= VN1432_data_out(2);
    CN183_sign_in(23) <= VN1432_sign_out(2);
    CN183_data_in(24) <= VN1491_data_out(2);
    CN183_sign_in(24) <= VN1491_sign_out(2);
    CN183_data_in(25) <= VN1530_data_out(2);
    CN183_sign_in(25) <= VN1530_sign_out(2);
    CN183_data_in(26) <= VN1598_data_out(2);
    CN183_sign_in(26) <= VN1598_sign_out(2);
    CN183_data_in(27) <= VN1659_data_out(2);
    CN183_sign_in(27) <= VN1659_sign_out(2);
    CN183_data_in(28) <= VN1776_data_out(2);
    CN183_sign_in(28) <= VN1776_sign_out(2);
    CN183_data_in(29) <= VN1860_data_out(2);
    CN183_sign_in(29) <= VN1860_sign_out(2);
    CN183_data_in(30) <= VN1926_data_out(2);
    CN183_sign_in(30) <= VN1926_sign_out(2);
    CN183_data_in(31) <= VN1931_data_out(2);
    CN183_sign_in(31) <= VN1931_sign_out(2);
    CN184_data_in(0) <= VN0_data_out(2);
    CN184_sign_in(0) <= VN0_sign_out(2);
    CN184_data_in(1) <= VN106_data_out(2);
    CN184_sign_in(1) <= VN106_sign_out(2);
    CN184_data_in(2) <= VN153_data_out(2);
    CN184_sign_in(2) <= VN153_sign_out(2);
    CN184_data_in(3) <= VN193_data_out(2);
    CN184_sign_in(3) <= VN193_sign_out(2);
    CN184_data_in(4) <= VN226_data_out(2);
    CN184_sign_in(4) <= VN226_sign_out(2);
    CN184_data_in(5) <= VN318_data_out(2);
    CN184_sign_in(5) <= VN318_sign_out(2);
    CN184_data_in(6) <= VN354_data_out(2);
    CN184_sign_in(6) <= VN354_sign_out(2);
    CN184_data_in(7) <= VN444_data_out(2);
    CN184_sign_in(7) <= VN444_sign_out(2);
    CN184_data_in(8) <= VN484_data_out(2);
    CN184_sign_in(8) <= VN484_sign_out(2);
    CN184_data_in(9) <= VN545_data_out(2);
    CN184_sign_in(9) <= VN545_sign_out(2);
    CN184_data_in(10) <= VN603_data_out(2);
    CN184_sign_in(10) <= VN603_sign_out(2);
    CN184_data_in(11) <= VN658_data_out(2);
    CN184_sign_in(11) <= VN658_sign_out(2);
    CN184_data_in(12) <= VN689_data_out(2);
    CN184_sign_in(12) <= VN689_sign_out(2);
    CN184_data_in(13) <= VN726_data_out(2);
    CN184_sign_in(13) <= VN726_sign_out(2);
    CN184_data_in(14) <= VN783_data_out(2);
    CN184_sign_in(14) <= VN783_sign_out(2);
    CN184_data_in(15) <= VN850_data_out(2);
    CN184_sign_in(15) <= VN850_sign_out(2);
    CN184_data_in(16) <= VN909_data_out(2);
    CN184_sign_in(16) <= VN909_sign_out(2);
    CN184_data_in(17) <= VN1001_data_out(2);
    CN184_sign_in(17) <= VN1001_sign_out(2);
    CN184_data_in(18) <= VN1055_data_out(2);
    CN184_sign_in(18) <= VN1055_sign_out(2);
    CN184_data_in(19) <= VN1080_data_out(2);
    CN184_sign_in(19) <= VN1080_sign_out(2);
    CN184_data_in(20) <= VN1125_data_out(2);
    CN184_sign_in(20) <= VN1125_sign_out(2);
    CN184_data_in(21) <= VN1176_data_out(2);
    CN184_sign_in(21) <= VN1176_sign_out(2);
    CN184_data_in(22) <= VN1305_data_out(2);
    CN184_sign_in(22) <= VN1305_sign_out(2);
    CN184_data_in(23) <= VN1358_data_out(2);
    CN184_sign_in(23) <= VN1358_sign_out(2);
    CN184_data_in(24) <= VN1412_data_out(2);
    CN184_sign_in(24) <= VN1412_sign_out(2);
    CN184_data_in(25) <= VN1426_data_out(2);
    CN184_sign_in(25) <= VN1426_sign_out(2);
    CN184_data_in(26) <= VN1463_data_out(2);
    CN184_sign_in(26) <= VN1463_sign_out(2);
    CN184_data_in(27) <= VN1521_data_out(2);
    CN184_sign_in(27) <= VN1521_sign_out(2);
    CN184_data_in(28) <= VN1558_data_out(2);
    CN184_sign_in(28) <= VN1558_sign_out(2);
    CN184_data_in(29) <= VN1648_data_out(2);
    CN184_sign_in(29) <= VN1648_sign_out(2);
    CN184_data_in(30) <= VN1652_data_out(2);
    CN184_sign_in(30) <= VN1652_sign_out(2);
    CN184_data_in(31) <= VN1767_data_out(2);
    CN184_sign_in(31) <= VN1767_sign_out(2);
    CN185_data_in(0) <= VN121_data_out(2);
    CN185_sign_in(0) <= VN121_sign_out(2);
    CN185_data_in(1) <= VN272_data_out(2);
    CN185_sign_in(1) <= VN272_sign_out(2);
    CN185_data_in(2) <= VN320_data_out(2);
    CN185_sign_in(2) <= VN320_sign_out(2);
    CN185_data_in(3) <= VN359_data_out(2);
    CN185_sign_in(3) <= VN359_sign_out(2);
    CN185_data_in(4) <= VN501_data_out(2);
    CN185_sign_in(4) <= VN501_sign_out(2);
    CN185_data_in(5) <= VN577_data_out(2);
    CN185_sign_in(5) <= VN577_sign_out(2);
    CN185_data_in(6) <= VN680_data_out(2);
    CN185_sign_in(6) <= VN680_sign_out(2);
    CN185_data_in(7) <= VN804_data_out(2);
    CN185_sign_in(7) <= VN804_sign_out(2);
    CN185_data_in(8) <= VN926_data_out(2);
    CN185_sign_in(8) <= VN926_sign_out(2);
    CN185_data_in(9) <= VN979_data_out(2);
    CN185_sign_in(9) <= VN979_sign_out(2);
    CN185_data_in(10) <= VN1039_data_out(2);
    CN185_sign_in(10) <= VN1039_sign_out(2);
    CN185_data_in(11) <= VN1174_data_out(2);
    CN185_sign_in(11) <= VN1174_sign_out(2);
    CN185_data_in(12) <= VN1251_data_out(2);
    CN185_sign_in(12) <= VN1251_sign_out(2);
    CN185_data_in(13) <= VN1319_data_out(2);
    CN185_sign_in(13) <= VN1319_sign_out(2);
    CN185_data_in(14) <= VN1361_data_out(2);
    CN185_sign_in(14) <= VN1361_sign_out(2);
    CN185_data_in(15) <= VN1406_data_out(2);
    CN185_sign_in(15) <= VN1406_sign_out(2);
    CN185_data_in(16) <= VN1449_data_out(2);
    CN185_sign_in(16) <= VN1449_sign_out(2);
    CN185_data_in(17) <= VN1490_data_out(2);
    CN185_sign_in(17) <= VN1490_sign_out(2);
    CN185_data_in(18) <= VN1561_data_out(2);
    CN185_sign_in(18) <= VN1561_sign_out(2);
    CN185_data_in(19) <= VN1677_data_out(2);
    CN185_sign_in(19) <= VN1677_sign_out(2);
    CN185_data_in(20) <= VN1715_data_out(2);
    CN185_sign_in(20) <= VN1715_sign_out(2);
    CN185_data_in(21) <= VN1723_data_out(2);
    CN185_sign_in(21) <= VN1723_sign_out(2);
    CN185_data_in(22) <= VN1865_data_out(2);
    CN185_sign_in(22) <= VN1865_sign_out(2);
    CN185_data_in(23) <= VN1876_data_out(2);
    CN185_sign_in(23) <= VN1876_sign_out(2);
    CN185_data_in(24) <= VN1903_data_out(2);
    CN185_sign_in(24) <= VN1903_sign_out(2);
    CN185_data_in(25) <= VN1943_data_out(2);
    CN185_sign_in(25) <= VN1943_sign_out(2);
    CN185_data_in(26) <= VN1954_data_out(2);
    CN185_sign_in(26) <= VN1954_sign_out(2);
    CN185_data_in(27) <= VN1981_data_out(2);
    CN185_sign_in(27) <= VN1981_sign_out(2);
    CN185_data_in(28) <= VN2007_data_out(2);
    CN185_sign_in(28) <= VN2007_sign_out(2);
    CN185_data_in(29) <= VN2012_data_out(2);
    CN185_sign_in(29) <= VN2012_sign_out(2);
    CN185_data_in(30) <= VN2028_data_out(2);
    CN185_sign_in(30) <= VN2028_sign_out(2);
    CN185_data_in(31) <= VN2036_data_out(2);
    CN185_sign_in(31) <= VN2036_sign_out(2);
    CN186_data_in(0) <= VN63_data_out(2);
    CN186_sign_in(0) <= VN63_sign_out(2);
    CN186_data_in(1) <= VN160_data_out(2);
    CN186_sign_in(1) <= VN160_sign_out(2);
    CN186_data_in(2) <= VN216_data_out(2);
    CN186_sign_in(2) <= VN216_sign_out(2);
    CN186_data_in(3) <= VN235_data_out(2);
    CN186_sign_in(3) <= VN235_sign_out(2);
    CN186_data_in(4) <= VN290_data_out(2);
    CN186_sign_in(4) <= VN290_sign_out(2);
    CN186_data_in(5) <= VN349_data_out(2);
    CN186_sign_in(5) <= VN349_sign_out(2);
    CN186_data_in(6) <= VN410_data_out(2);
    CN186_sign_in(6) <= VN410_sign_out(2);
    CN186_data_in(7) <= VN465_data_out(2);
    CN186_sign_in(7) <= VN465_sign_out(2);
    CN186_data_in(8) <= VN507_data_out(2);
    CN186_sign_in(8) <= VN507_sign_out(2);
    CN186_data_in(9) <= VN565_data_out(2);
    CN186_sign_in(9) <= VN565_sign_out(2);
    CN186_data_in(10) <= VN627_data_out(2);
    CN186_sign_in(10) <= VN627_sign_out(2);
    CN186_data_in(11) <= VN669_data_out(2);
    CN186_sign_in(11) <= VN669_sign_out(2);
    CN186_data_in(12) <= VN766_data_out(2);
    CN186_sign_in(12) <= VN766_sign_out(2);
    CN186_data_in(13) <= VN818_data_out(2);
    CN186_sign_in(13) <= VN818_sign_out(2);
    CN186_data_in(14) <= VN900_data_out(2);
    CN186_sign_in(14) <= VN900_sign_out(2);
    CN186_data_in(15) <= VN958_data_out(2);
    CN186_sign_in(15) <= VN958_sign_out(2);
    CN186_data_in(16) <= VN1016_data_out(2);
    CN186_sign_in(16) <= VN1016_sign_out(2);
    CN186_data_in(17) <= VN1082_data_out(2);
    CN186_sign_in(17) <= VN1082_sign_out(2);
    CN186_data_in(18) <= VN1136_data_out(2);
    CN186_sign_in(18) <= VN1136_sign_out(2);
    CN186_data_in(19) <= VN1188_data_out(2);
    CN186_sign_in(19) <= VN1188_sign_out(2);
    CN186_data_in(20) <= VN1222_data_out(2);
    CN186_sign_in(20) <= VN1222_sign_out(2);
    CN186_data_in(21) <= VN1248_data_out(2);
    CN186_sign_in(21) <= VN1248_sign_out(2);
    CN186_data_in(22) <= VN1295_data_out(2);
    CN186_sign_in(22) <= VN1295_sign_out(2);
    CN186_data_in(23) <= VN1347_data_out(2);
    CN186_sign_in(23) <= VN1347_sign_out(2);
    CN186_data_in(24) <= VN1410_data_out(2);
    CN186_sign_in(24) <= VN1410_sign_out(2);
    CN186_data_in(25) <= VN1478_data_out(2);
    CN186_sign_in(25) <= VN1478_sign_out(2);
    CN186_data_in(26) <= VN1501_data_out(2);
    CN186_sign_in(26) <= VN1501_sign_out(2);
    CN186_data_in(27) <= VN1571_data_out(2);
    CN186_sign_in(27) <= VN1571_sign_out(2);
    CN186_data_in(28) <= VN1645_data_out(2);
    CN186_sign_in(28) <= VN1645_sign_out(2);
    CN186_data_in(29) <= VN1666_data_out(2);
    CN186_sign_in(29) <= VN1666_sign_out(2);
    CN186_data_in(30) <= VN1928_data_out(2);
    CN186_sign_in(30) <= VN1928_sign_out(2);
    CN186_data_in(31) <= VN1932_data_out(2);
    CN186_sign_in(31) <= VN1932_sign_out(2);
    CN187_data_in(0) <= VN90_data_out(2);
    CN187_sign_in(0) <= VN90_sign_out(2);
    CN187_data_in(1) <= VN113_data_out(2);
    CN187_sign_in(1) <= VN113_sign_out(2);
    CN187_data_in(2) <= VN200_data_out(2);
    CN187_sign_in(2) <= VN200_sign_out(2);
    CN187_data_in(3) <= VN240_data_out(2);
    CN187_sign_in(3) <= VN240_sign_out(2);
    CN187_data_in(4) <= VN326_data_out(2);
    CN187_sign_in(4) <= VN326_sign_out(2);
    CN187_data_in(5) <= VN374_data_out(2);
    CN187_sign_in(5) <= VN374_sign_out(2);
    CN187_data_in(6) <= VN439_data_out(2);
    CN187_sign_in(6) <= VN439_sign_out(2);
    CN187_data_in(7) <= VN474_data_out(2);
    CN187_sign_in(7) <= VN474_sign_out(2);
    CN187_data_in(8) <= VN550_data_out(2);
    CN187_sign_in(8) <= VN550_sign_out(2);
    CN187_data_in(9) <= VN606_data_out(2);
    CN187_sign_in(9) <= VN606_sign_out(2);
    CN187_data_in(10) <= VN636_data_out(2);
    CN187_sign_in(10) <= VN636_sign_out(2);
    CN187_data_in(11) <= VN685_data_out(2);
    CN187_sign_in(11) <= VN685_sign_out(2);
    CN187_data_in(12) <= VN767_data_out(2);
    CN187_sign_in(12) <= VN767_sign_out(2);
    CN187_data_in(13) <= VN814_data_out(2);
    CN187_sign_in(13) <= VN814_sign_out(2);
    CN187_data_in(14) <= VN854_data_out(2);
    CN187_sign_in(14) <= VN854_sign_out(2);
    CN187_data_in(15) <= VN897_data_out(2);
    CN187_sign_in(15) <= VN897_sign_out(2);
    CN187_data_in(16) <= VN961_data_out(2);
    CN187_sign_in(16) <= VN961_sign_out(2);
    CN187_data_in(17) <= VN1035_data_out(2);
    CN187_sign_in(17) <= VN1035_sign_out(2);
    CN187_data_in(18) <= VN1094_data_out(2);
    CN187_sign_in(18) <= VN1094_sign_out(2);
    CN187_data_in(19) <= VN1127_data_out(2);
    CN187_sign_in(19) <= VN1127_sign_out(2);
    CN187_data_in(20) <= VN1181_data_out(2);
    CN187_sign_in(20) <= VN1181_sign_out(2);
    CN187_data_in(21) <= VN1263_data_out(2);
    CN187_sign_in(21) <= VN1263_sign_out(2);
    CN187_data_in(22) <= VN1327_data_out(2);
    CN187_sign_in(22) <= VN1327_sign_out(2);
    CN187_data_in(23) <= VN1378_data_out(2);
    CN187_sign_in(23) <= VN1378_sign_out(2);
    CN187_data_in(24) <= VN1399_data_out(2);
    CN187_sign_in(24) <= VN1399_sign_out(2);
    CN187_data_in(25) <= VN1554_data_out(2);
    CN187_sign_in(25) <= VN1554_sign_out(2);
    CN187_data_in(26) <= VN1564_data_out(2);
    CN187_sign_in(26) <= VN1564_sign_out(2);
    CN187_data_in(27) <= VN1590_data_out(2);
    CN187_sign_in(27) <= VN1590_sign_out(2);
    CN187_data_in(28) <= VN1629_data_out(2);
    CN187_sign_in(28) <= VN1629_sign_out(2);
    CN187_data_in(29) <= VN1672_data_out(2);
    CN187_sign_in(29) <= VN1672_sign_out(2);
    CN187_data_in(30) <= VN1722_data_out(2);
    CN187_sign_in(30) <= VN1722_sign_out(2);
    CN187_data_in(31) <= VN1768_data_out(2);
    CN187_sign_in(31) <= VN1768_sign_out(2);
    CN188_data_in(0) <= VN81_data_out(2);
    CN188_sign_in(0) <= VN81_sign_out(2);
    CN188_data_in(1) <= VN212_data_out(2);
    CN188_sign_in(1) <= VN212_sign_out(2);
    CN188_data_in(2) <= VN279_data_out(2);
    CN188_sign_in(2) <= VN279_sign_out(2);
    CN188_data_in(3) <= VN284_data_out(2);
    CN188_sign_in(3) <= VN284_sign_out(2);
    CN188_data_in(4) <= VN381_data_out(2);
    CN188_sign_in(4) <= VN381_sign_out(2);
    CN188_data_in(5) <= VN427_data_out(2);
    CN188_sign_in(5) <= VN427_sign_out(2);
    CN188_data_in(6) <= VN469_data_out(2);
    CN188_sign_in(6) <= VN469_sign_out(2);
    CN188_data_in(7) <= VN511_data_out(2);
    CN188_sign_in(7) <= VN511_sign_out(2);
    CN188_data_in(8) <= VN568_data_out(2);
    CN188_sign_in(8) <= VN568_sign_out(2);
    CN188_data_in(9) <= VN715_data_out(2);
    CN188_sign_in(9) <= VN715_sign_out(2);
    CN188_data_in(10) <= VN744_data_out(2);
    CN188_sign_in(10) <= VN744_sign_out(2);
    CN188_data_in(11) <= VN779_data_out(2);
    CN188_sign_in(11) <= VN779_sign_out(2);
    CN188_data_in(12) <= VN848_data_out(2);
    CN188_sign_in(12) <= VN848_sign_out(2);
    CN188_data_in(13) <= VN913_data_out(2);
    CN188_sign_in(13) <= VN913_sign_out(2);
    CN188_data_in(14) <= VN945_data_out(2);
    CN188_sign_in(14) <= VN945_sign_out(2);
    CN188_data_in(15) <= VN1090_data_out(2);
    CN188_sign_in(15) <= VN1090_sign_out(2);
    CN188_data_in(16) <= VN1108_data_out(2);
    CN188_sign_in(16) <= VN1108_sign_out(2);
    CN188_data_in(17) <= VN1212_data_out(2);
    CN188_sign_in(17) <= VN1212_sign_out(2);
    CN188_data_in(18) <= VN1256_data_out(2);
    CN188_sign_in(18) <= VN1256_sign_out(2);
    CN188_data_in(19) <= VN1343_data_out(2);
    CN188_sign_in(19) <= VN1343_sign_out(2);
    CN188_data_in(20) <= VN1542_data_out(2);
    CN188_sign_in(20) <= VN1542_sign_out(2);
    CN188_data_in(21) <= VN1568_data_out(2);
    CN188_sign_in(21) <= VN1568_sign_out(2);
    CN188_data_in(22) <= VN1721_data_out(2);
    CN188_sign_in(22) <= VN1721_sign_out(2);
    CN188_data_in(23) <= VN1737_data_out(2);
    CN188_sign_in(23) <= VN1737_sign_out(2);
    CN188_data_in(24) <= VN1774_data_out(2);
    CN188_sign_in(24) <= VN1774_sign_out(2);
    CN188_data_in(25) <= VN1783_data_out(2);
    CN188_sign_in(25) <= VN1783_sign_out(2);
    CN188_data_in(26) <= VN1812_data_out(2);
    CN188_sign_in(26) <= VN1812_sign_out(2);
    CN188_data_in(27) <= VN1825_data_out(2);
    CN188_sign_in(27) <= VN1825_sign_out(2);
    CN188_data_in(28) <= VN1828_data_out(2);
    CN188_sign_in(28) <= VN1828_sign_out(2);
    CN188_data_in(29) <= VN1852_data_out(2);
    CN188_sign_in(29) <= VN1852_sign_out(2);
    CN188_data_in(30) <= VN1870_data_out(2);
    CN188_sign_in(30) <= VN1870_sign_out(2);
    CN188_data_in(31) <= VN1884_data_out(2);
    CN188_sign_in(31) <= VN1884_sign_out(2);
    CN189_data_in(0) <= VN68_data_out(2);
    CN189_sign_in(0) <= VN68_sign_out(2);
    CN189_data_in(1) <= VN152_data_out(2);
    CN189_sign_in(1) <= VN152_sign_out(2);
    CN189_data_in(2) <= VN223_data_out(2);
    CN189_sign_in(2) <= VN223_sign_out(2);
    CN189_data_in(3) <= VN239_data_out(2);
    CN189_sign_in(3) <= VN239_sign_out(2);
    CN189_data_in(4) <= VN291_data_out(2);
    CN189_sign_in(4) <= VN291_sign_out(2);
    CN189_data_in(5) <= VN363_data_out(2);
    CN189_sign_in(5) <= VN363_sign_out(2);
    CN189_data_in(6) <= VN413_data_out(2);
    CN189_sign_in(6) <= VN413_sign_out(2);
    CN189_data_in(7) <= VN475_data_out(2);
    CN189_sign_in(7) <= VN475_sign_out(2);
    CN189_data_in(8) <= VN541_data_out(2);
    CN189_sign_in(8) <= VN541_sign_out(2);
    CN189_data_in(9) <= VN587_data_out(2);
    CN189_sign_in(9) <= VN587_sign_out(2);
    CN189_data_in(10) <= VN633_data_out(2);
    CN189_sign_in(10) <= VN633_sign_out(2);
    CN189_data_in(11) <= VN713_data_out(2);
    CN189_sign_in(11) <= VN713_sign_out(2);
    CN189_data_in(12) <= VN736_data_out(2);
    CN189_sign_in(12) <= VN736_sign_out(2);
    CN189_data_in(13) <= VN799_data_out(2);
    CN189_sign_in(13) <= VN799_sign_out(2);
    CN189_data_in(14) <= VN885_data_out(2);
    CN189_sign_in(14) <= VN885_sign_out(2);
    CN189_data_in(15) <= VN906_data_out(2);
    CN189_sign_in(15) <= VN906_sign_out(2);
    CN189_data_in(16) <= VN980_data_out(2);
    CN189_sign_in(16) <= VN980_sign_out(2);
    CN189_data_in(17) <= VN1048_data_out(2);
    CN189_sign_in(17) <= VN1048_sign_out(2);
    CN189_data_in(18) <= VN1132_data_out(2);
    CN189_sign_in(18) <= VN1132_sign_out(2);
    CN189_data_in(19) <= VN1233_data_out(2);
    CN189_sign_in(19) <= VN1233_sign_out(2);
    CN189_data_in(20) <= VN1307_data_out(2);
    CN189_sign_in(20) <= VN1307_sign_out(2);
    CN189_data_in(21) <= VN1418_data_out(2);
    CN189_sign_in(21) <= VN1418_sign_out(2);
    CN189_data_in(22) <= VN1444_data_out(2);
    CN189_sign_in(22) <= VN1444_sign_out(2);
    CN189_data_in(23) <= VN1506_data_out(2);
    CN189_sign_in(23) <= VN1506_sign_out(2);
    CN189_data_in(24) <= VN1559_data_out(2);
    CN189_sign_in(24) <= VN1559_sign_out(2);
    CN189_data_in(25) <= VN1596_data_out(2);
    CN189_sign_in(25) <= VN1596_sign_out(2);
    CN189_data_in(26) <= VN1662_data_out(2);
    CN189_sign_in(26) <= VN1662_sign_out(2);
    CN189_data_in(27) <= VN1719_data_out(2);
    CN189_sign_in(27) <= VN1719_sign_out(2);
    CN189_data_in(28) <= VN1740_data_out(2);
    CN189_sign_in(28) <= VN1740_sign_out(2);
    CN189_data_in(29) <= VN1748_data_out(2);
    CN189_sign_in(29) <= VN1748_sign_out(2);
    CN189_data_in(30) <= VN1793_data_out(2);
    CN189_sign_in(30) <= VN1793_sign_out(2);
    CN189_data_in(31) <= VN1844_data_out(2);
    CN189_sign_in(31) <= VN1844_sign_out(2);
    CN190_data_in(0) <= VN168_data_out(2);
    CN190_sign_in(0) <= VN168_sign_out(2);
    CN190_data_in(1) <= VN196_data_out(2);
    CN190_sign_in(1) <= VN196_sign_out(2);
    CN190_data_in(2) <= VN234_data_out(2);
    CN190_sign_in(2) <= VN234_sign_out(2);
    CN190_data_in(3) <= VN319_data_out(2);
    CN190_sign_in(3) <= VN319_sign_out(2);
    CN190_data_in(4) <= VN365_data_out(2);
    CN190_sign_in(4) <= VN365_sign_out(2);
    CN190_data_in(5) <= VN430_data_out(2);
    CN190_sign_in(5) <= VN430_sign_out(2);
    CN190_data_in(6) <= VN464_data_out(2);
    CN190_sign_in(6) <= VN464_sign_out(2);
    CN190_data_in(7) <= VN538_data_out(2);
    CN190_sign_in(7) <= VN538_sign_out(2);
    CN190_data_in(8) <= VN595_data_out(2);
    CN190_sign_in(8) <= VN595_sign_out(2);
    CN190_data_in(9) <= VN673_data_out(2);
    CN190_sign_in(9) <= VN673_sign_out(2);
    CN190_data_in(10) <= VN752_data_out(2);
    CN190_sign_in(10) <= VN752_sign_out(2);
    CN190_data_in(11) <= VN836_data_out(2);
    CN190_sign_in(11) <= VN836_sign_out(2);
    CN190_data_in(12) <= VN935_data_out(2);
    CN190_sign_in(12) <= VN935_sign_out(2);
    CN190_data_in(13) <= VN1000_data_out(2);
    CN190_sign_in(13) <= VN1000_sign_out(2);
    CN190_data_in(14) <= VN1018_data_out(2);
    CN190_sign_in(14) <= VN1018_sign_out(2);
    CN190_data_in(15) <= VN1112_data_out(2);
    CN190_sign_in(15) <= VN1112_sign_out(2);
    CN190_data_in(16) <= VN1241_data_out(2);
    CN190_sign_in(16) <= VN1241_sign_out(2);
    CN190_data_in(17) <= VN1355_data_out(2);
    CN190_sign_in(17) <= VN1355_sign_out(2);
    CN190_data_in(18) <= VN1433_data_out(2);
    CN190_sign_in(18) <= VN1433_sign_out(2);
    CN190_data_in(19) <= VN1466_data_out(2);
    CN190_sign_in(19) <= VN1466_sign_out(2);
    CN190_data_in(20) <= VN1485_data_out(2);
    CN190_sign_in(20) <= VN1485_sign_out(2);
    CN190_data_in(21) <= VN1653_data_out(2);
    CN190_sign_in(21) <= VN1653_sign_out(2);
    CN190_data_in(22) <= VN1720_data_out(2);
    CN190_sign_in(22) <= VN1720_sign_out(2);
    CN190_data_in(23) <= VN1753_data_out(2);
    CN190_sign_in(23) <= VN1753_sign_out(2);
    CN190_data_in(24) <= VN1782_data_out(2);
    CN190_sign_in(24) <= VN1782_sign_out(2);
    CN190_data_in(25) <= VN1821_data_out(2);
    CN190_sign_in(25) <= VN1821_sign_out(2);
    CN190_data_in(26) <= VN1905_data_out(2);
    CN190_sign_in(26) <= VN1905_sign_out(2);
    CN190_data_in(27) <= VN1968_data_out(2);
    CN190_sign_in(27) <= VN1968_sign_out(2);
    CN190_data_in(28) <= VN2002_data_out(2);
    CN190_sign_in(28) <= VN2002_sign_out(2);
    CN190_data_in(29) <= VN2004_data_out(2);
    CN190_sign_in(29) <= VN2004_sign_out(2);
    CN190_data_in(30) <= VN2038_data_out(2);
    CN190_sign_in(30) <= VN2038_sign_out(2);
    CN190_data_in(31) <= VN2040_data_out(2);
    CN190_sign_in(31) <= VN2040_sign_out(2);
    CN191_data_in(0) <= VN52_data_out(2);
    CN191_sign_in(0) <= VN52_sign_out(2);
    CN191_data_in(1) <= VN59_data_out(2);
    CN191_sign_in(1) <= VN59_sign_out(2);
    CN191_data_in(2) <= VN138_data_out(2);
    CN191_sign_in(2) <= VN138_sign_out(2);
    CN191_data_in(3) <= VN185_data_out(2);
    CN191_sign_in(3) <= VN185_sign_out(2);
    CN191_data_in(4) <= VN270_data_out(2);
    CN191_sign_in(4) <= VN270_sign_out(2);
    CN191_data_in(5) <= VN280_data_out(2);
    CN191_sign_in(5) <= VN280_sign_out(2);
    CN191_data_in(6) <= VN393_data_out(2);
    CN191_sign_in(6) <= VN393_sign_out(2);
    CN191_data_in(7) <= VN486_data_out(2);
    CN191_sign_in(7) <= VN486_sign_out(2);
    CN191_data_in(8) <= VN554_data_out(2);
    CN191_sign_in(8) <= VN554_sign_out(2);
    CN191_data_in(9) <= VN591_data_out(2);
    CN191_sign_in(9) <= VN591_sign_out(2);
    CN191_data_in(10) <= VN659_data_out(2);
    CN191_sign_in(10) <= VN659_sign_out(2);
    CN191_data_in(11) <= VN719_data_out(2);
    CN191_sign_in(11) <= VN719_sign_out(2);
    CN191_data_in(12) <= VN757_data_out(2);
    CN191_sign_in(12) <= VN757_sign_out(2);
    CN191_data_in(13) <= VN778_data_out(2);
    CN191_sign_in(13) <= VN778_sign_out(2);
    CN191_data_in(14) <= VN859_data_out(2);
    CN191_sign_in(14) <= VN859_sign_out(2);
    CN191_data_in(15) <= VN889_data_out(2);
    CN191_sign_in(15) <= VN889_sign_out(2);
    CN191_data_in(16) <= VN970_data_out(2);
    CN191_sign_in(16) <= VN970_sign_out(2);
    CN191_data_in(17) <= VN1009_data_out(2);
    CN191_sign_in(17) <= VN1009_sign_out(2);
    CN191_data_in(18) <= VN1078_data_out(2);
    CN191_sign_in(18) <= VN1078_sign_out(2);
    CN191_data_in(19) <= VN1161_data_out(2);
    CN191_sign_in(19) <= VN1161_sign_out(2);
    CN191_data_in(20) <= VN1217_data_out(2);
    CN191_sign_in(20) <= VN1217_sign_out(2);
    CN191_data_in(21) <= VN1224_data_out(2);
    CN191_sign_in(21) <= VN1224_sign_out(2);
    CN191_data_in(22) <= VN1236_data_out(2);
    CN191_sign_in(22) <= VN1236_sign_out(2);
    CN191_data_in(23) <= VN1322_data_out(2);
    CN191_sign_in(23) <= VN1322_sign_out(2);
    CN191_data_in(24) <= VN1333_data_out(2);
    CN191_sign_in(24) <= VN1333_sign_out(2);
    CN191_data_in(25) <= VN1380_data_out(2);
    CN191_sign_in(25) <= VN1380_sign_out(2);
    CN191_data_in(26) <= VN1548_data_out(2);
    CN191_sign_in(26) <= VN1548_sign_out(2);
    CN191_data_in(27) <= VN1585_data_out(2);
    CN191_sign_in(27) <= VN1585_sign_out(2);
    CN191_data_in(28) <= VN1634_data_out(2);
    CN191_sign_in(28) <= VN1634_sign_out(2);
    CN191_data_in(29) <= VN1684_data_out(2);
    CN191_sign_in(29) <= VN1684_sign_out(2);
    CN191_data_in(30) <= VN1703_data_out(2);
    CN191_sign_in(30) <= VN1703_sign_out(2);
    CN191_data_in(31) <= VN1769_data_out(2);
    CN191_sign_in(31) <= VN1769_sign_out(2);
    CN192_data_in(0) <= VN53_data_out(3);
    CN192_sign_in(0) <= VN53_sign_out(3);
    CN192_data_in(1) <= VN107_data_out(3);
    CN192_sign_in(1) <= VN107_sign_out(3);
    CN192_data_in(2) <= VN128_data_out(3);
    CN192_sign_in(2) <= VN128_sign_out(3);
    CN192_data_in(3) <= VN197_data_out(3);
    CN192_sign_in(3) <= VN197_sign_out(3);
    CN192_data_in(4) <= VN243_data_out(3);
    CN192_sign_in(4) <= VN243_sign_out(3);
    CN192_data_in(5) <= VN297_data_out(3);
    CN192_sign_in(5) <= VN297_sign_out(3);
    CN192_data_in(6) <= VN340_data_out(3);
    CN192_sign_in(6) <= VN340_sign_out(3);
    CN192_data_in(7) <= VN440_data_out(3);
    CN192_sign_in(7) <= VN440_sign_out(3);
    CN192_data_in(8) <= VN456_data_out(3);
    CN192_sign_in(8) <= VN456_sign_out(3);
    CN192_data_in(9) <= VN533_data_out(3);
    CN192_sign_in(9) <= VN533_sign_out(3);
    CN192_data_in(10) <= VN578_data_out(3);
    CN192_sign_in(10) <= VN578_sign_out(3);
    CN192_data_in(11) <= VN639_data_out(3);
    CN192_sign_in(11) <= VN639_sign_out(3);
    CN192_data_in(12) <= VN709_data_out(3);
    CN192_sign_in(12) <= VN709_sign_out(3);
    CN192_data_in(13) <= VN761_data_out(3);
    CN192_sign_in(13) <= VN761_sign_out(3);
    CN192_data_in(14) <= VN794_data_out(3);
    CN192_sign_in(14) <= VN794_sign_out(3);
    CN192_data_in(15) <= VN857_data_out(3);
    CN192_sign_in(15) <= VN857_sign_out(3);
    CN192_data_in(16) <= VN892_data_out(3);
    CN192_sign_in(16) <= VN892_sign_out(3);
    CN192_data_in(17) <= VN1001_data_out(3);
    CN192_sign_in(17) <= VN1001_sign_out(3);
    CN192_data_in(18) <= VN1036_data_out(3);
    CN192_sign_in(18) <= VN1036_sign_out(3);
    CN192_data_in(19) <= VN1072_data_out(3);
    CN192_sign_in(19) <= VN1072_sign_out(3);
    CN192_data_in(20) <= VN1156_data_out(3);
    CN192_sign_in(20) <= VN1156_sign_out(3);
    CN192_data_in(21) <= VN1243_data_out(3);
    CN192_sign_in(21) <= VN1243_sign_out(3);
    CN192_data_in(22) <= VN1344_data_out(3);
    CN192_sign_in(22) <= VN1344_sign_out(3);
    CN192_data_in(23) <= VN1415_data_out(3);
    CN192_sign_in(23) <= VN1415_sign_out(3);
    CN192_data_in(24) <= VN1455_data_out(3);
    CN192_sign_in(24) <= VN1455_sign_out(3);
    CN192_data_in(25) <= VN1485_data_out(3);
    CN192_sign_in(25) <= VN1485_sign_out(3);
    CN192_data_in(26) <= VN1518_data_out(3);
    CN192_sign_in(26) <= VN1518_sign_out(3);
    CN192_data_in(27) <= VN1580_data_out(3);
    CN192_sign_in(27) <= VN1580_sign_out(3);
    CN192_data_in(28) <= VN1663_data_out(3);
    CN192_sign_in(28) <= VN1663_sign_out(3);
    CN192_data_in(29) <= VN1734_data_out(3);
    CN192_sign_in(29) <= VN1734_sign_out(3);
    CN192_data_in(30) <= VN1788_data_out(3);
    CN192_sign_in(30) <= VN1788_sign_out(3);
    CN192_data_in(31) <= VN1845_data_out(3);
    CN192_sign_in(31) <= VN1845_sign_out(3);
    CN193_data_in(0) <= VN51_data_out(3);
    CN193_sign_in(0) <= VN51_sign_out(3);
    CN193_data_in(1) <= VN58_data_out(3);
    CN193_sign_in(1) <= VN58_sign_out(3);
    CN193_data_in(2) <= VN137_data_out(3);
    CN193_sign_in(2) <= VN137_sign_out(3);
    CN193_data_in(3) <= VN269_data_out(3);
    CN193_sign_in(3) <= VN269_sign_out(3);
    CN193_data_in(4) <= VN333_data_out(3);
    CN193_sign_in(4) <= VN333_sign_out(3);
    CN193_data_in(5) <= VN485_data_out(3);
    CN193_sign_in(5) <= VN485_sign_out(3);
    CN193_data_in(6) <= VN590_data_out(3);
    CN193_sign_in(6) <= VN590_sign_out(3);
    CN193_data_in(7) <= VN658_data_out(3);
    CN193_sign_in(7) <= VN658_sign_out(3);
    CN193_data_in(8) <= VN756_data_out(3);
    CN193_sign_in(8) <= VN756_sign_out(3);
    CN193_data_in(9) <= VN858_data_out(3);
    CN193_sign_in(9) <= VN858_sign_out(3);
    CN193_data_in(10) <= VN888_data_out(3);
    CN193_sign_in(10) <= VN888_sign_out(3);
    CN193_data_in(11) <= VN969_data_out(3);
    CN193_sign_in(11) <= VN969_sign_out(3);
    CN193_data_in(12) <= VN1008_data_out(3);
    CN193_sign_in(12) <= VN1008_sign_out(3);
    CN193_data_in(13) <= VN1160_data_out(3);
    CN193_sign_in(13) <= VN1160_sign_out(3);
    CN193_data_in(14) <= VN1216_data_out(3);
    CN193_sign_in(14) <= VN1216_sign_out(3);
    CN193_data_in(15) <= VN1223_data_out(3);
    CN193_sign_in(15) <= VN1223_sign_out(3);
    CN193_data_in(16) <= VN1235_data_out(3);
    CN193_sign_in(16) <= VN1235_sign_out(3);
    CN193_data_in(17) <= VN1321_data_out(3);
    CN193_sign_in(17) <= VN1321_sign_out(3);
    CN193_data_in(18) <= VN1379_data_out(3);
    CN193_sign_in(18) <= VN1379_sign_out(3);
    CN193_data_in(19) <= VN1584_data_out(3);
    CN193_sign_in(19) <= VN1584_sign_out(3);
    CN193_data_in(20) <= VN1633_data_out(3);
    CN193_sign_in(20) <= VN1633_sign_out(3);
    CN193_data_in(21) <= VN1683_data_out(3);
    CN193_sign_in(21) <= VN1683_sign_out(3);
    CN193_data_in(22) <= VN1702_data_out(3);
    CN193_sign_in(22) <= VN1702_sign_out(3);
    CN193_data_in(23) <= VN1877_data_out(3);
    CN193_sign_in(23) <= VN1877_sign_out(3);
    CN193_data_in(24) <= VN1899_data_out(3);
    CN193_sign_in(24) <= VN1899_sign_out(3);
    CN193_data_in(25) <= VN1944_data_out(3);
    CN193_sign_in(25) <= VN1944_sign_out(3);
    CN193_data_in(26) <= VN1985_data_out(3);
    CN193_sign_in(26) <= VN1985_sign_out(3);
    CN193_data_in(27) <= VN2022_data_out(3);
    CN193_sign_in(27) <= VN2022_sign_out(3);
    CN193_data_in(28) <= VN2027_data_out(3);
    CN193_sign_in(28) <= VN2027_sign_out(3);
    CN193_data_in(29) <= VN2032_data_out(3);
    CN193_sign_in(29) <= VN2032_sign_out(3);
    CN193_data_in(30) <= VN2040_data_out(3);
    CN193_sign_in(30) <= VN2040_sign_out(3);
    CN193_data_in(31) <= VN2042_data_out(3);
    CN193_sign_in(31) <= VN2042_sign_out(3);
    CN194_data_in(0) <= VN50_data_out(3);
    CN194_sign_in(0) <= VN50_sign_out(3);
    CN194_data_in(1) <= VN55_data_out(3);
    CN194_sign_in(1) <= VN55_sign_out(3);
    CN194_data_in(2) <= VN115_data_out(3);
    CN194_sign_in(2) <= VN115_sign_out(3);
    CN194_data_in(3) <= VN171_data_out(3);
    CN194_sign_in(3) <= VN171_sign_out(3);
    CN194_data_in(4) <= VN275_data_out(3);
    CN194_sign_in(4) <= VN275_sign_out(3);
    CN194_data_in(5) <= VN304_data_out(3);
    CN194_sign_in(5) <= VN304_sign_out(3);
    CN194_data_in(6) <= VN371_data_out(3);
    CN194_sign_in(6) <= VN371_sign_out(3);
    CN194_data_in(7) <= VN401_data_out(3);
    CN194_sign_in(7) <= VN401_sign_out(3);
    CN194_data_in(8) <= VN492_data_out(3);
    CN194_sign_in(8) <= VN492_sign_out(3);
    CN194_data_in(9) <= VN546_data_out(3);
    CN194_sign_in(9) <= VN546_sign_out(3);
    CN194_data_in(10) <= VN595_data_out(3);
    CN194_sign_in(10) <= VN595_sign_out(3);
    CN194_data_in(11) <= VN642_data_out(3);
    CN194_sign_in(11) <= VN642_sign_out(3);
    CN194_data_in(12) <= VN695_data_out(3);
    CN194_sign_in(12) <= VN695_sign_out(3);
    CN194_data_in(13) <= VN823_data_out(3);
    CN194_sign_in(13) <= VN823_sign_out(3);
    CN194_data_in(14) <= VN938_data_out(3);
    CN194_sign_in(14) <= VN938_sign_out(3);
    CN194_data_in(15) <= VN953_data_out(3);
    CN194_sign_in(15) <= VN953_sign_out(3);
    CN194_data_in(16) <= VN1052_data_out(3);
    CN194_sign_in(16) <= VN1052_sign_out(3);
    CN194_data_in(17) <= VN1106_data_out(3);
    CN194_sign_in(17) <= VN1106_sign_out(3);
    CN194_data_in(18) <= VN1118_data_out(3);
    CN194_sign_in(18) <= VN1118_sign_out(3);
    CN194_data_in(19) <= VN1208_data_out(3);
    CN194_sign_in(19) <= VN1208_sign_out(3);
    CN194_data_in(20) <= VN1219_data_out(3);
    CN194_sign_in(20) <= VN1219_sign_out(3);
    CN194_data_in(21) <= VN1239_data_out(3);
    CN194_sign_in(21) <= VN1239_sign_out(3);
    CN194_data_in(22) <= VN1290_data_out(3);
    CN194_sign_in(22) <= VN1290_sign_out(3);
    CN194_data_in(23) <= VN1370_data_out(3);
    CN194_sign_in(23) <= VN1370_sign_out(3);
    CN194_data_in(24) <= VN1412_data_out(3);
    CN194_sign_in(24) <= VN1412_sign_out(3);
    CN194_data_in(25) <= VN1428_data_out(3);
    CN194_sign_in(25) <= VN1428_sign_out(3);
    CN194_data_in(26) <= VN1499_data_out(3);
    CN194_sign_in(26) <= VN1499_sign_out(3);
    CN194_data_in(27) <= VN1585_data_out(3);
    CN194_sign_in(27) <= VN1585_sign_out(3);
    CN194_data_in(28) <= VN1616_data_out(3);
    CN194_sign_in(28) <= VN1616_sign_out(3);
    CN194_data_in(29) <= VN1654_data_out(3);
    CN194_sign_in(29) <= VN1654_sign_out(3);
    CN194_data_in(30) <= VN1792_data_out(3);
    CN194_sign_in(30) <= VN1792_sign_out(3);
    CN194_data_in(31) <= VN1846_data_out(3);
    CN194_sign_in(31) <= VN1846_sign_out(3);
    CN195_data_in(0) <= VN72_data_out(3);
    CN195_sign_in(0) <= VN72_sign_out(3);
    CN195_data_in(1) <= VN139_data_out(3);
    CN195_sign_in(1) <= VN139_sign_out(3);
    CN195_data_in(2) <= VN187_data_out(3);
    CN195_sign_in(2) <= VN187_sign_out(3);
    CN195_data_in(3) <= VN244_data_out(3);
    CN195_sign_in(3) <= VN244_sign_out(3);
    CN195_data_in(4) <= VN384_data_out(3);
    CN195_sign_in(4) <= VN384_sign_out(3);
    CN195_data_in(5) <= VN397_data_out(3);
    CN195_sign_in(5) <= VN397_sign_out(3);
    CN195_data_in(6) <= VN519_data_out(3);
    CN195_sign_in(6) <= VN519_sign_out(3);
    CN195_data_in(7) <= VN585_data_out(3);
    CN195_sign_in(7) <= VN585_sign_out(3);
    CN195_data_in(8) <= VN705_data_out(3);
    CN195_sign_in(8) <= VN705_sign_out(3);
    CN195_data_in(9) <= VN755_data_out(3);
    CN195_sign_in(9) <= VN755_sign_out(3);
    CN195_data_in(10) <= VN785_data_out(3);
    CN195_sign_in(10) <= VN785_sign_out(3);
    CN195_data_in(11) <= VN834_data_out(3);
    CN195_sign_in(11) <= VN834_sign_out(3);
    CN195_data_in(12) <= VN942_data_out(3);
    CN195_sign_in(12) <= VN942_sign_out(3);
    CN195_data_in(13) <= VN1098_data_out(3);
    CN195_sign_in(13) <= VN1098_sign_out(3);
    CN195_data_in(14) <= VN1188_data_out(3);
    CN195_sign_in(14) <= VN1188_sign_out(3);
    CN195_data_in(15) <= VN1229_data_out(3);
    CN195_sign_in(15) <= VN1229_sign_out(3);
    CN195_data_in(16) <= VN1291_data_out(3);
    CN195_sign_in(16) <= VN1291_sign_out(3);
    CN195_data_in(17) <= VN1358_data_out(3);
    CN195_sign_in(17) <= VN1358_sign_out(3);
    CN195_data_in(18) <= VN1400_data_out(3);
    CN195_sign_in(18) <= VN1400_sign_out(3);
    CN195_data_in(19) <= VN1438_data_out(3);
    CN195_sign_in(19) <= VN1438_sign_out(3);
    CN195_data_in(20) <= VN1464_data_out(3);
    CN195_sign_in(20) <= VN1464_sign_out(3);
    CN195_data_in(21) <= VN1555_data_out(3);
    CN195_sign_in(21) <= VN1555_sign_out(3);
    CN195_data_in(22) <= VN1619_data_out(3);
    CN195_sign_in(22) <= VN1619_sign_out(3);
    CN195_data_in(23) <= VN1668_data_out(3);
    CN195_sign_in(23) <= VN1668_sign_out(3);
    CN195_data_in(24) <= VN1718_data_out(3);
    CN195_sign_in(24) <= VN1718_sign_out(3);
    CN195_data_in(25) <= VN1729_data_out(3);
    CN195_sign_in(25) <= VN1729_sign_out(3);
    CN195_data_in(26) <= VN1732_data_out(3);
    CN195_sign_in(26) <= VN1732_sign_out(3);
    CN195_data_in(27) <= VN1790_data_out(3);
    CN195_sign_in(27) <= VN1790_sign_out(3);
    CN195_data_in(28) <= VN1827_data_out(3);
    CN195_sign_in(28) <= VN1827_sign_out(3);
    CN195_data_in(29) <= VN1833_data_out(3);
    CN195_sign_in(29) <= VN1833_sign_out(3);
    CN195_data_in(30) <= VN1843_data_out(3);
    CN195_sign_in(30) <= VN1843_sign_out(3);
    CN195_data_in(31) <= VN1885_data_out(3);
    CN195_sign_in(31) <= VN1885_sign_out(3);
    CN196_data_in(0) <= VN49_data_out(3);
    CN196_sign_in(0) <= VN49_sign_out(3);
    CN196_data_in(1) <= VN64_data_out(3);
    CN196_sign_in(1) <= VN64_sign_out(3);
    CN196_data_in(2) <= VN153_data_out(3);
    CN196_sign_in(2) <= VN153_sign_out(3);
    CN196_data_in(3) <= VN205_data_out(3);
    CN196_sign_in(3) <= VN205_sign_out(3);
    CN196_data_in(4) <= VN242_data_out(3);
    CN196_sign_in(4) <= VN242_sign_out(3);
    CN196_data_in(5) <= VN306_data_out(3);
    CN196_sign_in(5) <= VN306_sign_out(3);
    CN196_data_in(6) <= VN402_data_out(3);
    CN196_sign_in(6) <= VN402_sign_out(3);
    CN196_data_in(7) <= VN478_data_out(3);
    CN196_sign_in(7) <= VN478_sign_out(3);
    CN196_data_in(8) <= VN529_data_out(3);
    CN196_sign_in(8) <= VN529_sign_out(3);
    CN196_data_in(9) <= VN664_data_out(3);
    CN196_sign_in(9) <= VN664_sign_out(3);
    CN196_data_in(10) <= VN699_data_out(3);
    CN196_sign_in(10) <= VN699_sign_out(3);
    CN196_data_in(11) <= VN749_data_out(3);
    CN196_sign_in(11) <= VN749_sign_out(3);
    CN196_data_in(12) <= VN790_data_out(3);
    CN196_sign_in(12) <= VN790_sign_out(3);
    CN196_data_in(13) <= VN830_data_out(3);
    CN196_sign_in(13) <= VN830_sign_out(3);
    CN196_data_in(14) <= VN869_data_out(3);
    CN196_sign_in(14) <= VN869_sign_out(3);
    CN196_data_in(15) <= VN931_data_out(3);
    CN196_sign_in(15) <= VN931_sign_out(3);
    CN196_data_in(16) <= VN971_data_out(3);
    CN196_sign_in(16) <= VN971_sign_out(3);
    CN196_data_in(17) <= VN1043_data_out(3);
    CN196_sign_in(17) <= VN1043_sign_out(3);
    CN196_data_in(18) <= VN1063_data_out(3);
    CN196_sign_in(18) <= VN1063_sign_out(3);
    CN196_data_in(19) <= VN1142_data_out(3);
    CN196_sign_in(19) <= VN1142_sign_out(3);
    CN196_data_in(20) <= VN1172_data_out(3);
    CN196_sign_in(20) <= VN1172_sign_out(3);
    CN196_data_in(21) <= VN1263_data_out(3);
    CN196_sign_in(21) <= VN1263_sign_out(3);
    CN196_data_in(22) <= VN1320_data_out(3);
    CN196_sign_in(22) <= VN1320_sign_out(3);
    CN196_data_in(23) <= VN1376_data_out(3);
    CN196_sign_in(23) <= VN1376_sign_out(3);
    CN196_data_in(24) <= VN1550_data_out(3);
    CN196_sign_in(24) <= VN1550_sign_out(3);
    CN196_data_in(25) <= VN1571_data_out(3);
    CN196_sign_in(25) <= VN1571_sign_out(3);
    CN196_data_in(26) <= VN1604_data_out(3);
    CN196_sign_in(26) <= VN1604_sign_out(3);
    CN196_data_in(27) <= VN1673_data_out(3);
    CN196_sign_in(27) <= VN1673_sign_out(3);
    CN196_data_in(28) <= VN1728_data_out(3);
    CN196_sign_in(28) <= VN1728_sign_out(3);
    CN196_data_in(29) <= VN1740_data_out(3);
    CN196_sign_in(29) <= VN1740_sign_out(3);
    CN196_data_in(30) <= VN1769_data_out(3);
    CN196_sign_in(30) <= VN1769_sign_out(3);
    CN196_data_in(31) <= VN1847_data_out(3);
    CN196_sign_in(31) <= VN1847_sign_out(3);
    CN197_data_in(0) <= VN48_data_out(3);
    CN197_sign_in(0) <= VN48_sign_out(3);
    CN197_data_in(1) <= VN96_data_out(3);
    CN197_sign_in(1) <= VN96_sign_out(3);
    CN197_data_in(2) <= VN150_data_out(3);
    CN197_sign_in(2) <= VN150_sign_out(3);
    CN197_data_in(3) <= VN213_data_out(3);
    CN197_sign_in(3) <= VN213_sign_out(3);
    CN197_data_in(4) <= VN273_data_out(3);
    CN197_sign_in(4) <= VN273_sign_out(3);
    CN197_data_in(5) <= VN320_data_out(3);
    CN197_sign_in(5) <= VN320_sign_out(3);
    CN197_data_in(6) <= VN363_data_out(3);
    CN197_sign_in(6) <= VN363_sign_out(3);
    CN197_data_in(7) <= VN504_data_out(3);
    CN197_sign_in(7) <= VN504_sign_out(3);
    CN197_data_in(8) <= VN523_data_out(3);
    CN197_sign_in(8) <= VN523_sign_out(3);
    CN197_data_in(9) <= VN614_data_out(3);
    CN197_sign_in(9) <= VN614_sign_out(3);
    CN197_data_in(10) <= VN636_data_out(3);
    CN197_sign_in(10) <= VN636_sign_out(3);
    CN197_data_in(11) <= VN703_data_out(3);
    CN197_sign_in(11) <= VN703_sign_out(3);
    CN197_data_in(12) <= VN732_data_out(3);
    CN197_sign_in(12) <= VN732_sign_out(3);
    CN197_data_in(13) <= VN872_data_out(3);
    CN197_sign_in(13) <= VN872_sign_out(3);
    CN197_data_in(14) <= VN887_data_out(3);
    CN197_sign_in(14) <= VN887_sign_out(3);
    CN197_data_in(15) <= VN913_data_out(3);
    CN197_sign_in(15) <= VN913_sign_out(3);
    CN197_data_in(16) <= VN958_data_out(3);
    CN197_sign_in(16) <= VN958_sign_out(3);
    CN197_data_in(17) <= VN1040_data_out(3);
    CN197_sign_in(17) <= VN1040_sign_out(3);
    CN197_data_in(18) <= VN1068_data_out(3);
    CN197_sign_in(18) <= VN1068_sign_out(3);
    CN197_data_in(19) <= VN1153_data_out(3);
    CN197_sign_in(19) <= VN1153_sign_out(3);
    CN197_data_in(20) <= VN1184_data_out(3);
    CN197_sign_in(20) <= VN1184_sign_out(3);
    CN197_data_in(21) <= VN1246_data_out(3);
    CN197_sign_in(21) <= VN1246_sign_out(3);
    CN197_data_in(22) <= VN1312_data_out(3);
    CN197_sign_in(22) <= VN1312_sign_out(3);
    CN197_data_in(23) <= VN1351_data_out(3);
    CN197_sign_in(23) <= VN1351_sign_out(3);
    CN197_data_in(24) <= VN1403_data_out(3);
    CN197_sign_in(24) <= VN1403_sign_out(3);
    CN197_data_in(25) <= VN1457_data_out(3);
    CN197_sign_in(25) <= VN1457_sign_out(3);
    CN197_data_in(26) <= VN1481_data_out(3);
    CN197_sign_in(26) <= VN1481_sign_out(3);
    CN197_data_in(27) <= VN1500_data_out(3);
    CN197_sign_in(27) <= VN1500_sign_out(3);
    CN197_data_in(28) <= VN1634_data_out(3);
    CN197_sign_in(28) <= VN1634_sign_out(3);
    CN197_data_in(29) <= VN1670_data_out(3);
    CN197_sign_in(29) <= VN1670_sign_out(3);
    CN197_data_in(30) <= VN1701_data_out(3);
    CN197_sign_in(30) <= VN1701_sign_out(3);
    CN197_data_in(31) <= VN1770_data_out(3);
    CN197_sign_in(31) <= VN1770_sign_out(3);
    CN198_data_in(0) <= VN47_data_out(3);
    CN198_sign_in(0) <= VN47_sign_out(3);
    CN198_data_in(1) <= VN105_data_out(3);
    CN198_sign_in(1) <= VN105_sign_out(3);
    CN198_data_in(2) <= VN111_data_out(3);
    CN198_sign_in(2) <= VN111_sign_out(3);
    CN198_data_in(3) <= VN208_data_out(3);
    CN198_sign_in(3) <= VN208_sign_out(3);
    CN198_data_in(4) <= VN254_data_out(3);
    CN198_sign_in(4) <= VN254_sign_out(3);
    CN198_data_in(5) <= VN316_data_out(3);
    CN198_sign_in(5) <= VN316_sign_out(3);
    CN198_data_in(6) <= VN379_data_out(3);
    CN198_sign_in(6) <= VN379_sign_out(3);
    CN198_data_in(7) <= VN415_data_out(3);
    CN198_sign_in(7) <= VN415_sign_out(3);
    CN198_data_in(8) <= VN484_data_out(3);
    CN198_sign_in(8) <= VN484_sign_out(3);
    CN198_data_in(9) <= VN526_data_out(3);
    CN198_sign_in(9) <= VN526_sign_out(3);
    CN198_data_in(10) <= VN599_data_out(3);
    CN198_sign_in(10) <= VN599_sign_out(3);
    CN198_data_in(11) <= VN625_data_out(3);
    CN198_sign_in(11) <= VN625_sign_out(3);
    CN198_data_in(12) <= VN692_data_out(3);
    CN198_sign_in(12) <= VN692_sign_out(3);
    CN198_data_in(13) <= VN739_data_out(3);
    CN198_sign_in(13) <= VN739_sign_out(3);
    CN198_data_in(14) <= VN789_data_out(3);
    CN198_sign_in(14) <= VN789_sign_out(3);
    CN198_data_in(15) <= VN859_data_out(3);
    CN198_sign_in(15) <= VN859_sign_out(3);
    CN198_data_in(16) <= VN895_data_out(3);
    CN198_sign_in(16) <= VN895_sign_out(3);
    CN198_data_in(17) <= VN977_data_out(3);
    CN198_sign_in(17) <= VN977_sign_out(3);
    CN198_data_in(18) <= VN1057_data_out(3);
    CN198_sign_in(18) <= VN1057_sign_out(3);
    CN198_data_in(19) <= VN1146_data_out(3);
    CN198_sign_in(19) <= VN1146_sign_out(3);
    CN198_data_in(20) <= VN1193_data_out(3);
    CN198_sign_in(20) <= VN1193_sign_out(3);
    CN198_data_in(21) <= VN1258_data_out(3);
    CN198_sign_in(21) <= VN1258_sign_out(3);
    CN198_data_in(22) <= VN1348_data_out(3);
    CN198_sign_in(22) <= VN1348_sign_out(3);
    CN198_data_in(23) <= VN1422_data_out(3);
    CN198_sign_in(23) <= VN1422_sign_out(3);
    CN198_data_in(24) <= VN1440_data_out(3);
    CN198_sign_in(24) <= VN1440_sign_out(3);
    CN198_data_in(25) <= VN1484_data_out(3);
    CN198_sign_in(25) <= VN1484_sign_out(3);
    CN198_data_in(26) <= VN1487_data_out(3);
    CN198_sign_in(26) <= VN1487_sign_out(3);
    CN198_data_in(27) <= VN1509_data_out(3);
    CN198_sign_in(27) <= VN1509_sign_out(3);
    CN198_data_in(28) <= VN1527_data_out(3);
    CN198_sign_in(28) <= VN1527_sign_out(3);
    CN198_data_in(29) <= VN1674_data_out(3);
    CN198_sign_in(29) <= VN1674_sign_out(3);
    CN198_data_in(30) <= VN1689_data_out(3);
    CN198_sign_in(30) <= VN1689_sign_out(3);
    CN198_data_in(31) <= VN1771_data_out(3);
    CN198_sign_in(31) <= VN1771_sign_out(3);
    CN199_data_in(0) <= VN46_data_out(3);
    CN199_sign_in(0) <= VN46_sign_out(3);
    CN199_data_in(1) <= VN99_data_out(3);
    CN199_sign_in(1) <= VN99_sign_out(3);
    CN199_data_in(2) <= VN133_data_out(3);
    CN199_sign_in(2) <= VN133_sign_out(3);
    CN199_data_in(3) <= VN214_data_out(3);
    CN199_sign_in(3) <= VN214_sign_out(3);
    CN199_data_in(4) <= VN257_data_out(3);
    CN199_sign_in(4) <= VN257_sign_out(3);
    CN199_data_in(5) <= VN282_data_out(3);
    CN199_sign_in(5) <= VN282_sign_out(3);
    CN199_data_in(6) <= VN350_data_out(3);
    CN199_sign_in(6) <= VN350_sign_out(3);
    CN199_data_in(7) <= VN422_data_out(3);
    CN199_sign_in(7) <= VN422_sign_out(3);
    CN199_data_in(8) <= VN496_data_out(3);
    CN199_sign_in(8) <= VN496_sign_out(3);
    CN199_data_in(9) <= VN517_data_out(3);
    CN199_sign_in(9) <= VN517_sign_out(3);
    CN199_data_in(10) <= VN601_data_out(3);
    CN199_sign_in(10) <= VN601_sign_out(3);
    CN199_data_in(11) <= VN667_data_out(3);
    CN199_sign_in(11) <= VN667_sign_out(3);
    CN199_data_in(12) <= VN673_data_out(3);
    CN199_sign_in(12) <= VN673_sign_out(3);
    CN199_data_in(13) <= VN762_data_out(3);
    CN199_sign_in(13) <= VN762_sign_out(3);
    CN199_data_in(14) <= VN784_data_out(3);
    CN199_sign_in(14) <= VN784_sign_out(3);
    CN199_data_in(15) <= VN835_data_out(3);
    CN199_sign_in(15) <= VN835_sign_out(3);
    CN199_data_in(16) <= VN909_data_out(3);
    CN199_sign_in(16) <= VN909_sign_out(3);
    CN199_data_in(17) <= VN949_data_out(3);
    CN199_sign_in(17) <= VN949_sign_out(3);
    CN199_data_in(18) <= VN1049_data_out(3);
    CN199_sign_in(18) <= VN1049_sign_out(3);
    CN199_data_in(19) <= VN1067_data_out(3);
    CN199_sign_in(19) <= VN1067_sign_out(3);
    CN199_data_in(20) <= VN1150_data_out(3);
    CN199_sign_in(20) <= VN1150_sign_out(3);
    CN199_data_in(21) <= VN1270_data_out(3);
    CN199_sign_in(21) <= VN1270_sign_out(3);
    CN199_data_in(22) <= VN1280_data_out(3);
    CN199_sign_in(22) <= VN1280_sign_out(3);
    CN199_data_in(23) <= VN1283_data_out(3);
    CN199_sign_in(23) <= VN1283_sign_out(3);
    CN199_data_in(24) <= VN1363_data_out(3);
    CN199_sign_in(24) <= VN1363_sign_out(3);
    CN199_data_in(25) <= VN1539_data_out(3);
    CN199_sign_in(25) <= VN1539_sign_out(3);
    CN199_data_in(26) <= VN1562_data_out(3);
    CN199_sign_in(26) <= VN1562_sign_out(3);
    CN199_data_in(27) <= VN1607_data_out(3);
    CN199_sign_in(27) <= VN1607_sign_out(3);
    CN199_data_in(28) <= VN1627_data_out(3);
    CN199_sign_in(28) <= VN1627_sign_out(3);
    CN199_data_in(29) <= VN1748_data_out(3);
    CN199_sign_in(29) <= VN1748_sign_out(3);
    CN199_data_in(30) <= VN1765_data_out(3);
    CN199_sign_in(30) <= VN1765_sign_out(3);
    CN199_data_in(31) <= VN1848_data_out(3);
    CN199_sign_in(31) <= VN1848_sign_out(3);
    CN200_data_in(0) <= VN45_data_out(3);
    CN200_sign_in(0) <= VN45_sign_out(3);
    CN200_data_in(1) <= VN102_data_out(3);
    CN200_sign_in(1) <= VN102_sign_out(3);
    CN200_data_in(2) <= VN134_data_out(3);
    CN200_sign_in(2) <= VN134_sign_out(3);
    CN200_data_in(3) <= VN204_data_out(3);
    CN200_sign_in(3) <= VN204_sign_out(3);
    CN200_data_in(4) <= VN245_data_out(3);
    CN200_sign_in(4) <= VN245_sign_out(3);
    CN200_data_in(5) <= VN300_data_out(3);
    CN200_sign_in(5) <= VN300_sign_out(3);
    CN200_data_in(6) <= VN387_data_out(3);
    CN200_sign_in(6) <= VN387_sign_out(3);
    CN200_data_in(7) <= VN406_data_out(3);
    CN200_sign_in(7) <= VN406_sign_out(3);
    CN200_data_in(8) <= VN448_data_out(3);
    CN200_sign_in(8) <= VN448_sign_out(3);
    CN200_data_in(9) <= VN554_data_out(3);
    CN200_sign_in(9) <= VN554_sign_out(3);
    CN200_data_in(10) <= VN570_data_out(3);
    CN200_sign_in(10) <= VN570_sign_out(3);
    CN200_data_in(11) <= VN628_data_out(3);
    CN200_sign_in(11) <= VN628_sign_out(3);
    CN200_data_in(12) <= VN711_data_out(3);
    CN200_sign_in(12) <= VN711_sign_out(3);
    CN200_data_in(13) <= VN760_data_out(3);
    CN200_sign_in(13) <= VN760_sign_out(3);
    CN200_data_in(14) <= VN820_data_out(3);
    CN200_sign_in(14) <= VN820_sign_out(3);
    CN200_data_in(15) <= VN856_data_out(3);
    CN200_sign_in(15) <= VN856_sign_out(3);
    CN200_data_in(16) <= VN919_data_out(3);
    CN200_sign_in(16) <= VN919_sign_out(3);
    CN200_data_in(17) <= VN946_data_out(3);
    CN200_sign_in(17) <= VN946_sign_out(3);
    CN200_data_in(18) <= VN1024_data_out(3);
    CN200_sign_in(18) <= VN1024_sign_out(3);
    CN200_data_in(19) <= VN1061_data_out(3);
    CN200_sign_in(19) <= VN1061_sign_out(3);
    CN200_data_in(20) <= VN1139_data_out(3);
    CN200_sign_in(20) <= VN1139_sign_out(3);
    CN200_data_in(21) <= VN1210_data_out(3);
    CN200_sign_in(21) <= VN1210_sign_out(3);
    CN200_data_in(22) <= VN1241_data_out(3);
    CN200_sign_in(22) <= VN1241_sign_out(3);
    CN200_data_in(23) <= VN1356_data_out(3);
    CN200_sign_in(23) <= VN1356_sign_out(3);
    CN200_data_in(24) <= VN1386_data_out(3);
    CN200_sign_in(24) <= VN1386_sign_out(3);
    CN200_data_in(25) <= VN1446_data_out(3);
    CN200_sign_in(25) <= VN1446_sign_out(3);
    CN200_data_in(26) <= VN1532_data_out(3);
    CN200_sign_in(26) <= VN1532_sign_out(3);
    CN200_data_in(27) <= VN1576_data_out(3);
    CN200_sign_in(27) <= VN1576_sign_out(3);
    CN200_data_in(28) <= VN1613_data_out(3);
    CN200_sign_in(28) <= VN1613_sign_out(3);
    CN200_data_in(29) <= VN1685_data_out(3);
    CN200_sign_in(29) <= VN1685_sign_out(3);
    CN200_data_in(30) <= VN1707_data_out(3);
    CN200_sign_in(30) <= VN1707_sign_out(3);
    CN200_data_in(31) <= VN1772_data_out(3);
    CN200_sign_in(31) <= VN1772_sign_out(3);
    CN201_data_in(0) <= VN44_data_out(3);
    CN201_sign_in(0) <= VN44_sign_out(3);
    CN201_data_in(1) <= VN93_data_out(3);
    CN201_sign_in(1) <= VN93_sign_out(3);
    CN201_data_in(2) <= VN169_data_out(3);
    CN201_sign_in(2) <= VN169_sign_out(3);
    CN201_data_in(3) <= VN174_data_out(3);
    CN201_sign_in(3) <= VN174_sign_out(3);
    CN201_data_in(4) <= VN274_data_out(3);
    CN201_sign_in(4) <= VN274_sign_out(3);
    CN201_data_in(5) <= VN351_data_out(3);
    CN201_sign_in(5) <= VN351_sign_out(3);
    CN201_data_in(6) <= VN407_data_out(3);
    CN201_sign_in(6) <= VN407_sign_out(3);
    CN201_data_in(7) <= VN477_data_out(3);
    CN201_sign_in(7) <= VN477_sign_out(3);
    CN201_data_in(8) <= VN536_data_out(3);
    CN201_sign_in(8) <= VN536_sign_out(3);
    CN201_data_in(9) <= VN606_data_out(3);
    CN201_sign_in(9) <= VN606_sign_out(3);
    CN201_data_in(10) <= VN648_data_out(3);
    CN201_sign_in(10) <= VN648_sign_out(3);
    CN201_data_in(11) <= VN669_data_out(3);
    CN201_sign_in(11) <= VN669_sign_out(3);
    CN201_data_in(12) <= VN737_data_out(3);
    CN201_sign_in(12) <= VN737_sign_out(3);
    CN201_data_in(13) <= VN881_data_out(3);
    CN201_sign_in(13) <= VN881_sign_out(3);
    CN201_data_in(14) <= VN889_data_out(3);
    CN201_sign_in(14) <= VN889_sign_out(3);
    CN201_data_in(15) <= VN963_data_out(3);
    CN201_sign_in(15) <= VN963_sign_out(3);
    CN201_data_in(16) <= VN1033_data_out(3);
    CN201_sign_in(16) <= VN1033_sign_out(3);
    CN201_data_in(17) <= VN1096_data_out(3);
    CN201_sign_in(17) <= VN1096_sign_out(3);
    CN201_data_in(18) <= VN1119_data_out(3);
    CN201_sign_in(18) <= VN1119_sign_out(3);
    CN201_data_in(19) <= VN1196_data_out(3);
    CN201_sign_in(19) <= VN1196_sign_out(3);
    CN201_data_in(20) <= VN1231_data_out(3);
    CN201_sign_in(20) <= VN1231_sign_out(3);
    CN201_data_in(21) <= VN1430_data_out(3);
    CN201_sign_in(21) <= VN1430_sign_out(3);
    CN201_data_in(22) <= VN1450_data_out(3);
    CN201_sign_in(22) <= VN1450_sign_out(3);
    CN201_data_in(23) <= VN1479_data_out(3);
    CN201_sign_in(23) <= VN1479_sign_out(3);
    CN201_data_in(24) <= VN1531_data_out(3);
    CN201_sign_in(24) <= VN1531_sign_out(3);
    CN201_data_in(25) <= VN1535_data_out(3);
    CN201_sign_in(25) <= VN1535_sign_out(3);
    CN201_data_in(26) <= VN1747_data_out(3);
    CN201_sign_in(26) <= VN1747_sign_out(3);
    CN201_data_in(27) <= VN1750_data_out(3);
    CN201_sign_in(27) <= VN1750_sign_out(3);
    CN201_data_in(28) <= VN1758_data_out(3);
    CN201_sign_in(28) <= VN1758_sign_out(3);
    CN201_data_in(29) <= VN1812_data_out(3);
    CN201_sign_in(29) <= VN1812_sign_out(3);
    CN201_data_in(30) <= VN1835_data_out(3);
    CN201_sign_in(30) <= VN1835_sign_out(3);
    CN201_data_in(31) <= VN1886_data_out(3);
    CN201_sign_in(31) <= VN1886_sign_out(3);
    CN202_data_in(0) <= VN43_data_out(3);
    CN202_sign_in(0) <= VN43_sign_out(3);
    CN202_data_in(1) <= VN73_data_out(3);
    CN202_sign_in(1) <= VN73_sign_out(3);
    CN202_data_in(2) <= VN160_data_out(3);
    CN202_sign_in(2) <= VN160_sign_out(3);
    CN202_data_in(3) <= VN181_data_out(3);
    CN202_sign_in(3) <= VN181_sign_out(3);
    CN202_data_in(4) <= VN281_data_out(3);
    CN202_sign_in(4) <= VN281_sign_out(3);
    CN202_data_in(5) <= VN365_data_out(3);
    CN202_sign_in(5) <= VN365_sign_out(3);
    CN202_data_in(6) <= VN433_data_out(3);
    CN202_sign_in(6) <= VN433_sign_out(3);
    CN202_data_in(7) <= VN491_data_out(3);
    CN202_sign_in(7) <= VN491_sign_out(3);
    CN202_data_in(8) <= VN550_data_out(3);
    CN202_sign_in(8) <= VN550_sign_out(3);
    CN202_data_in(9) <= VN563_data_out(3);
    CN202_sign_in(9) <= VN563_sign_out(3);
    CN202_data_in(10) <= VN655_data_out(3);
    CN202_sign_in(10) <= VN655_sign_out(3);
    CN202_data_in(11) <= VN678_data_out(3);
    CN202_sign_in(11) <= VN678_sign_out(3);
    CN202_data_in(12) <= VN773_data_out(3);
    CN202_sign_in(12) <= VN773_sign_out(3);
    CN202_data_in(13) <= VN795_data_out(3);
    CN202_sign_in(13) <= VN795_sign_out(3);
    CN202_data_in(14) <= VN933_data_out(3);
    CN202_sign_in(14) <= VN933_sign_out(3);
    CN202_data_in(15) <= VN955_data_out(3);
    CN202_sign_in(15) <= VN955_sign_out(3);
    CN202_data_in(16) <= VN1027_data_out(3);
    CN202_sign_in(16) <= VN1027_sign_out(3);
    CN202_data_in(17) <= VN1102_data_out(3);
    CN202_sign_in(17) <= VN1102_sign_out(3);
    CN202_data_in(18) <= VN1159_data_out(3);
    CN202_sign_in(18) <= VN1159_sign_out(3);
    CN202_data_in(19) <= VN1273_data_out(3);
    CN202_sign_in(19) <= VN1273_sign_out(3);
    CN202_data_in(20) <= VN1328_data_out(3);
    CN202_sign_in(20) <= VN1328_sign_out(3);
    CN202_data_in(21) <= VN1340_data_out(3);
    CN202_sign_in(21) <= VN1340_sign_out(3);
    CN202_data_in(22) <= VN1426_data_out(3);
    CN202_sign_in(22) <= VN1426_sign_out(3);
    CN202_data_in(23) <= VN1602_data_out(3);
    CN202_sign_in(23) <= VN1602_sign_out(3);
    CN202_data_in(24) <= VN1724_data_out(3);
    CN202_sign_in(24) <= VN1724_sign_out(3);
    CN202_data_in(25) <= VN1726_data_out(3);
    CN202_sign_in(25) <= VN1726_sign_out(3);
    CN202_data_in(26) <= VN1761_data_out(3);
    CN202_sign_in(26) <= VN1761_sign_out(3);
    CN202_data_in(27) <= VN1803_data_out(3);
    CN202_sign_in(27) <= VN1803_sign_out(3);
    CN202_data_in(28) <= VN1839_data_out(3);
    CN202_sign_in(28) <= VN1839_sign_out(3);
    CN202_data_in(29) <= VN1841_data_out(3);
    CN202_sign_in(29) <= VN1841_sign_out(3);
    CN202_data_in(30) <= VN1868_data_out(3);
    CN202_sign_in(30) <= VN1868_sign_out(3);
    CN202_data_in(31) <= VN1887_data_out(3);
    CN202_sign_in(31) <= VN1887_sign_out(3);
    CN203_data_in(0) <= VN42_data_out(3);
    CN203_sign_in(0) <= VN42_sign_out(3);
    CN203_data_in(1) <= VN54_data_out(3);
    CN203_sign_in(1) <= VN54_sign_out(3);
    CN203_data_in(2) <= VN119_data_out(3);
    CN203_sign_in(2) <= VN119_sign_out(3);
    CN203_data_in(3) <= VN217_data_out(3);
    CN203_sign_in(3) <= VN217_sign_out(3);
    CN203_data_in(4) <= VN267_data_out(3);
    CN203_sign_in(4) <= VN267_sign_out(3);
    CN203_data_in(5) <= VN326_data_out(3);
    CN203_sign_in(5) <= VN326_sign_out(3);
    CN203_data_in(6) <= VN361_data_out(3);
    CN203_sign_in(6) <= VN361_sign_out(3);
    CN203_data_in(7) <= VN413_data_out(3);
    CN203_sign_in(7) <= VN413_sign_out(3);
    CN203_data_in(8) <= VN465_data_out(3);
    CN203_sign_in(8) <= VN465_sign_out(3);
    CN203_data_in(9) <= VN560_data_out(3);
    CN203_sign_in(9) <= VN560_sign_out(3);
    CN203_data_in(10) <= VN571_data_out(3);
    CN203_sign_in(10) <= VN571_sign_out(3);
    CN203_data_in(11) <= VN706_data_out(3);
    CN203_sign_in(11) <= VN706_sign_out(3);
    CN203_data_in(12) <= VN793_data_out(3);
    CN203_sign_in(12) <= VN793_sign_out(3);
    CN203_data_in(13) <= VN836_data_out(3);
    CN203_sign_in(13) <= VN836_sign_out(3);
    CN203_data_in(14) <= VN988_data_out(3);
    CN203_sign_in(14) <= VN988_sign_out(3);
    CN203_data_in(15) <= VN1030_data_out(3);
    CN203_sign_in(15) <= VN1030_sign_out(3);
    CN203_data_in(16) <= VN1073_data_out(3);
    CN203_sign_in(16) <= VN1073_sign_out(3);
    CN203_data_in(17) <= VN1234_data_out(3);
    CN203_sign_in(17) <= VN1234_sign_out(3);
    CN203_data_in(18) <= VN1392_data_out(3);
    CN203_sign_in(18) <= VN1392_sign_out(3);
    CN203_data_in(19) <= VN1460_data_out(3);
    CN203_sign_in(19) <= VN1460_sign_out(3);
    CN203_data_in(20) <= VN1617_data_out(3);
    CN203_sign_in(20) <= VN1617_sign_out(3);
    CN203_data_in(21) <= VN1679_data_out(3);
    CN203_sign_in(21) <= VN1679_sign_out(3);
    CN203_data_in(22) <= VN1828_data_out(3);
    CN203_sign_in(22) <= VN1828_sign_out(3);
    CN203_data_in(23) <= VN1871_data_out(3);
    CN203_sign_in(23) <= VN1871_sign_out(3);
    CN203_data_in(24) <= VN1903_data_out(3);
    CN203_sign_in(24) <= VN1903_sign_out(3);
    CN203_data_in(25) <= VN1912_data_out(3);
    CN203_sign_in(25) <= VN1912_sign_out(3);
    CN203_data_in(26) <= VN1924_data_out(3);
    CN203_sign_in(26) <= VN1924_sign_out(3);
    CN203_data_in(27) <= VN1953_data_out(3);
    CN203_sign_in(27) <= VN1953_sign_out(3);
    CN203_data_in(28) <= VN1955_data_out(3);
    CN203_sign_in(28) <= VN1955_sign_out(3);
    CN203_data_in(29) <= VN1956_data_out(3);
    CN203_sign_in(29) <= VN1956_sign_out(3);
    CN203_data_in(30) <= VN2000_data_out(3);
    CN203_sign_in(30) <= VN2000_sign_out(3);
    CN203_data_in(31) <= VN2006_data_out(3);
    CN203_sign_in(31) <= VN2006_sign_out(3);
    CN204_data_in(0) <= VN41_data_out(3);
    CN204_sign_in(0) <= VN41_sign_out(3);
    CN204_data_in(1) <= VN68_data_out(3);
    CN204_sign_in(1) <= VN68_sign_out(3);
    CN204_data_in(2) <= VN123_data_out(3);
    CN204_sign_in(2) <= VN123_sign_out(3);
    CN204_data_in(3) <= VN219_data_out(3);
    CN204_sign_in(3) <= VN219_sign_out(3);
    CN204_data_in(4) <= VN251_data_out(3);
    CN204_sign_in(4) <= VN251_sign_out(3);
    CN204_data_in(5) <= VN288_data_out(3);
    CN204_sign_in(5) <= VN288_sign_out(3);
    CN204_data_in(6) <= VN382_data_out(3);
    CN204_sign_in(6) <= VN382_sign_out(3);
    CN204_data_in(7) <= VN425_data_out(3);
    CN204_sign_in(7) <= VN425_sign_out(3);
    CN204_data_in(8) <= VN499_data_out(3);
    CN204_sign_in(8) <= VN499_sign_out(3);
    CN204_data_in(9) <= VN530_data_out(3);
    CN204_sign_in(9) <= VN530_sign_out(3);
    CN204_data_in(10) <= VN600_data_out(3);
    CN204_sign_in(10) <= VN600_sign_out(3);
    CN204_data_in(11) <= VN656_data_out(3);
    CN204_sign_in(11) <= VN656_sign_out(3);
    CN204_data_in(12) <= VN694_data_out(3);
    CN204_sign_in(12) <= VN694_sign_out(3);
    CN204_data_in(13) <= VN763_data_out(3);
    CN204_sign_in(13) <= VN763_sign_out(3);
    CN204_data_in(14) <= VN826_data_out(3);
    CN204_sign_in(14) <= VN826_sign_out(3);
    CN204_data_in(15) <= VN883_data_out(3);
    CN204_sign_in(15) <= VN883_sign_out(3);
    CN204_data_in(16) <= VN936_data_out(3);
    CN204_sign_in(16) <= VN936_sign_out(3);
    CN204_data_in(17) <= VN998_data_out(3);
    CN204_sign_in(17) <= VN998_sign_out(3);
    CN204_data_in(18) <= VN1021_data_out(3);
    CN204_sign_in(18) <= VN1021_sign_out(3);
    CN204_data_in(19) <= VN1071_data_out(3);
    CN204_sign_in(19) <= VN1071_sign_out(3);
    CN204_data_in(20) <= VN1125_data_out(3);
    CN204_sign_in(20) <= VN1125_sign_out(3);
    CN204_data_in(21) <= VN1252_data_out(3);
    CN204_sign_in(21) <= VN1252_sign_out(3);
    CN204_data_in(22) <= VN1316_data_out(3);
    CN204_sign_in(22) <= VN1316_sign_out(3);
    CN204_data_in(23) <= VN1385_data_out(3);
    CN204_sign_in(23) <= VN1385_sign_out(3);
    CN204_data_in(24) <= VN1581_data_out(3);
    CN204_sign_in(24) <= VN1581_sign_out(3);
    CN204_data_in(25) <= VN1632_data_out(3);
    CN204_sign_in(25) <= VN1632_sign_out(3);
    CN204_data_in(26) <= VN1657_data_out(3);
    CN204_sign_in(26) <= VN1657_sign_out(3);
    CN204_data_in(27) <= VN1745_data_out(3);
    CN204_sign_in(27) <= VN1745_sign_out(3);
    CN204_data_in(28) <= VN1752_data_out(3);
    CN204_sign_in(28) <= VN1752_sign_out(3);
    CN204_data_in(29) <= VN1763_data_out(3);
    CN204_sign_in(29) <= VN1763_sign_out(3);
    CN204_data_in(30) <= VN1795_data_out(3);
    CN204_sign_in(30) <= VN1795_sign_out(3);
    CN204_data_in(31) <= VN1849_data_out(3);
    CN204_sign_in(31) <= VN1849_sign_out(3);
    CN205_data_in(0) <= VN170_data_out(3);
    CN205_sign_in(0) <= VN170_sign_out(3);
    CN205_data_in(1) <= VN276_data_out(3);
    CN205_sign_in(1) <= VN276_sign_out(3);
    CN205_data_in(2) <= VN345_data_out(3);
    CN205_sign_in(2) <= VN345_sign_out(3);
    CN205_data_in(3) <= VN434_data_out(3);
    CN205_sign_in(3) <= VN434_sign_out(3);
    CN205_data_in(4) <= VN613_data_out(3);
    CN205_sign_in(4) <= VN613_sign_out(3);
    CN205_data_in(5) <= VN647_data_out(3);
    CN205_sign_in(5) <= VN647_sign_out(3);
    CN205_data_in(6) <= VN738_data_out(3);
    CN205_sign_in(6) <= VN738_sign_out(3);
    CN205_data_in(7) <= VN870_data_out(3);
    CN205_sign_in(7) <= VN870_sign_out(3);
    CN205_data_in(8) <= VN901_data_out(3);
    CN205_sign_in(8) <= VN901_sign_out(3);
    CN205_data_in(9) <= VN1058_data_out(3);
    CN205_sign_in(9) <= VN1058_sign_out(3);
    CN205_data_in(10) <= VN1181_data_out(3);
    CN205_sign_in(10) <= VN1181_sign_out(3);
    CN205_data_in(11) <= VN1260_data_out(3);
    CN205_sign_in(11) <= VN1260_sign_out(3);
    CN205_data_in(12) <= VN1286_data_out(3);
    CN205_sign_in(12) <= VN1286_sign_out(3);
    CN205_data_in(13) <= VN1543_data_out(3);
    CN205_sign_in(13) <= VN1543_sign_out(3);
    CN205_data_in(14) <= VN1553_data_out(3);
    CN205_sign_in(14) <= VN1553_sign_out(3);
    CN205_data_in(15) <= VN1610_data_out(3);
    CN205_sign_in(15) <= VN1610_sign_out(3);
    CN205_data_in(16) <= VN1684_data_out(3);
    CN205_sign_in(16) <= VN1684_sign_out(3);
    CN205_data_in(17) <= VN1810_data_out(3);
    CN205_sign_in(17) <= VN1810_sign_out(3);
    CN205_data_in(18) <= VN1914_data_out(3);
    CN205_sign_in(18) <= VN1914_sign_out(3);
    CN205_data_in(19) <= VN1967_data_out(3);
    CN205_sign_in(19) <= VN1967_sign_out(3);
    CN205_data_in(20) <= VN1977_data_out(3);
    CN205_sign_in(20) <= VN1977_sign_out(3);
    CN205_data_in(21) <= VN1984_data_out(3);
    CN205_sign_in(21) <= VN1984_sign_out(3);
    CN205_data_in(22) <= VN1989_data_out(3);
    CN205_sign_in(22) <= VN1989_sign_out(3);
    CN205_data_in(23) <= VN1994_data_out(3);
    CN205_sign_in(23) <= VN1994_sign_out(3);
    CN205_data_in(24) <= VN1997_data_out(3);
    CN205_sign_in(24) <= VN1997_sign_out(3);
    CN205_data_in(25) <= VN2009_data_out(3);
    CN205_sign_in(25) <= VN2009_sign_out(3);
    CN205_data_in(26) <= VN2015_data_out(3);
    CN205_sign_in(26) <= VN2015_sign_out(3);
    CN205_data_in(27) <= VN2016_data_out(3);
    CN205_sign_in(27) <= VN2016_sign_out(3);
    CN205_data_in(28) <= VN2025_data_out(3);
    CN205_sign_in(28) <= VN2025_sign_out(3);
    CN205_data_in(29) <= VN2029_data_out(3);
    CN205_sign_in(29) <= VN2029_sign_out(3);
    CN205_data_in(30) <= VN2036_data_out(3);
    CN205_sign_in(30) <= VN2036_sign_out(3);
    CN205_data_in(31) <= VN2044_data_out(3);
    CN205_sign_in(31) <= VN2044_sign_out(3);
    CN206_data_in(0) <= VN40_data_out(3);
    CN206_sign_in(0) <= VN40_sign_out(3);
    CN206_data_in(1) <= VN122_data_out(3);
    CN206_sign_in(1) <= VN122_sign_out(3);
    CN206_data_in(2) <= VN172_data_out(3);
    CN206_sign_in(2) <= VN172_sign_out(3);
    CN206_data_in(3) <= VN332_data_out(3);
    CN206_sign_in(3) <= VN332_sign_out(3);
    CN206_data_in(4) <= VN346_data_out(3);
    CN206_sign_in(4) <= VN346_sign_out(3);
    CN206_data_in(5) <= VN479_data_out(3);
    CN206_sign_in(5) <= VN479_sign_out(3);
    CN206_data_in(6) <= VN587_data_out(3);
    CN206_sign_in(6) <= VN587_sign_out(3);
    CN206_data_in(7) <= VN617_data_out(3);
    CN206_sign_in(7) <= VN617_sign_out(3);
    CN206_data_in(8) <= VN697_data_out(3);
    CN206_sign_in(8) <= VN697_sign_out(3);
    CN206_data_in(9) <= VN759_data_out(3);
    CN206_sign_in(9) <= VN759_sign_out(3);
    CN206_data_in(10) <= VN808_data_out(3);
    CN206_sign_in(10) <= VN808_sign_out(3);
    CN206_data_in(11) <= VN833_data_out(3);
    CN206_sign_in(11) <= VN833_sign_out(3);
    CN206_data_in(12) <= VN910_data_out(3);
    CN206_sign_in(12) <= VN910_sign_out(3);
    CN206_data_in(13) <= VN995_data_out(3);
    CN206_sign_in(13) <= VN995_sign_out(3);
    CN206_data_in(14) <= VN1039_data_out(3);
    CN206_sign_in(14) <= VN1039_sign_out(3);
    CN206_data_in(15) <= VN1084_data_out(3);
    CN206_sign_in(15) <= VN1084_sign_out(3);
    CN206_data_in(16) <= VN1141_data_out(3);
    CN206_sign_in(16) <= VN1141_sign_out(3);
    CN206_data_in(17) <= VN1186_data_out(3);
    CN206_sign_in(17) <= VN1186_sign_out(3);
    CN206_data_in(18) <= VN1256_data_out(3);
    CN206_sign_in(18) <= VN1256_sign_out(3);
    CN206_data_in(19) <= VN1285_data_out(3);
    CN206_sign_in(19) <= VN1285_sign_out(3);
    CN206_data_in(20) <= VN1331_data_out(3);
    CN206_sign_in(20) <= VN1331_sign_out(3);
    CN206_data_in(21) <= VN1458_data_out(3);
    CN206_sign_in(21) <= VN1458_sign_out(3);
    CN206_data_in(22) <= VN1473_data_out(3);
    CN206_sign_in(22) <= VN1473_sign_out(3);
    CN206_data_in(23) <= VN1545_data_out(3);
    CN206_sign_in(23) <= VN1545_sign_out(3);
    CN206_data_in(24) <= VN1652_data_out(3);
    CN206_sign_in(24) <= VN1652_sign_out(3);
    CN206_data_in(25) <= VN1693_data_out(3);
    CN206_sign_in(25) <= VN1693_sign_out(3);
    CN206_data_in(26) <= VN1824_data_out(3);
    CN206_sign_in(26) <= VN1824_sign_out(3);
    CN206_data_in(27) <= VN1829_data_out(3);
    CN206_sign_in(27) <= VN1829_sign_out(3);
    CN206_data_in(28) <= VN1869_data_out(3);
    CN206_sign_in(28) <= VN1869_sign_out(3);
    CN206_data_in(29) <= VN1921_data_out(3);
    CN206_sign_in(29) <= VN1921_sign_out(3);
    CN206_data_in(30) <= VN1930_data_out(3);
    CN206_sign_in(30) <= VN1930_sign_out(3);
    CN206_data_in(31) <= VN1938_data_out(3);
    CN206_sign_in(31) <= VN1938_sign_out(3);
    CN207_data_in(0) <= VN39_data_out(3);
    CN207_sign_in(0) <= VN39_sign_out(3);
    CN207_data_in(1) <= VN95_data_out(3);
    CN207_sign_in(1) <= VN95_sign_out(3);
    CN207_data_in(2) <= VN117_data_out(3);
    CN207_sign_in(2) <= VN117_sign_out(3);
    CN207_data_in(3) <= VN255_data_out(3);
    CN207_sign_in(3) <= VN255_sign_out(3);
    CN207_data_in(4) <= VN292_data_out(3);
    CN207_sign_in(4) <= VN292_sign_out(3);
    CN207_data_in(5) <= VN381_data_out(3);
    CN207_sign_in(5) <= VN381_sign_out(3);
    CN207_data_in(6) <= VN391_data_out(3);
    CN207_sign_in(6) <= VN391_sign_out(3);
    CN207_data_in(7) <= VN421_data_out(3);
    CN207_sign_in(7) <= VN421_sign_out(3);
    CN207_data_in(8) <= VN521_data_out(3);
    CN207_sign_in(8) <= VN521_sign_out(3);
    CN207_data_in(9) <= VN566_data_out(3);
    CN207_sign_in(9) <= VN566_sign_out(3);
    CN207_data_in(10) <= VN622_data_out(3);
    CN207_sign_in(10) <= VN622_sign_out(3);
    CN207_data_in(11) <= VN716_data_out(3);
    CN207_sign_in(11) <= VN716_sign_out(3);
    CN207_data_in(12) <= VN730_data_out(3);
    CN207_sign_in(12) <= VN730_sign_out(3);
    CN207_data_in(13) <= VN796_data_out(3);
    CN207_sign_in(13) <= VN796_sign_out(3);
    CN207_data_in(14) <= VN864_data_out(3);
    CN207_sign_in(14) <= VN864_sign_out(3);
    CN207_data_in(15) <= VN906_data_out(3);
    CN207_sign_in(15) <= VN906_sign_out(3);
    CN207_data_in(16) <= VN985_data_out(3);
    CN207_sign_in(16) <= VN985_sign_out(3);
    CN207_data_in(17) <= VN1053_data_out(3);
    CN207_sign_in(17) <= VN1053_sign_out(3);
    CN207_data_in(18) <= VN1087_data_out(3);
    CN207_sign_in(18) <= VN1087_sign_out(3);
    CN207_data_in(19) <= VN1128_data_out(3);
    CN207_sign_in(19) <= VN1128_sign_out(3);
    CN207_data_in(20) <= VN1176_data_out(3);
    CN207_sign_in(20) <= VN1176_sign_out(3);
    CN207_data_in(21) <= VN1261_data_out(3);
    CN207_sign_in(21) <= VN1261_sign_out(3);
    CN207_data_in(22) <= VN1314_data_out(3);
    CN207_sign_in(22) <= VN1314_sign_out(3);
    CN207_data_in(23) <= VN1347_data_out(3);
    CN207_sign_in(23) <= VN1347_sign_out(3);
    CN207_data_in(24) <= VN1407_data_out(3);
    CN207_sign_in(24) <= VN1407_sign_out(3);
    CN207_data_in(25) <= VN1434_data_out(3);
    CN207_sign_in(25) <= VN1434_sign_out(3);
    CN207_data_in(26) <= VN1591_data_out(3);
    CN207_sign_in(26) <= VN1591_sign_out(3);
    CN207_data_in(27) <= VN1622_data_out(3);
    CN207_sign_in(27) <= VN1622_sign_out(3);
    CN207_data_in(28) <= VN1725_data_out(3);
    CN207_sign_in(28) <= VN1725_sign_out(3);
    CN207_data_in(29) <= VN1881_data_out(3);
    CN207_sign_in(29) <= VN1881_sign_out(3);
    CN207_data_in(30) <= VN1954_data_out(3);
    CN207_sign_in(30) <= VN1954_sign_out(3);
    CN207_data_in(31) <= VN1963_data_out(3);
    CN207_sign_in(31) <= VN1963_sign_out(3);
    CN208_data_in(0) <= VN38_data_out(3);
    CN208_sign_in(0) <= VN38_sign_out(3);
    CN208_data_in(1) <= VN82_data_out(3);
    CN208_sign_in(1) <= VN82_sign_out(3);
    CN208_data_in(2) <= VN157_data_out(3);
    CN208_sign_in(2) <= VN157_sign_out(3);
    CN208_data_in(3) <= VN191_data_out(3);
    CN208_sign_in(3) <= VN191_sign_out(3);
    CN208_data_in(4) <= VN286_data_out(3);
    CN208_sign_in(4) <= VN286_sign_out(3);
    CN208_data_in(5) <= VN372_data_out(3);
    CN208_sign_in(5) <= VN372_sign_out(3);
    CN208_data_in(6) <= VN393_data_out(3);
    CN208_sign_in(6) <= VN393_sign_out(3);
    CN208_data_in(7) <= VN494_data_out(3);
    CN208_sign_in(7) <= VN494_sign_out(3);
    CN208_data_in(8) <= VN542_data_out(3);
    CN208_sign_in(8) <= VN542_sign_out(3);
    CN208_data_in(9) <= VN588_data_out(3);
    CN208_sign_in(9) <= VN588_sign_out(3);
    CN208_data_in(10) <= VN660_data_out(3);
    CN208_sign_in(10) <= VN660_sign_out(3);
    CN208_data_in(11) <= VN770_data_out(3);
    CN208_sign_in(11) <= VN770_sign_out(3);
    CN208_data_in(12) <= VN861_data_out(3);
    CN208_sign_in(12) <= VN861_sign_out(3);
    CN208_data_in(13) <= VN911_data_out(3);
    CN208_sign_in(13) <= VN911_sign_out(3);
    CN208_data_in(14) <= VN1074_data_out(3);
    CN208_sign_in(14) <= VN1074_sign_out(3);
    CN208_data_in(15) <= VN1144_data_out(3);
    CN208_sign_in(15) <= VN1144_sign_out(3);
    CN208_data_in(16) <= VN1251_data_out(3);
    CN208_sign_in(16) <= VN1251_sign_out(3);
    CN208_data_in(17) <= VN1298_data_out(3);
    CN208_sign_in(17) <= VN1298_sign_out(3);
    CN208_data_in(18) <= VN1359_data_out(3);
    CN208_sign_in(18) <= VN1359_sign_out(3);
    CN208_data_in(19) <= VN1435_data_out(3);
    CN208_sign_in(19) <= VN1435_sign_out(3);
    CN208_data_in(20) <= VN1454_data_out(3);
    CN208_sign_in(20) <= VN1454_sign_out(3);
    CN208_data_in(21) <= VN1551_data_out(3);
    CN208_sign_in(21) <= VN1551_sign_out(3);
    CN208_data_in(22) <= VN1614_data_out(3);
    CN208_sign_in(22) <= VN1614_sign_out(3);
    CN208_data_in(23) <= VN1678_data_out(3);
    CN208_sign_in(23) <= VN1678_sign_out(3);
    CN208_data_in(24) <= VN1767_data_out(3);
    CN208_sign_in(24) <= VN1767_sign_out(3);
    CN208_data_in(25) <= VN1813_data_out(3);
    CN208_sign_in(25) <= VN1813_sign_out(3);
    CN208_data_in(26) <= VN1815_data_out(3);
    CN208_sign_in(26) <= VN1815_sign_out(3);
    CN208_data_in(27) <= VN1862_data_out(3);
    CN208_sign_in(27) <= VN1862_sign_out(3);
    CN208_data_in(28) <= VN1884_data_out(3);
    CN208_sign_in(28) <= VN1884_sign_out(3);
    CN208_data_in(29) <= VN1894_data_out(3);
    CN208_sign_in(29) <= VN1894_sign_out(3);
    CN208_data_in(30) <= VN1916_data_out(3);
    CN208_sign_in(30) <= VN1916_sign_out(3);
    CN208_data_in(31) <= VN1919_data_out(3);
    CN208_sign_in(31) <= VN1919_sign_out(3);
    CN209_data_in(0) <= VN37_data_out(3);
    CN209_sign_in(0) <= VN37_sign_out(3);
    CN209_data_in(1) <= VN97_data_out(3);
    CN209_sign_in(1) <= VN97_sign_out(3);
    CN209_data_in(2) <= VN165_data_out(3);
    CN209_sign_in(2) <= VN165_sign_out(3);
    CN209_data_in(3) <= VN218_data_out(3);
    CN209_sign_in(3) <= VN218_sign_out(3);
    CN209_data_in(4) <= VN323_data_out(3);
    CN209_sign_in(4) <= VN323_sign_out(3);
    CN209_data_in(5) <= VN428_data_out(3);
    CN209_sign_in(5) <= VN428_sign_out(3);
    CN209_data_in(6) <= VN461_data_out(3);
    CN209_sign_in(6) <= VN461_sign_out(3);
    CN209_data_in(7) <= VN552_data_out(3);
    CN209_sign_in(7) <= VN552_sign_out(3);
    CN209_data_in(8) <= VN662_data_out(3);
    CN209_sign_in(8) <= VN662_sign_out(3);
    CN209_data_in(9) <= VN719_data_out(3);
    CN209_sign_in(9) <= VN719_sign_out(3);
    CN209_data_in(10) <= VN740_data_out(3);
    CN209_sign_in(10) <= VN740_sign_out(3);
    CN209_data_in(11) <= VN792_data_out(3);
    CN209_sign_in(11) <= VN792_sign_out(3);
    CN209_data_in(12) <= VN875_data_out(3);
    CN209_sign_in(12) <= VN875_sign_out(3);
    CN209_data_in(13) <= VN900_data_out(3);
    CN209_sign_in(13) <= VN900_sign_out(3);
    CN209_data_in(14) <= VN945_data_out(3);
    CN209_sign_in(14) <= VN945_sign_out(3);
    CN209_data_in(15) <= VN1101_data_out(3);
    CN209_sign_in(15) <= VN1101_sign_out(3);
    CN209_data_in(16) <= VN1205_data_out(3);
    CN209_sign_in(16) <= VN1205_sign_out(3);
    CN209_data_in(17) <= VN1329_data_out(3);
    CN209_sign_in(17) <= VN1329_sign_out(3);
    CN209_data_in(18) <= VN1399_data_out(3);
    CN209_sign_in(18) <= VN1399_sign_out(3);
    CN209_data_in(19) <= VN1510_data_out(3);
    CN209_sign_in(19) <= VN1510_sign_out(3);
    CN209_data_in(20) <= VN1565_data_out(3);
    CN209_sign_in(20) <= VN1565_sign_out(3);
    CN209_data_in(21) <= VN1582_data_out(3);
    CN209_sign_in(21) <= VN1582_sign_out(3);
    CN209_data_in(22) <= VN1642_data_out(3);
    CN209_sign_in(22) <= VN1642_sign_out(3);
    CN209_data_in(23) <= VN1710_data_out(3);
    CN209_sign_in(23) <= VN1710_sign_out(3);
    CN209_data_in(24) <= VN1844_data_out(3);
    CN209_sign_in(24) <= VN1844_sign_out(3);
    CN209_data_in(25) <= VN1880_data_out(3);
    CN209_sign_in(25) <= VN1880_sign_out(3);
    CN209_data_in(26) <= VN1907_data_out(3);
    CN209_sign_in(26) <= VN1907_sign_out(3);
    CN209_data_in(27) <= VN1908_data_out(3);
    CN209_sign_in(27) <= VN1908_sign_out(3);
    CN209_data_in(28) <= VN1917_data_out(3);
    CN209_sign_in(28) <= VN1917_sign_out(3);
    CN209_data_in(29) <= VN1922_data_out(3);
    CN209_sign_in(29) <= VN1922_sign_out(3);
    CN209_data_in(30) <= VN1931_data_out(3);
    CN209_sign_in(30) <= VN1931_sign_out(3);
    CN209_data_in(31) <= VN1939_data_out(3);
    CN209_sign_in(31) <= VN1939_sign_out(3);
    CN210_data_in(0) <= VN36_data_out(3);
    CN210_sign_in(0) <= VN36_sign_out(3);
    CN210_data_in(1) <= VN60_data_out(3);
    CN210_sign_in(1) <= VN60_sign_out(3);
    CN210_data_in(2) <= VN129_data_out(3);
    CN210_sign_in(2) <= VN129_sign_out(3);
    CN210_data_in(3) <= VN180_data_out(3);
    CN210_sign_in(3) <= VN180_sign_out(3);
    CN210_data_in(4) <= VN246_data_out(3);
    CN210_sign_in(4) <= VN246_sign_out(3);
    CN210_data_in(5) <= VN330_data_out(3);
    CN210_sign_in(5) <= VN330_sign_out(3);
    CN210_data_in(6) <= VN335_data_out(3);
    CN210_sign_in(6) <= VN335_sign_out(3);
    CN210_data_in(7) <= VN395_data_out(3);
    CN210_sign_in(7) <= VN395_sign_out(3);
    CN210_data_in(8) <= VN462_data_out(3);
    CN210_sign_in(8) <= VN462_sign_out(3);
    CN210_data_in(9) <= VN547_data_out(3);
    CN210_sign_in(9) <= VN547_sign_out(3);
    CN210_data_in(10) <= VN598_data_out(3);
    CN210_sign_in(10) <= VN598_sign_out(3);
    CN210_data_in(11) <= VN630_data_out(3);
    CN210_sign_in(11) <= VN630_sign_out(3);
    CN210_data_in(12) <= VN671_data_out(3);
    CN210_sign_in(12) <= VN671_sign_out(3);
    CN210_data_in(13) <= VN731_data_out(3);
    CN210_sign_in(13) <= VN731_sign_out(3);
    CN210_data_in(14) <= VN818_data_out(3);
    CN210_sign_in(14) <= VN818_sign_out(3);
    CN210_data_in(15) <= VN867_data_out(3);
    CN210_sign_in(15) <= VN867_sign_out(3);
    CN210_data_in(16) <= VN924_data_out(3);
    CN210_sign_in(16) <= VN924_sign_out(3);
    CN210_data_in(17) <= VN959_data_out(3);
    CN210_sign_in(17) <= VN959_sign_out(3);
    CN210_data_in(18) <= VN1023_data_out(3);
    CN210_sign_in(18) <= VN1023_sign_out(3);
    CN210_data_in(19) <= VN1070_data_out(3);
    CN210_sign_in(19) <= VN1070_sign_out(3);
    CN210_data_in(20) <= VN1116_data_out(3);
    CN210_sign_in(20) <= VN1116_sign_out(3);
    CN210_data_in(21) <= VN1164_data_out(3);
    CN210_sign_in(21) <= VN1164_sign_out(3);
    CN210_data_in(22) <= VN1190_data_out(3);
    CN210_sign_in(22) <= VN1190_sign_out(3);
    CN210_data_in(23) <= VN1226_data_out(3);
    CN210_sign_in(23) <= VN1226_sign_out(3);
    CN210_data_in(24) <= VN1287_data_out(3);
    CN210_sign_in(24) <= VN1287_sign_out(3);
    CN210_data_in(25) <= VN1341_data_out(3);
    CN210_sign_in(25) <= VN1341_sign_out(3);
    CN210_data_in(26) <= VN1408_data_out(3);
    CN210_sign_in(26) <= VN1408_sign_out(3);
    CN210_data_in(27) <= VN1441_data_out(3);
    CN210_sign_in(27) <= VN1441_sign_out(3);
    CN210_data_in(28) <= VN1459_data_out(3);
    CN210_sign_in(28) <= VN1459_sign_out(3);
    CN210_data_in(29) <= VN1491_data_out(3);
    CN210_sign_in(29) <= VN1491_sign_out(3);
    CN210_data_in(30) <= VN1694_data_out(3);
    CN210_sign_in(30) <= VN1694_sign_out(3);
    CN210_data_in(31) <= VN1773_data_out(3);
    CN210_sign_in(31) <= VN1773_sign_out(3);
    CN211_data_in(0) <= VN35_data_out(3);
    CN211_sign_in(0) <= VN35_sign_out(3);
    CN211_data_in(1) <= VN70_data_out(3);
    CN211_sign_in(1) <= VN70_sign_out(3);
    CN211_data_in(2) <= VN127_data_out(3);
    CN211_sign_in(2) <= VN127_sign_out(3);
    CN211_data_in(3) <= VN206_data_out(3);
    CN211_sign_in(3) <= VN206_sign_out(3);
    CN211_data_in(4) <= VN260_data_out(3);
    CN211_sign_in(4) <= VN260_sign_out(3);
    CN211_data_in(5) <= VN298_data_out(3);
    CN211_sign_in(5) <= VN298_sign_out(3);
    CN211_data_in(6) <= VN408_data_out(3);
    CN211_sign_in(6) <= VN408_sign_out(3);
    CN211_data_in(7) <= VN493_data_out(3);
    CN211_sign_in(7) <= VN493_sign_out(3);
    CN211_data_in(8) <= VN553_data_out(3);
    CN211_sign_in(8) <= VN553_sign_out(3);
    CN211_data_in(9) <= VN561_data_out(3);
    CN211_sign_in(9) <= VN561_sign_out(3);
    CN211_data_in(10) <= VN715_data_out(3);
    CN211_sign_in(10) <= VN715_sign_out(3);
    CN211_data_in(11) <= VN774_data_out(3);
    CN211_sign_in(11) <= VN774_sign_out(3);
    CN211_data_in(12) <= VN802_data_out(3);
    CN211_sign_in(12) <= VN802_sign_out(3);
    CN211_data_in(13) <= VN844_data_out(3);
    CN211_sign_in(13) <= VN844_sign_out(3);
    CN211_data_in(14) <= VN930_data_out(3);
    CN211_sign_in(14) <= VN930_sign_out(3);
    CN211_data_in(15) <= VN970_data_out(3);
    CN211_sign_in(15) <= VN970_sign_out(3);
    CN211_data_in(16) <= VN1010_data_out(3);
    CN211_sign_in(16) <= VN1010_sign_out(3);
    CN211_data_in(17) <= VN1094_data_out(3);
    CN211_sign_in(17) <= VN1094_sign_out(3);
    CN211_data_in(18) <= VN1167_data_out(3);
    CN211_sign_in(18) <= VN1167_sign_out(3);
    CN211_data_in(19) <= VN1192_data_out(3);
    CN211_sign_in(19) <= VN1192_sign_out(3);
    CN211_data_in(20) <= VN1265_data_out(3);
    CN211_sign_in(20) <= VN1265_sign_out(3);
    CN211_data_in(21) <= VN1315_data_out(3);
    CN211_sign_in(21) <= VN1315_sign_out(3);
    CN211_data_in(22) <= VN1496_data_out(3);
    CN211_sign_in(22) <= VN1496_sign_out(3);
    CN211_data_in(23) <= VN1513_data_out(3);
    CN211_sign_in(23) <= VN1513_sign_out(3);
    CN211_data_in(24) <= VN1534_data_out(3);
    CN211_sign_in(24) <= VN1534_sign_out(3);
    CN211_data_in(25) <= VN1544_data_out(3);
    CN211_sign_in(25) <= VN1544_sign_out(3);
    CN211_data_in(26) <= VN1559_data_out(3);
    CN211_sign_in(26) <= VN1559_sign_out(3);
    CN211_data_in(27) <= VN1579_data_out(3);
    CN211_sign_in(27) <= VN1579_sign_out(3);
    CN211_data_in(28) <= VN1645_data_out(3);
    CN211_sign_in(28) <= VN1645_sign_out(3);
    CN211_data_in(29) <= VN1738_data_out(3);
    CN211_sign_in(29) <= VN1738_sign_out(3);
    CN211_data_in(30) <= VN1743_data_out(3);
    CN211_sign_in(30) <= VN1743_sign_out(3);
    CN211_data_in(31) <= VN1850_data_out(3);
    CN211_sign_in(31) <= VN1850_sign_out(3);
    CN212_data_in(0) <= VN34_data_out(3);
    CN212_sign_in(0) <= VN34_sign_out(3);
    CN212_data_in(1) <= VN65_data_out(3);
    CN212_sign_in(1) <= VN65_sign_out(3);
    CN212_data_in(2) <= VN163_data_out(3);
    CN212_sign_in(2) <= VN163_sign_out(3);
    CN212_data_in(3) <= VN186_data_out(3);
    CN212_sign_in(3) <= VN186_sign_out(3);
    CN212_data_in(4) <= VN296_data_out(3);
    CN212_sign_in(4) <= VN296_sign_out(3);
    CN212_data_in(5) <= VN405_data_out(3);
    CN212_sign_in(5) <= VN405_sign_out(3);
    CN212_data_in(6) <= VN541_data_out(3);
    CN212_sign_in(6) <= VN541_sign_out(3);
    CN212_data_in(7) <= VN683_data_out(3);
    CN212_sign_in(7) <= VN683_sign_out(3);
    CN212_data_in(8) <= VN827_data_out(3);
    CN212_sign_in(8) <= VN827_sign_out(3);
    CN212_data_in(9) <= VN999_data_out(3);
    CN212_sign_in(9) <= VN999_sign_out(3);
    CN212_data_in(10) <= VN1025_data_out(3);
    CN212_sign_in(10) <= VN1025_sign_out(3);
    CN212_data_in(11) <= VN1080_data_out(3);
    CN212_sign_in(11) <= VN1080_sign_out(3);
    CN212_data_in(12) <= VN1117_data_out(3);
    CN212_sign_in(12) <= VN1117_sign_out(3);
    CN212_data_in(13) <= VN1267_data_out(3);
    CN212_sign_in(13) <= VN1267_sign_out(3);
    CN212_data_in(14) <= VN1372_data_out(3);
    CN212_sign_in(14) <= VN1372_sign_out(3);
    CN212_data_in(15) <= VN1395_data_out(3);
    CN212_sign_in(15) <= VN1395_sign_out(3);
    CN212_data_in(16) <= VN1488_data_out(3);
    CN212_sign_in(16) <= VN1488_sign_out(3);
    CN212_data_in(17) <= VN1566_data_out(3);
    CN212_sign_in(17) <= VN1566_sign_out(3);
    CN212_data_in(18) <= VN1712_data_out(3);
    CN212_sign_in(18) <= VN1712_sign_out(3);
    CN212_data_in(19) <= VN1730_data_out(3);
    CN212_sign_in(19) <= VN1730_sign_out(3);
    CN212_data_in(20) <= VN1737_data_out(3);
    CN212_sign_in(20) <= VN1737_sign_out(3);
    CN212_data_in(21) <= VN1796_data_out(3);
    CN212_sign_in(21) <= VN1796_sign_out(3);
    CN212_data_in(22) <= VN1865_data_out(3);
    CN212_sign_in(22) <= VN1865_sign_out(3);
    CN212_data_in(23) <= VN1875_data_out(3);
    CN212_sign_in(23) <= VN1875_sign_out(3);
    CN212_data_in(24) <= VN1895_data_out(3);
    CN212_sign_in(24) <= VN1895_sign_out(3);
    CN212_data_in(25) <= VN1896_data_out(3);
    CN212_sign_in(25) <= VN1896_sign_out(3);
    CN212_data_in(26) <= VN1898_data_out(3);
    CN212_sign_in(26) <= VN1898_sign_out(3);
    CN212_data_in(27) <= VN1900_data_out(3);
    CN212_sign_in(27) <= VN1900_sign_out(3);
    CN212_data_in(28) <= VN1902_data_out(3);
    CN212_sign_in(28) <= VN1902_sign_out(3);
    CN212_data_in(29) <= VN1905_data_out(3);
    CN212_sign_in(29) <= VN1905_sign_out(3);
    CN212_data_in(30) <= VN1934_data_out(3);
    CN212_sign_in(30) <= VN1934_sign_out(3);
    CN212_data_in(31) <= VN1945_data_out(3);
    CN212_sign_in(31) <= VN1945_sign_out(3);
    CN213_data_in(0) <= VN33_data_out(3);
    CN213_sign_in(0) <= VN33_sign_out(3);
    CN213_data_in(1) <= VN71_data_out(3);
    CN213_sign_in(1) <= VN71_sign_out(3);
    CN213_data_in(2) <= VN142_data_out(3);
    CN213_sign_in(2) <= VN142_sign_out(3);
    CN213_data_in(3) <= VN230_data_out(3);
    CN213_sign_in(3) <= VN230_sign_out(3);
    CN213_data_in(4) <= VN389_data_out(3);
    CN213_sign_in(4) <= VN389_sign_out(3);
    CN213_data_in(5) <= VN503_data_out(3);
    CN213_sign_in(5) <= VN503_sign_out(3);
    CN213_data_in(6) <= VN583_data_out(3);
    CN213_sign_in(6) <= VN583_sign_out(3);
    CN213_data_in(7) <= VN631_data_out(3);
    CN213_sign_in(7) <= VN631_sign_out(3);
    CN213_data_in(8) <= VN767_data_out(3);
    CN213_sign_in(8) <= VN767_sign_out(3);
    CN213_data_in(9) <= VN848_data_out(3);
    CN213_sign_in(9) <= VN848_sign_out(3);
    CN213_data_in(10) <= VN916_data_out(3);
    CN213_sign_in(10) <= VN916_sign_out(3);
    CN213_data_in(11) <= VN987_data_out(3);
    CN213_sign_in(11) <= VN987_sign_out(3);
    CN213_data_in(12) <= VN1045_data_out(3);
    CN213_sign_in(12) <= VN1045_sign_out(3);
    CN213_data_in(13) <= VN1103_data_out(3);
    CN213_sign_in(13) <= VN1103_sign_out(3);
    CN213_data_in(14) <= VN1197_data_out(3);
    CN213_sign_in(14) <= VN1197_sign_out(3);
    CN213_data_in(15) <= VN1237_data_out(3);
    CN213_sign_in(15) <= VN1237_sign_out(3);
    CN213_data_in(16) <= VN1307_data_out(3);
    CN213_sign_in(16) <= VN1307_sign_out(3);
    CN213_data_in(17) <= VN1330_data_out(3);
    CN213_sign_in(17) <= VN1330_sign_out(3);
    CN213_data_in(18) <= VN1423_data_out(3);
    CN213_sign_in(18) <= VN1423_sign_out(3);
    CN213_data_in(19) <= VN1639_data_out(3);
    CN213_sign_in(19) <= VN1639_sign_out(3);
    CN213_data_in(20) <= VN1680_data_out(3);
    CN213_sign_in(20) <= VN1680_sign_out(3);
    CN213_data_in(21) <= VN1692_data_out(3);
    CN213_sign_in(21) <= VN1692_sign_out(3);
    CN213_data_in(22) <= VN1915_data_out(3);
    CN213_sign_in(22) <= VN1915_sign_out(3);
    CN213_data_in(23) <= VN1918_data_out(3);
    CN213_sign_in(23) <= VN1918_sign_out(3);
    CN213_data_in(24) <= VN1957_data_out(3);
    CN213_sign_in(24) <= VN1957_sign_out(3);
    CN213_data_in(25) <= VN1974_data_out(3);
    CN213_sign_in(25) <= VN1974_sign_out(3);
    CN213_data_in(26) <= VN1975_data_out(3);
    CN213_sign_in(26) <= VN1975_sign_out(3);
    CN213_data_in(27) <= VN2002_data_out(3);
    CN213_sign_in(27) <= VN2002_sign_out(3);
    CN213_data_in(28) <= VN2012_data_out(3);
    CN213_sign_in(28) <= VN2012_sign_out(3);
    CN213_data_in(29) <= VN2018_data_out(3);
    CN213_sign_in(29) <= VN2018_sign_out(3);
    CN213_data_in(30) <= VN2021_data_out(3);
    CN213_sign_in(30) <= VN2021_sign_out(3);
    CN213_data_in(31) <= VN2037_data_out(3);
    CN213_sign_in(31) <= VN2037_sign_out(3);
    CN214_data_in(0) <= VN32_data_out(3);
    CN214_sign_in(0) <= VN32_sign_out(3);
    CN214_data_in(1) <= VN59_data_out(3);
    CN214_sign_in(1) <= VN59_sign_out(3);
    CN214_data_in(2) <= VN145_data_out(3);
    CN214_sign_in(2) <= VN145_sign_out(3);
    CN214_data_in(3) <= VN220_data_out(3);
    CN214_sign_in(3) <= VN220_sign_out(3);
    CN214_data_in(4) <= VN240_data_out(3);
    CN214_sign_in(4) <= VN240_sign_out(3);
    CN214_data_in(5) <= VN308_data_out(3);
    CN214_sign_in(5) <= VN308_sign_out(3);
    CN214_data_in(6) <= VN369_data_out(3);
    CN214_sign_in(6) <= VN369_sign_out(3);
    CN214_data_in(7) <= VN445_data_out(3);
    CN214_sign_in(7) <= VN445_sign_out(3);
    CN214_data_in(8) <= VN451_data_out(3);
    CN214_sign_in(8) <= VN451_sign_out(3);
    CN214_data_in(9) <= VN515_data_out(3);
    CN214_sign_in(9) <= VN515_sign_out(3);
    CN214_data_in(10) <= VN615_data_out(3);
    CN214_sign_in(10) <= VN615_sign_out(3);
    CN214_data_in(11) <= VN661_data_out(3);
    CN214_sign_in(11) <= VN661_sign_out(3);
    CN214_data_in(12) <= VN674_data_out(3);
    CN214_sign_in(12) <= VN674_sign_out(3);
    CN214_data_in(13) <= VN764_data_out(3);
    CN214_sign_in(13) <= VN764_sign_out(3);
    CN214_data_in(14) <= VN806_data_out(3);
    CN214_sign_in(14) <= VN806_sign_out(3);
    CN214_data_in(15) <= VN852_data_out(3);
    CN214_sign_in(15) <= VN852_sign_out(3);
    CN214_data_in(16) <= VN940_data_out(3);
    CN214_sign_in(16) <= VN940_sign_out(3);
    CN214_data_in(17) <= VN973_data_out(3);
    CN214_sign_in(17) <= VN973_sign_out(3);
    CN214_data_in(18) <= VN1055_data_out(3);
    CN214_sign_in(18) <= VN1055_sign_out(3);
    CN214_data_in(19) <= VN1095_data_out(3);
    CN214_sign_in(19) <= VN1095_sign_out(3);
    CN214_data_in(20) <= VN1130_data_out(3);
    CN214_sign_in(20) <= VN1130_sign_out(3);
    CN214_data_in(21) <= VN1209_data_out(3);
    CN214_sign_in(21) <= VN1209_sign_out(3);
    CN214_data_in(22) <= VN1274_data_out(3);
    CN214_sign_in(22) <= VN1274_sign_out(3);
    CN214_data_in(23) <= VN1295_data_out(3);
    CN214_sign_in(23) <= VN1295_sign_out(3);
    CN214_data_in(24) <= VN1353_data_out(3);
    CN214_sign_in(24) <= VN1353_sign_out(3);
    CN214_data_in(25) <= VN1402_data_out(3);
    CN214_sign_in(25) <= VN1402_sign_out(3);
    CN214_data_in(26) <= VN1453_data_out(3);
    CN214_sign_in(26) <= VN1453_sign_out(3);
    CN214_data_in(27) <= VN1461_data_out(3);
    CN214_sign_in(27) <= VN1461_sign_out(3);
    CN214_data_in(28) <= VN1472_data_out(3);
    CN214_sign_in(28) <= VN1472_sign_out(3);
    CN214_data_in(29) <= VN1623_data_out(3);
    CN214_sign_in(29) <= VN1623_sign_out(3);
    CN214_data_in(30) <= VN1677_data_out(3);
    CN214_sign_in(30) <= VN1677_sign_out(3);
    CN214_data_in(31) <= VN1774_data_out(3);
    CN214_sign_in(31) <= VN1774_sign_out(3);
    CN215_data_in(0) <= VN31_data_out(3);
    CN215_sign_in(0) <= VN31_sign_out(3);
    CN215_data_in(1) <= VN85_data_out(3);
    CN215_sign_in(1) <= VN85_sign_out(3);
    CN215_data_in(2) <= VN130_data_out(3);
    CN215_sign_in(2) <= VN130_sign_out(3);
    CN215_data_in(3) <= VN216_data_out(3);
    CN215_sign_in(3) <= VN216_sign_out(3);
    CN215_data_in(4) <= VN234_data_out(3);
    CN215_sign_in(4) <= VN234_sign_out(3);
    CN215_data_in(5) <= VN311_data_out(3);
    CN215_sign_in(5) <= VN311_sign_out(3);
    CN215_data_in(6) <= VN377_data_out(3);
    CN215_sign_in(6) <= VN377_sign_out(3);
    CN215_data_in(7) <= VN446_data_out(3);
    CN215_sign_in(7) <= VN446_sign_out(3);
    CN215_data_in(8) <= VN505_data_out(3);
    CN215_sign_in(8) <= VN505_sign_out(3);
    CN215_data_in(9) <= VN556_data_out(3);
    CN215_sign_in(9) <= VN556_sign_out(3);
    CN215_data_in(10) <= VN607_data_out(3);
    CN215_sign_in(10) <= VN607_sign_out(3);
    CN215_data_in(11) <= VN621_data_out(3);
    CN215_sign_in(11) <= VN621_sign_out(3);
    CN215_data_in(12) <= VN676_data_out(3);
    CN215_sign_in(12) <= VN676_sign_out(3);
    CN215_data_in(13) <= VN724_data_out(3);
    CN215_sign_in(13) <= VN724_sign_out(3);
    CN215_data_in(14) <= VN825_data_out(3);
    CN215_sign_in(14) <= VN825_sign_out(3);
    CN215_data_in(15) <= VN841_data_out(3);
    CN215_sign_in(15) <= VN841_sign_out(3);
    CN215_data_in(16) <= VN922_data_out(3);
    CN215_sign_in(16) <= VN922_sign_out(3);
    CN215_data_in(17) <= VN990_data_out(3);
    CN215_sign_in(17) <= VN990_sign_out(3);
    CN215_data_in(18) <= VN1050_data_out(3);
    CN215_sign_in(18) <= VN1050_sign_out(3);
    CN215_data_in(19) <= VN1085_data_out(3);
    CN215_sign_in(19) <= VN1085_sign_out(3);
    CN215_data_in(20) <= VN1137_data_out(3);
    CN215_sign_in(20) <= VN1137_sign_out(3);
    CN215_data_in(21) <= VN1215_data_out(3);
    CN215_sign_in(21) <= VN1215_sign_out(3);
    CN215_data_in(22) <= VN1224_data_out(3);
    CN215_sign_in(22) <= VN1224_sign_out(3);
    CN215_data_in(23) <= VN1230_data_out(3);
    CN215_sign_in(23) <= VN1230_sign_out(3);
    CN215_data_in(24) <= VN1317_data_out(3);
    CN215_sign_in(24) <= VN1317_sign_out(3);
    CN215_data_in(25) <= VN1361_data_out(3);
    CN215_sign_in(25) <= VN1361_sign_out(3);
    CN215_data_in(26) <= VN1387_data_out(3);
    CN215_sign_in(26) <= VN1387_sign_out(3);
    CN215_data_in(27) <= VN1425_data_out(3);
    CN215_sign_in(27) <= VN1425_sign_out(3);
    CN215_data_in(28) <= VN1601_data_out(3);
    CN215_sign_in(28) <= VN1601_sign_out(3);
    CN215_data_in(29) <= VN1608_data_out(3);
    CN215_sign_in(29) <= VN1608_sign_out(3);
    CN215_data_in(30) <= VN1651_data_out(3);
    CN215_sign_in(30) <= VN1651_sign_out(3);
    CN215_data_in(31) <= VN1775_data_out(3);
    CN215_sign_in(31) <= VN1775_sign_out(3);
    CN216_data_in(0) <= VN30_data_out(3);
    CN216_sign_in(0) <= VN30_sign_out(3);
    CN216_data_in(1) <= VN91_data_out(3);
    CN216_sign_in(1) <= VN91_sign_out(3);
    CN216_data_in(2) <= VN164_data_out(3);
    CN216_sign_in(2) <= VN164_sign_out(3);
    CN216_data_in(3) <= VN183_data_out(3);
    CN216_sign_in(3) <= VN183_sign_out(3);
    CN216_data_in(4) <= VN237_data_out(3);
    CN216_sign_in(4) <= VN237_sign_out(3);
    CN216_data_in(5) <= VN299_data_out(3);
    CN216_sign_in(5) <= VN299_sign_out(3);
    CN216_data_in(6) <= VN341_data_out(3);
    CN216_sign_in(6) <= VN341_sign_out(3);
    CN216_data_in(7) <= VN423_data_out(3);
    CN216_sign_in(7) <= VN423_sign_out(3);
    CN216_data_in(8) <= VN450_data_out(3);
    CN216_sign_in(8) <= VN450_sign_out(3);
    CN216_data_in(9) <= VN558_data_out(3);
    CN216_sign_in(9) <= VN558_sign_out(3);
    CN216_data_in(10) <= VN649_data_out(3);
    CN216_sign_in(10) <= VN649_sign_out(3);
    CN216_data_in(11) <= VN701_data_out(3);
    CN216_sign_in(11) <= VN701_sign_out(3);
    CN216_data_in(12) <= VN772_data_out(3);
    CN216_sign_in(12) <= VN772_sign_out(3);
    CN216_data_in(13) <= VN876_data_out(3);
    CN216_sign_in(13) <= VN876_sign_out(3);
    CN216_data_in(14) <= VN932_data_out(3);
    CN216_sign_in(14) <= VN932_sign_out(3);
    CN216_data_in(15) <= VN951_data_out(3);
    CN216_sign_in(15) <= VN951_sign_out(3);
    CN216_data_in(16) <= VN1056_data_out(3);
    CN216_sign_in(16) <= VN1056_sign_out(3);
    CN216_data_in(17) <= VN1100_data_out(3);
    CN216_sign_in(17) <= VN1100_sign_out(3);
    CN216_data_in(18) <= VN1108_data_out(3);
    CN216_sign_in(18) <= VN1108_sign_out(3);
    CN216_data_in(19) <= VN1121_data_out(3);
    CN216_sign_in(19) <= VN1121_sign_out(3);
    CN216_data_in(20) <= VN1191_data_out(3);
    CN216_sign_in(20) <= VN1191_sign_out(3);
    CN216_data_in(21) <= VN1238_data_out(3);
    CN216_sign_in(21) <= VN1238_sign_out(3);
    CN216_data_in(22) <= VN1309_data_out(3);
    CN216_sign_in(22) <= VN1309_sign_out(3);
    CN216_data_in(23) <= VN1357_data_out(3);
    CN216_sign_in(23) <= VN1357_sign_out(3);
    CN216_data_in(24) <= VN1546_data_out(3);
    CN216_sign_in(24) <= VN1546_sign_out(3);
    CN216_data_in(25) <= VN1561_data_out(3);
    CN216_sign_in(25) <= VN1561_sign_out(3);
    CN216_data_in(26) <= VN1618_data_out(3);
    CN216_sign_in(26) <= VN1618_sign_out(3);
    CN216_data_in(27) <= VN1713_data_out(3);
    CN216_sign_in(27) <= VN1713_sign_out(3);
    CN216_data_in(28) <= VN1766_data_out(3);
    CN216_sign_in(28) <= VN1766_sign_out(3);
    CN216_data_in(29) <= VN1797_data_out(3);
    CN216_sign_in(29) <= VN1797_sign_out(3);
    CN216_data_in(30) <= VN1821_data_out(3);
    CN216_sign_in(30) <= VN1821_sign_out(3);
    CN216_data_in(31) <= VN1888_data_out(3);
    CN216_sign_in(31) <= VN1888_sign_out(3);
    CN217_data_in(0) <= VN29_data_out(3);
    CN217_sign_in(0) <= VN29_sign_out(3);
    CN217_data_in(1) <= VN75_data_out(3);
    CN217_sign_in(1) <= VN75_sign_out(3);
    CN217_data_in(2) <= VN126_data_out(3);
    CN217_sign_in(2) <= VN126_sign_out(3);
    CN217_data_in(3) <= VN201_data_out(3);
    CN217_sign_in(3) <= VN201_sign_out(3);
    CN217_data_in(4) <= VN227_data_out(3);
    CN217_sign_in(4) <= VN227_sign_out(3);
    CN217_data_in(5) <= VN329_data_out(3);
    CN217_sign_in(5) <= VN329_sign_out(3);
    CN217_data_in(6) <= VN339_data_out(3);
    CN217_sign_in(6) <= VN339_sign_out(3);
    CN217_data_in(7) <= VN414_data_out(3);
    CN217_sign_in(7) <= VN414_sign_out(3);
    CN217_data_in(8) <= VN501_data_out(3);
    CN217_sign_in(8) <= VN501_sign_out(3);
    CN217_data_in(9) <= VN524_data_out(3);
    CN217_sign_in(9) <= VN524_sign_out(3);
    CN217_data_in(10) <= VN574_data_out(3);
    CN217_sign_in(10) <= VN574_sign_out(3);
    CN217_data_in(11) <= VN627_data_out(3);
    CN217_sign_in(11) <= VN627_sign_out(3);
    CN217_data_in(12) <= VN681_data_out(3);
    CN217_sign_in(12) <= VN681_sign_out(3);
    CN217_data_in(13) <= VN747_data_out(3);
    CN217_sign_in(13) <= VN747_sign_out(3);
    CN217_data_in(14) <= VN797_data_out(3);
    CN217_sign_in(14) <= VN797_sign_out(3);
    CN217_data_in(15) <= VN860_data_out(3);
    CN217_sign_in(15) <= VN860_sign_out(3);
    CN217_data_in(16) <= VN941_data_out(3);
    CN217_sign_in(16) <= VN941_sign_out(3);
    CN217_data_in(17) <= VN961_data_out(3);
    CN217_sign_in(17) <= VN961_sign_out(3);
    CN217_data_in(18) <= VN1044_data_out(3);
    CN217_sign_in(18) <= VN1044_sign_out(3);
    CN217_data_in(19) <= VN1078_data_out(3);
    CN217_sign_in(19) <= VN1078_sign_out(3);
    CN217_data_in(20) <= VN1122_data_out(3);
    CN217_sign_in(20) <= VN1122_sign_out(3);
    CN217_data_in(21) <= VN1204_data_out(3);
    CN217_sign_in(21) <= VN1204_sign_out(3);
    CN217_data_in(22) <= VN1266_data_out(3);
    CN217_sign_in(22) <= VN1266_sign_out(3);
    CN217_data_in(23) <= VN1299_data_out(3);
    CN217_sign_in(23) <= VN1299_sign_out(3);
    CN217_data_in(24) <= VN1332_data_out(3);
    CN217_sign_in(24) <= VN1332_sign_out(3);
    CN217_data_in(25) <= VN1362_data_out(3);
    CN217_sign_in(25) <= VN1362_sign_out(3);
    CN217_data_in(26) <= VN1389_data_out(3);
    CN217_sign_in(26) <= VN1389_sign_out(3);
    CN217_data_in(27) <= VN1542_data_out(3);
    CN217_sign_in(27) <= VN1542_sign_out(3);
    CN217_data_in(28) <= VN1606_data_out(3);
    CN217_sign_in(28) <= VN1606_sign_out(3);
    CN217_data_in(29) <= VN1628_data_out(3);
    CN217_sign_in(29) <= VN1628_sign_out(3);
    CN217_data_in(30) <= VN1667_data_out(3);
    CN217_sign_in(30) <= VN1667_sign_out(3);
    CN217_data_in(31) <= VN1776_data_out(3);
    CN217_sign_in(31) <= VN1776_sign_out(3);
    CN218_data_in(0) <= VN28_data_out(3);
    CN218_sign_in(0) <= VN28_sign_out(3);
    CN218_data_in(1) <= VN77_data_out(3);
    CN218_sign_in(1) <= VN77_sign_out(3);
    CN218_data_in(2) <= VN154_data_out(3);
    CN218_sign_in(2) <= VN154_sign_out(3);
    CN218_data_in(3) <= VN202_data_out(3);
    CN218_sign_in(3) <= VN202_sign_out(3);
    CN218_data_in(4) <= VN261_data_out(3);
    CN218_sign_in(4) <= VN261_sign_out(3);
    CN218_data_in(5) <= VN295_data_out(3);
    CN218_sign_in(5) <= VN295_sign_out(3);
    CN218_data_in(6) <= VN375_data_out(3);
    CN218_sign_in(6) <= VN375_sign_out(3);
    CN218_data_in(7) <= VN432_data_out(3);
    CN218_sign_in(7) <= VN432_sign_out(3);
    CN218_data_in(8) <= VN483_data_out(3);
    CN218_sign_in(8) <= VN483_sign_out(3);
    CN218_data_in(9) <= VN508_data_out(3);
    CN218_sign_in(9) <= VN508_sign_out(3);
    CN218_data_in(10) <= VN616_data_out(3);
    CN218_sign_in(10) <= VN616_sign_out(3);
    CN218_data_in(11) <= VN651_data_out(3);
    CN218_sign_in(11) <= VN651_sign_out(3);
    CN218_data_in(12) <= VN693_data_out(3);
    CN218_sign_in(12) <= VN693_sign_out(3);
    CN218_data_in(13) <= VN757_data_out(3);
    CN218_sign_in(13) <= VN757_sign_out(3);
    CN218_data_in(14) <= VN811_data_out(3);
    CN218_sign_in(14) <= VN811_sign_out(3);
    CN218_data_in(15) <= VN871_data_out(3);
    CN218_sign_in(15) <= VN871_sign_out(3);
    CN218_data_in(16) <= VN915_data_out(3);
    CN218_sign_in(16) <= VN915_sign_out(3);
    CN218_data_in(17) <= VN956_data_out(3);
    CN218_sign_in(17) <= VN956_sign_out(3);
    CN218_data_in(18) <= VN1013_data_out(3);
    CN218_sign_in(18) <= VN1013_sign_out(3);
    CN218_data_in(19) <= VN1076_data_out(3);
    CN218_sign_in(19) <= VN1076_sign_out(3);
    CN218_data_in(20) <= VN1148_data_out(3);
    CN218_sign_in(20) <= VN1148_sign_out(3);
    CN218_data_in(21) <= VN1177_data_out(3);
    CN218_sign_in(21) <= VN1177_sign_out(3);
    CN218_data_in(22) <= VN1225_data_out(3);
    CN218_sign_in(22) <= VN1225_sign_out(3);
    CN218_data_in(23) <= VN1277_data_out(3);
    CN218_sign_in(23) <= VN1277_sign_out(3);
    CN218_data_in(24) <= VN1313_data_out(3);
    CN218_sign_in(24) <= VN1313_sign_out(3);
    CN218_data_in(25) <= VN1352_data_out(3);
    CN218_sign_in(25) <= VN1352_sign_out(3);
    CN218_data_in(26) <= VN1397_data_out(3);
    CN218_sign_in(26) <= VN1397_sign_out(3);
    CN218_data_in(27) <= VN1436_data_out(3);
    CN218_sign_in(27) <= VN1436_sign_out(3);
    CN218_data_in(28) <= VN1492_data_out(3);
    CN218_sign_in(28) <= VN1492_sign_out(3);
    CN218_data_in(29) <= VN1586_data_out(3);
    CN218_sign_in(29) <= VN1586_sign_out(3);
    CN218_data_in(30) <= VN1698_data_out(3);
    CN218_sign_in(30) <= VN1698_sign_out(3);
    CN218_data_in(31) <= VN1777_data_out(3);
    CN218_sign_in(31) <= VN1777_sign_out(3);
    CN219_data_in(0) <= VN27_data_out(3);
    CN219_sign_in(0) <= VN27_sign_out(3);
    CN219_data_in(1) <= VN101_data_out(3);
    CN219_sign_in(1) <= VN101_sign_out(3);
    CN219_data_in(2) <= VN138_data_out(3);
    CN219_sign_in(2) <= VN138_sign_out(3);
    CN219_data_in(3) <= VN182_data_out(3);
    CN219_sign_in(3) <= VN182_sign_out(3);
    CN219_data_in(4) <= VN321_data_out(3);
    CN219_sign_in(4) <= VN321_sign_out(3);
    CN219_data_in(5) <= VN354_data_out(3);
    CN219_sign_in(5) <= VN354_sign_out(3);
    CN219_data_in(6) <= VN437_data_out(3);
    CN219_sign_in(6) <= VN437_sign_out(3);
    CN219_data_in(7) <= VN489_data_out(3);
    CN219_sign_in(7) <= VN489_sign_out(3);
    CN219_data_in(8) <= VN518_data_out(3);
    CN219_sign_in(8) <= VN518_sign_out(3);
    CN219_data_in(9) <= VN573_data_out(3);
    CN219_sign_in(9) <= VN573_sign_out(3);
    CN219_data_in(10) <= VN663_data_out(3);
    CN219_sign_in(10) <= VN663_sign_out(3);
    CN219_data_in(11) <= VN702_data_out(3);
    CN219_sign_in(11) <= VN702_sign_out(3);
    CN219_data_in(12) <= VN750_data_out(3);
    CN219_sign_in(12) <= VN750_sign_out(3);
    CN219_data_in(13) <= VN804_data_out(3);
    CN219_sign_in(13) <= VN804_sign_out(3);
    CN219_data_in(14) <= VN882_data_out(3);
    CN219_sign_in(14) <= VN882_sign_out(3);
    CN219_data_in(15) <= VN929_data_out(3);
    CN219_sign_in(15) <= VN929_sign_out(3);
    CN219_data_in(16) <= VN962_data_out(3);
    CN219_sign_in(16) <= VN962_sign_out(3);
    CN219_data_in(17) <= VN1019_data_out(3);
    CN219_sign_in(17) <= VN1019_sign_out(3);
    CN219_data_in(18) <= VN1089_data_out(3);
    CN219_sign_in(18) <= VN1089_sign_out(3);
    CN219_data_in(19) <= VN1129_data_out(3);
    CN219_sign_in(19) <= VN1129_sign_out(3);
    CN219_data_in(20) <= VN1165_data_out(3);
    CN219_sign_in(20) <= VN1165_sign_out(3);
    CN219_data_in(21) <= VN1212_data_out(3);
    CN219_sign_in(21) <= VN1212_sign_out(3);
    CN219_data_in(22) <= VN1253_data_out(3);
    CN219_sign_in(22) <= VN1253_sign_out(3);
    CN219_data_in(23) <= VN1292_data_out(3);
    CN219_sign_in(23) <= VN1292_sign_out(3);
    CN219_data_in(24) <= VN1375_data_out(3);
    CN219_sign_in(24) <= VN1375_sign_out(3);
    CN219_data_in(25) <= VN1419_data_out(3);
    CN219_sign_in(25) <= VN1419_sign_out(3);
    CN219_data_in(26) <= VN1433_data_out(3);
    CN219_sign_in(26) <= VN1433_sign_out(3);
    CN219_data_in(27) <= VN1641_data_out(3);
    CN219_sign_in(27) <= VN1641_sign_out(3);
    CN219_data_in(28) <= VN1705_data_out(3);
    CN219_sign_in(28) <= VN1705_sign_out(3);
    CN219_data_in(29) <= VN1757_data_out(3);
    CN219_sign_in(29) <= VN1757_sign_out(3);
    CN219_data_in(30) <= VN1801_data_out(3);
    CN219_sign_in(30) <= VN1801_sign_out(3);
    CN219_data_in(31) <= VN1851_data_out(3);
    CN219_sign_in(31) <= VN1851_sign_out(3);
    CN220_data_in(0) <= VN26_data_out(3);
    CN220_sign_in(0) <= VN26_sign_out(3);
    CN220_data_in(1) <= VN83_data_out(3);
    CN220_sign_in(1) <= VN83_sign_out(3);
    CN220_data_in(2) <= VN166_data_out(3);
    CN220_sign_in(2) <= VN166_sign_out(3);
    CN220_data_in(3) <= VN173_data_out(3);
    CN220_sign_in(3) <= VN173_sign_out(3);
    CN220_data_in(4) <= VN256_data_out(3);
    CN220_sign_in(4) <= VN256_sign_out(3);
    CN220_data_in(5) <= VN305_data_out(3);
    CN220_sign_in(5) <= VN305_sign_out(3);
    CN220_data_in(6) <= VN356_data_out(3);
    CN220_sign_in(6) <= VN356_sign_out(3);
    CN220_data_in(7) <= VN447_data_out(3);
    CN220_sign_in(7) <= VN447_sign_out(3);
    CN220_data_in(8) <= VN457_data_out(3);
    CN220_sign_in(8) <= VN457_sign_out(3);
    CN220_data_in(9) <= VN525_data_out(3);
    CN220_sign_in(9) <= VN525_sign_out(3);
    CN220_data_in(10) <= VN568_data_out(3);
    CN220_sign_in(10) <= VN568_sign_out(3);
    CN220_data_in(11) <= VN659_data_out(3);
    CN220_sign_in(11) <= VN659_sign_out(3);
    CN220_data_in(12) <= VN675_data_out(3);
    CN220_sign_in(12) <= VN675_sign_out(3);
    CN220_data_in(13) <= VN754_data_out(3);
    CN220_sign_in(13) <= VN754_sign_out(3);
    CN220_data_in(14) <= VN781_data_out(3);
    CN220_sign_in(14) <= VN781_sign_out(3);
    CN220_data_in(15) <= VN855_data_out(3);
    CN220_sign_in(15) <= VN855_sign_out(3);
    CN220_data_in(16) <= VN902_data_out(3);
    CN220_sign_in(16) <= VN902_sign_out(3);
    CN220_data_in(17) <= VN950_data_out(3);
    CN220_sign_in(17) <= VN950_sign_out(3);
    CN220_data_in(18) <= VN1004_data_out(3);
    CN220_sign_in(18) <= VN1004_sign_out(3);
    CN220_data_in(19) <= VN1082_data_out(3);
    CN220_sign_in(19) <= VN1082_sign_out(3);
    CN220_data_in(20) <= VN1140_data_out(3);
    CN220_sign_in(20) <= VN1140_sign_out(3);
    CN220_data_in(21) <= VN1179_data_out(3);
    CN220_sign_in(21) <= VN1179_sign_out(3);
    CN220_data_in(22) <= VN1233_data_out(3);
    CN220_sign_in(22) <= VN1233_sign_out(3);
    CN220_data_in(23) <= VN1282_data_out(3);
    CN220_sign_in(23) <= VN1282_sign_out(3);
    CN220_data_in(24) <= VN1289_data_out(3);
    CN220_sign_in(24) <= VN1289_sign_out(3);
    CN220_data_in(25) <= VN1381_data_out(3);
    CN220_sign_in(25) <= VN1381_sign_out(3);
    CN220_data_in(26) <= VN1420_data_out(3);
    CN220_sign_in(26) <= VN1420_sign_out(3);
    CN220_data_in(27) <= VN1475_data_out(3);
    CN220_sign_in(27) <= VN1475_sign_out(3);
    CN220_data_in(28) <= VN1594_data_out(3);
    CN220_sign_in(28) <= VN1594_sign_out(3);
    CN220_data_in(29) <= VN1629_data_out(3);
    CN220_sign_in(29) <= VN1629_sign_out(3);
    CN220_data_in(30) <= VN1656_data_out(3);
    CN220_sign_in(30) <= VN1656_sign_out(3);
    CN220_data_in(31) <= VN1778_data_out(3);
    CN220_sign_in(31) <= VN1778_sign_out(3);
    CN221_data_in(0) <= VN25_data_out(3);
    CN221_sign_in(0) <= VN25_sign_out(3);
    CN221_data_in(1) <= VN94_data_out(3);
    CN221_sign_in(1) <= VN94_sign_out(3);
    CN221_data_in(2) <= VN156_data_out(3);
    CN221_sign_in(2) <= VN156_sign_out(3);
    CN221_data_in(3) <= VN190_data_out(3);
    CN221_sign_in(3) <= VN190_sign_out(3);
    CN221_data_in(4) <= VN268_data_out(3);
    CN221_sign_in(4) <= VN268_sign_out(3);
    CN221_data_in(5) <= VN331_data_out(3);
    CN221_sign_in(5) <= VN331_sign_out(3);
    CN221_data_in(6) <= VN342_data_out(3);
    CN221_sign_in(6) <= VN342_sign_out(3);
    CN221_data_in(7) <= VN436_data_out(3);
    CN221_sign_in(7) <= VN436_sign_out(3);
    CN221_data_in(8) <= VN455_data_out(3);
    CN221_sign_in(8) <= VN455_sign_out(3);
    CN221_data_in(9) <= VN557_data_out(3);
    CN221_sign_in(9) <= VN557_sign_out(3);
    CN221_data_in(10) <= VN604_data_out(3);
    CN221_sign_in(10) <= VN604_sign_out(3);
    CN221_data_in(11) <= VN624_data_out(3);
    CN221_sign_in(11) <= VN624_sign_out(3);
    CN221_data_in(12) <= VN689_data_out(3);
    CN221_sign_in(12) <= VN689_sign_out(3);
    CN221_data_in(13) <= VN791_data_out(3);
    CN221_sign_in(13) <= VN791_sign_out(3);
    CN221_data_in(14) <= VN843_data_out(3);
    CN221_sign_in(14) <= VN843_sign_out(3);
    CN221_data_in(15) <= VN935_data_out(3);
    CN221_sign_in(15) <= VN935_sign_out(3);
    CN221_data_in(16) <= VN976_data_out(3);
    CN221_sign_in(16) <= VN976_sign_out(3);
    CN221_data_in(17) <= VN1111_data_out(3);
    CN221_sign_in(17) <= VN1111_sign_out(3);
    CN221_data_in(18) <= VN1149_data_out(3);
    CN221_sign_in(18) <= VN1149_sign_out(3);
    CN221_data_in(19) <= VN1302_data_out(3);
    CN221_sign_in(19) <= VN1302_sign_out(3);
    CN221_data_in(20) <= VN1334_data_out(3);
    CN221_sign_in(20) <= VN1334_sign_out(3);
    CN221_data_in(21) <= VN1365_data_out(3);
    CN221_sign_in(21) <= VN1365_sign_out(3);
    CN221_data_in(22) <= VN1396_data_out(3);
    CN221_sign_in(22) <= VN1396_sign_out(3);
    CN221_data_in(23) <= VN1590_data_out(3);
    CN221_sign_in(23) <= VN1590_sign_out(3);
    CN221_data_in(24) <= VN1660_data_out(3);
    CN221_sign_in(24) <= VN1660_sign_out(3);
    CN221_data_in(25) <= VN1704_data_out(3);
    CN221_sign_in(25) <= VN1704_sign_out(3);
    CN221_data_in(26) <= VN1727_data_out(3);
    CN221_sign_in(26) <= VN1727_sign_out(3);
    CN221_data_in(27) <= VN1876_data_out(3);
    CN221_sign_in(27) <= VN1876_sign_out(3);
    CN221_data_in(28) <= VN1882_data_out(3);
    CN221_sign_in(28) <= VN1882_sign_out(3);
    CN221_data_in(29) <= VN1935_data_out(3);
    CN221_sign_in(29) <= VN1935_sign_out(3);
    CN221_data_in(30) <= VN1940_data_out(3);
    CN221_sign_in(30) <= VN1940_sign_out(3);
    CN221_data_in(31) <= VN1946_data_out(3);
    CN221_sign_in(31) <= VN1946_sign_out(3);
    CN222_data_in(0) <= VN24_data_out(3);
    CN222_sign_in(0) <= VN24_sign_out(3);
    CN222_data_in(1) <= VN143_data_out(3);
    CN222_sign_in(1) <= VN143_sign_out(3);
    CN222_data_in(2) <= VN241_data_out(3);
    CN222_sign_in(2) <= VN241_sign_out(3);
    CN222_data_in(3) <= VN376_data_out(3);
    CN222_sign_in(3) <= VN376_sign_out(3);
    CN222_data_in(4) <= VN430_data_out(3);
    CN222_sign_in(4) <= VN430_sign_out(3);
    CN222_data_in(5) <= VN487_data_out(3);
    CN222_sign_in(5) <= VN487_sign_out(3);
    CN222_data_in(6) <= VN611_data_out(3);
    CN222_sign_in(6) <= VN611_sign_out(3);
    CN222_data_in(7) <= VN644_data_out(3);
    CN222_sign_in(7) <= VN644_sign_out(3);
    CN222_data_in(8) <= VN777_data_out(3);
    CN222_sign_in(8) <= VN777_sign_out(3);
    CN222_data_in(9) <= VN885_data_out(3);
    CN222_sign_in(9) <= VN885_sign_out(3);
    CN222_data_in(10) <= VN904_data_out(3);
    CN222_sign_in(10) <= VN904_sign_out(3);
    CN222_data_in(11) <= VN982_data_out(3);
    CN222_sign_in(11) <= VN982_sign_out(3);
    CN222_data_in(12) <= VN1189_data_out(3);
    CN222_sign_in(12) <= VN1189_sign_out(3);
    CN222_data_in(13) <= VN1268_data_out(3);
    CN222_sign_in(13) <= VN1268_sign_out(3);
    CN222_data_in(14) <= VN1367_data_out(3);
    CN222_sign_in(14) <= VN1367_sign_out(3);
    CN222_data_in(15) <= VN1391_data_out(3);
    CN222_sign_in(15) <= VN1391_sign_out(3);
    CN222_data_in(16) <= VN1687_data_out(3);
    CN222_sign_in(16) <= VN1687_sign_out(3);
    CN222_data_in(17) <= VN1749_data_out(3);
    CN222_sign_in(17) <= VN1749_sign_out(3);
    CN222_data_in(18) <= VN1820_data_out(3);
    CN222_sign_in(18) <= VN1820_sign_out(3);
    CN222_data_in(19) <= VN1823_data_out(3);
    CN222_sign_in(19) <= VN1823_sign_out(3);
    CN222_data_in(20) <= VN1870_data_out(3);
    CN222_sign_in(20) <= VN1870_sign_out(3);
    CN222_data_in(21) <= VN1913_data_out(3);
    CN222_sign_in(21) <= VN1913_sign_out(3);
    CN222_data_in(22) <= VN1932_data_out(3);
    CN222_sign_in(22) <= VN1932_sign_out(3);
    CN222_data_in(23) <= VN1969_data_out(3);
    CN222_sign_in(23) <= VN1969_sign_out(3);
    CN222_data_in(24) <= VN1973_data_out(3);
    CN222_sign_in(24) <= VN1973_sign_out(3);
    CN222_data_in(25) <= VN1982_data_out(3);
    CN222_sign_in(25) <= VN1982_sign_out(3);
    CN222_data_in(26) <= VN2007_data_out(3);
    CN222_sign_in(26) <= VN2007_sign_out(3);
    CN222_data_in(27) <= VN2023_data_out(3);
    CN222_sign_in(27) <= VN2023_sign_out(3);
    CN222_data_in(28) <= VN2033_data_out(3);
    CN222_sign_in(28) <= VN2033_sign_out(3);
    CN222_data_in(29) <= VN2035_data_out(3);
    CN222_sign_in(29) <= VN2035_sign_out(3);
    CN222_data_in(30) <= VN2041_data_out(3);
    CN222_sign_in(30) <= VN2041_sign_out(3);
    CN222_data_in(31) <= VN2046_data_out(3);
    CN222_sign_in(31) <= VN2046_sign_out(3);
    CN223_data_in(0) <= VN23_data_out(3);
    CN223_sign_in(0) <= VN23_sign_out(3);
    CN223_data_in(1) <= VN76_data_out(3);
    CN223_sign_in(1) <= VN76_sign_out(3);
    CN223_data_in(2) <= VN162_data_out(3);
    CN223_sign_in(2) <= VN162_sign_out(3);
    CN223_data_in(3) <= VN224_data_out(3);
    CN223_sign_in(3) <= VN224_sign_out(3);
    CN223_data_in(4) <= VN229_data_out(3);
    CN223_sign_in(4) <= VN229_sign_out(3);
    CN223_data_in(5) <= VN309_data_out(3);
    CN223_sign_in(5) <= VN309_sign_out(3);
    CN223_data_in(6) <= VN338_data_out(3);
    CN223_sign_in(6) <= VN338_sign_out(3);
    CN223_data_in(7) <= VN411_data_out(3);
    CN223_sign_in(7) <= VN411_sign_out(3);
    CN223_data_in(8) <= VN469_data_out(3);
    CN223_sign_in(8) <= VN469_sign_out(3);
    CN223_data_in(9) <= VN543_data_out(3);
    CN223_sign_in(9) <= VN543_sign_out(3);
    CN223_data_in(10) <= VN579_data_out(3);
    CN223_sign_in(10) <= VN579_sign_out(3);
    CN223_data_in(11) <= VN645_data_out(3);
    CN223_sign_in(11) <= VN645_sign_out(3);
    CN223_data_in(12) <= VN696_data_out(3);
    CN223_sign_in(12) <= VN696_sign_out(3);
    CN223_data_in(13) <= VN788_data_out(3);
    CN223_sign_in(13) <= VN788_sign_out(3);
    CN223_data_in(14) <= VN846_data_out(3);
    CN223_sign_in(14) <= VN846_sign_out(3);
    CN223_data_in(15) <= VN917_data_out(3);
    CN223_sign_in(15) <= VN917_sign_out(3);
    CN223_data_in(16) <= VN965_data_out(3);
    CN223_sign_in(16) <= VN965_sign_out(3);
    CN223_data_in(17) <= VN1011_data_out(3);
    CN223_sign_in(17) <= VN1011_sign_out(3);
    CN223_data_in(18) <= VN1062_data_out(3);
    CN223_sign_in(18) <= VN1062_sign_out(3);
    CN223_data_in(19) <= VN1136_data_out(3);
    CN223_sign_in(19) <= VN1136_sign_out(3);
    CN223_data_in(20) <= VN1169_data_out(3);
    CN223_sign_in(20) <= VN1169_sign_out(3);
    CN223_data_in(21) <= VN1207_data_out(3);
    CN223_sign_in(21) <= VN1207_sign_out(3);
    CN223_data_in(22) <= VN1264_data_out(3);
    CN223_sign_in(22) <= VN1264_sign_out(3);
    CN223_data_in(23) <= VN1325_data_out(3);
    CN223_sign_in(23) <= VN1325_sign_out(3);
    CN223_data_in(24) <= VN1336_data_out(3);
    CN223_sign_in(24) <= VN1336_sign_out(3);
    CN223_data_in(25) <= VN1406_data_out(3);
    CN223_sign_in(25) <= VN1406_sign_out(3);
    CN223_data_in(26) <= VN1474_data_out(3);
    CN223_sign_in(26) <= VN1474_sign_out(3);
    CN223_data_in(27) <= VN1577_data_out(3);
    CN223_sign_in(27) <= VN1577_sign_out(3);
    CN223_data_in(28) <= VN1620_data_out(3);
    CN223_sign_in(28) <= VN1620_sign_out(3);
    CN223_data_in(29) <= VN1659_data_out(3);
    CN223_sign_in(29) <= VN1659_sign_out(3);
    CN223_data_in(30) <= VN1714_data_out(3);
    CN223_sign_in(30) <= VN1714_sign_out(3);
    CN223_data_in(31) <= VN1779_data_out(3);
    CN223_sign_in(31) <= VN1779_sign_out(3);
    CN224_data_in(0) <= VN22_data_out(3);
    CN224_sign_in(0) <= VN22_sign_out(3);
    CN224_data_in(1) <= VN90_data_out(3);
    CN224_sign_in(1) <= VN90_sign_out(3);
    CN224_data_in(2) <= VN135_data_out(3);
    CN224_sign_in(2) <= VN135_sign_out(3);
    CN224_data_in(3) <= VN193_data_out(3);
    CN224_sign_in(3) <= VN193_sign_out(3);
    CN224_data_in(4) <= VN270_data_out(3);
    CN224_sign_in(4) <= VN270_sign_out(3);
    CN224_data_in(5) <= VN328_data_out(3);
    CN224_sign_in(5) <= VN328_sign_out(3);
    CN224_data_in(6) <= VN366_data_out(3);
    CN224_sign_in(6) <= VN366_sign_out(3);
    CN224_data_in(7) <= VN419_data_out(3);
    CN224_sign_in(7) <= VN419_sign_out(3);
    CN224_data_in(8) <= VN472_data_out(3);
    CN224_sign_in(8) <= VN472_sign_out(3);
    CN224_data_in(9) <= VN520_data_out(3);
    CN224_sign_in(9) <= VN520_sign_out(3);
    CN224_data_in(10) <= VN623_data_out(3);
    CN224_sign_in(10) <= VN623_sign_out(3);
    CN224_data_in(11) <= VN718_data_out(3);
    CN224_sign_in(11) <= VN718_sign_out(3);
    CN224_data_in(12) <= VN775_data_out(3);
    CN224_sign_in(12) <= VN775_sign_out(3);
    CN224_data_in(13) <= VN779_data_out(3);
    CN224_sign_in(13) <= VN779_sign_out(3);
    CN224_data_in(14) <= VN865_data_out(3);
    CN224_sign_in(14) <= VN865_sign_out(3);
    CN224_data_in(15) <= VN914_data_out(3);
    CN224_sign_in(15) <= VN914_sign_out(3);
    CN224_data_in(16) <= VN967_data_out(3);
    CN224_sign_in(16) <= VN967_sign_out(3);
    CN224_data_in(17) <= VN1022_data_out(3);
    CN224_sign_in(17) <= VN1022_sign_out(3);
    CN224_data_in(18) <= VN1066_data_out(3);
    CN224_sign_in(18) <= VN1066_sign_out(3);
    CN224_data_in(19) <= VN1112_data_out(3);
    CN224_sign_in(19) <= VN1112_sign_out(3);
    CN224_data_in(20) <= VN1174_data_out(3);
    CN224_sign_in(20) <= VN1174_sign_out(3);
    CN224_data_in(21) <= VN1228_data_out(3);
    CN224_sign_in(21) <= VN1228_sign_out(3);
    CN224_data_in(22) <= VN1284_data_out(3);
    CN224_sign_in(22) <= VN1284_sign_out(3);
    CN224_data_in(23) <= VN1373_data_out(3);
    CN224_sign_in(23) <= VN1373_sign_out(3);
    CN224_data_in(24) <= VN1411_data_out(3);
    CN224_sign_in(24) <= VN1411_sign_out(3);
    CN224_data_in(25) <= VN1442_data_out(3);
    CN224_sign_in(25) <= VN1442_sign_out(3);
    CN224_data_in(26) <= VN1480_data_out(3);
    CN224_sign_in(26) <= VN1480_sign_out(3);
    CN224_data_in(27) <= VN1511_data_out(3);
    CN224_sign_in(27) <= VN1511_sign_out(3);
    CN224_data_in(28) <= VN1615_data_out(3);
    CN224_sign_in(28) <= VN1615_sign_out(3);
    CN224_data_in(29) <= VN1655_data_out(3);
    CN224_sign_in(29) <= VN1655_sign_out(3);
    CN224_data_in(30) <= VN1708_data_out(3);
    CN224_sign_in(30) <= VN1708_sign_out(3);
    CN224_data_in(31) <= VN1780_data_out(3);
    CN224_sign_in(31) <= VN1780_sign_out(3);
    CN225_data_in(0) <= VN21_data_out(3);
    CN225_sign_in(0) <= VN21_sign_out(3);
    CN225_data_in(1) <= VN61_data_out(3);
    CN225_sign_in(1) <= VN61_sign_out(3);
    CN225_data_in(2) <= VN132_data_out(3);
    CN225_sign_in(2) <= VN132_sign_out(3);
    CN225_data_in(3) <= VN188_data_out(3);
    CN225_sign_in(3) <= VN188_sign_out(3);
    CN225_data_in(4) <= VN232_data_out(3);
    CN225_sign_in(4) <= VN232_sign_out(3);
    CN225_data_in(5) <= VN301_data_out(3);
    CN225_sign_in(5) <= VN301_sign_out(3);
    CN225_data_in(6) <= VN441_data_out(3);
    CN225_sign_in(6) <= VN441_sign_out(3);
    CN225_data_in(7) <= VN458_data_out(3);
    CN225_sign_in(7) <= VN458_sign_out(3);
    CN225_data_in(8) <= VN545_data_out(3);
    CN225_sign_in(8) <= VN545_sign_out(3);
    CN225_data_in(9) <= VN609_data_out(3);
    CN225_sign_in(9) <= VN609_sign_out(3);
    CN225_data_in(10) <= VN812_data_out(3);
    CN225_sign_in(10) <= VN812_sign_out(3);
    CN225_data_in(11) <= VN873_data_out(3);
    CN225_sign_in(11) <= VN873_sign_out(3);
    CN225_data_in(12) <= VN993_data_out(3);
    CN225_sign_in(12) <= VN993_sign_out(3);
    CN225_data_in(13) <= VN1029_data_out(3);
    CN225_sign_in(13) <= VN1029_sign_out(3);
    CN225_data_in(14) <= VN1143_data_out(3);
    CN225_sign_in(14) <= VN1143_sign_out(3);
    CN225_data_in(15) <= VN1248_data_out(3);
    CN225_sign_in(15) <= VN1248_sign_out(3);
    CN225_data_in(16) <= VN1486_data_out(3);
    CN225_sign_in(16) <= VN1486_sign_out(3);
    CN225_data_in(17) <= VN1506_data_out(3);
    CN225_sign_in(17) <= VN1506_sign_out(3);
    CN225_data_in(18) <= VN1526_data_out(3);
    CN225_sign_in(18) <= VN1526_sign_out(3);
    CN225_data_in(19) <= VN1533_data_out(3);
    CN225_sign_in(19) <= VN1533_sign_out(3);
    CN225_data_in(20) <= VN1552_data_out(3);
    CN225_sign_in(20) <= VN1552_sign_out(3);
    CN225_data_in(21) <= VN1564_data_out(3);
    CN225_sign_in(21) <= VN1564_sign_out(3);
    CN225_data_in(22) <= VN1621_data_out(3);
    CN225_sign_in(22) <= VN1621_sign_out(3);
    CN225_data_in(23) <= VN1682_data_out(3);
    CN225_sign_in(23) <= VN1682_sign_out(3);
    CN225_data_in(24) <= VN1739_data_out(3);
    CN225_sign_in(24) <= VN1739_sign_out(3);
    CN225_data_in(25) <= VN1800_data_out(3);
    CN225_sign_in(25) <= VN1800_sign_out(3);
    CN225_data_in(26) <= VN1873_data_out(3);
    CN225_sign_in(26) <= VN1873_sign_out(3);
    CN225_data_in(27) <= VN1874_data_out(3);
    CN225_sign_in(27) <= VN1874_sign_out(3);
    CN225_data_in(28) <= VN1925_data_out(3);
    CN225_sign_in(28) <= VN1925_sign_out(3);
    CN225_data_in(29) <= VN1948_data_out(3);
    CN225_sign_in(29) <= VN1948_sign_out(3);
    CN225_data_in(30) <= VN1958_data_out(3);
    CN225_sign_in(30) <= VN1958_sign_out(3);
    CN225_data_in(31) <= VN1965_data_out(3);
    CN225_sign_in(31) <= VN1965_sign_out(3);
    CN226_data_in(0) <= VN20_data_out(3);
    CN226_sign_in(0) <= VN20_sign_out(3);
    CN226_data_in(1) <= VN148_data_out(3);
    CN226_sign_in(1) <= VN148_sign_out(3);
    CN226_data_in(2) <= VN378_data_out(3);
    CN226_sign_in(2) <= VN378_sign_out(3);
    CN226_data_in(3) <= VN488_data_out(3);
    CN226_sign_in(3) <= VN488_sign_out(3);
    CN226_data_in(4) <= VN591_data_out(3);
    CN226_sign_in(4) <= VN591_sign_out(3);
    CN226_data_in(5) <= VN758_data_out(3);
    CN226_sign_in(5) <= VN758_sign_out(3);
    CN226_data_in(6) <= VN868_data_out(3);
    CN226_sign_in(6) <= VN868_sign_out(3);
    CN226_data_in(7) <= VN897_data_out(3);
    CN226_sign_in(7) <= VN897_sign_out(3);
    CN226_data_in(8) <= VN974_data_out(3);
    CN226_sign_in(8) <= VN974_sign_out(3);
    CN226_data_in(9) <= VN1005_data_out(3);
    CN226_sign_in(9) <= VN1005_sign_out(3);
    CN226_data_in(10) <= VN1206_data_out(3);
    CN226_sign_in(10) <= VN1206_sign_out(3);
    CN226_data_in(11) <= VN1249_data_out(3);
    CN226_sign_in(11) <= VN1249_sign_out(3);
    CN226_data_in(12) <= VN1337_data_out(3);
    CN226_sign_in(12) <= VN1337_sign_out(3);
    CN226_data_in(13) <= VN1410_data_out(3);
    CN226_sign_in(13) <= VN1410_sign_out(3);
    CN226_data_in(14) <= VN1451_data_out(3);
    CN226_sign_in(14) <= VN1451_sign_out(3);
    CN226_data_in(15) <= VN1466_data_out(3);
    CN226_sign_in(15) <= VN1466_sign_out(3);
    CN226_data_in(16) <= VN1530_data_out(3);
    CN226_sign_in(16) <= VN1530_sign_out(3);
    CN226_data_in(17) <= VN1569_data_out(3);
    CN226_sign_in(17) <= VN1569_sign_out(3);
    CN226_data_in(18) <= VN1611_data_out(3);
    CN226_sign_in(18) <= VN1611_sign_out(3);
    CN226_data_in(19) <= VN1649_data_out(3);
    CN226_sign_in(19) <= VN1649_sign_out(3);
    CN226_data_in(20) <= VN1688_data_out(3);
    CN226_sign_in(20) <= VN1688_sign_out(3);
    CN226_data_in(21) <= VN1825_data_out(3);
    CN226_sign_in(21) <= VN1825_sign_out(3);
    CN226_data_in(22) <= VN1943_data_out(3);
    CN226_sign_in(22) <= VN1943_sign_out(3);
    CN226_data_in(23) <= VN1964_data_out(3);
    CN226_sign_in(23) <= VN1964_sign_out(3);
    CN226_data_in(24) <= VN1970_data_out(3);
    CN226_sign_in(24) <= VN1970_sign_out(3);
    CN226_data_in(25) <= VN1990_data_out(3);
    CN226_sign_in(25) <= VN1990_sign_out(3);
    CN226_data_in(26) <= VN1993_data_out(3);
    CN226_sign_in(26) <= VN1993_sign_out(3);
    CN226_data_in(27) <= VN2003_data_out(3);
    CN226_sign_in(27) <= VN2003_sign_out(3);
    CN226_data_in(28) <= VN2017_data_out(3);
    CN226_sign_in(28) <= VN2017_sign_out(3);
    CN226_data_in(29) <= VN2026_data_out(3);
    CN226_sign_in(29) <= VN2026_sign_out(3);
    CN226_data_in(30) <= VN2034_data_out(3);
    CN226_sign_in(30) <= VN2034_sign_out(3);
    CN226_data_in(31) <= VN2045_data_out(3);
    CN226_sign_in(31) <= VN2045_sign_out(3);
    CN227_data_in(0) <= VN19_data_out(3);
    CN227_sign_in(0) <= VN19_sign_out(3);
    CN227_data_in(1) <= VN63_data_out(3);
    CN227_sign_in(1) <= VN63_sign_out(3);
    CN227_data_in(2) <= VN140_data_out(3);
    CN227_sign_in(2) <= VN140_sign_out(3);
    CN227_data_in(3) <= VN178_data_out(3);
    CN227_sign_in(3) <= VN178_sign_out(3);
    CN227_data_in(4) <= VN258_data_out(3);
    CN227_sign_in(4) <= VN258_sign_out(3);
    CN227_data_in(5) <= VN314_data_out(3);
    CN227_sign_in(5) <= VN314_sign_out(3);
    CN227_data_in(6) <= VN368_data_out(3);
    CN227_sign_in(6) <= VN368_sign_out(3);
    CN227_data_in(7) <= VN417_data_out(3);
    CN227_sign_in(7) <= VN417_sign_out(3);
    CN227_data_in(8) <= VN454_data_out(3);
    CN227_sign_in(8) <= VN454_sign_out(3);
    CN227_data_in(9) <= VN555_data_out(3);
    CN227_sign_in(9) <= VN555_sign_out(3);
    CN227_data_in(10) <= VN593_data_out(3);
    CN227_sign_in(10) <= VN593_sign_out(3);
    CN227_data_in(11) <= VN634_data_out(3);
    CN227_sign_in(11) <= VN634_sign_out(3);
    CN227_data_in(12) <= VN691_data_out(3);
    CN227_sign_in(12) <= VN691_sign_out(3);
    CN227_data_in(13) <= VN746_data_out(3);
    CN227_sign_in(13) <= VN746_sign_out(3);
    CN227_data_in(14) <= VN807_data_out(3);
    CN227_sign_in(14) <= VN807_sign_out(3);
    CN227_data_in(15) <= VN874_data_out(3);
    CN227_sign_in(15) <= VN874_sign_out(3);
    CN227_data_in(16) <= VN898_data_out(3);
    CN227_sign_in(16) <= VN898_sign_out(3);
    CN227_data_in(17) <= VN986_data_out(3);
    CN227_sign_in(17) <= VN986_sign_out(3);
    CN227_data_in(18) <= VN1018_data_out(3);
    CN227_sign_in(18) <= VN1018_sign_out(3);
    CN227_data_in(19) <= VN1075_data_out(3);
    CN227_sign_in(19) <= VN1075_sign_out(3);
    CN227_data_in(20) <= VN1123_data_out(3);
    CN227_sign_in(20) <= VN1123_sign_out(3);
    CN227_data_in(21) <= VN1198_data_out(3);
    CN227_sign_in(21) <= VN1198_sign_out(3);
    CN227_data_in(22) <= VN1227_data_out(3);
    CN227_sign_in(22) <= VN1227_sign_out(3);
    CN227_data_in(23) <= VN1322_data_out(3);
    CN227_sign_in(23) <= VN1322_sign_out(3);
    CN227_data_in(24) <= VN1366_data_out(3);
    CN227_sign_in(24) <= VN1366_sign_out(3);
    CN227_data_in(25) <= VN1404_data_out(3);
    CN227_sign_in(25) <= VN1404_sign_out(3);
    CN227_data_in(26) <= VN1445_data_out(3);
    CN227_sign_in(26) <= VN1445_sign_out(3);
    CN227_data_in(27) <= VN1575_data_out(3);
    CN227_sign_in(27) <= VN1575_sign_out(3);
    CN227_data_in(28) <= VN1595_data_out(3);
    CN227_sign_in(28) <= VN1595_sign_out(3);
    CN227_data_in(29) <= VN1631_data_out(3);
    CN227_sign_in(29) <= VN1631_sign_out(3);
    CN227_data_in(30) <= VN1706_data_out(3);
    CN227_sign_in(30) <= VN1706_sign_out(3);
    CN227_data_in(31) <= VN1781_data_out(3);
    CN227_sign_in(31) <= VN1781_sign_out(3);
    CN228_data_in(0) <= VN18_data_out(3);
    CN228_sign_in(0) <= VN18_sign_out(3);
    CN228_data_in(1) <= VN78_data_out(3);
    CN228_sign_in(1) <= VN78_sign_out(3);
    CN228_data_in(2) <= VN114_data_out(3);
    CN228_sign_in(2) <= VN114_sign_out(3);
    CN228_data_in(3) <= VN198_data_out(3);
    CN228_sign_in(3) <= VN198_sign_out(3);
    CN228_data_in(4) <= VN253_data_out(3);
    CN228_sign_in(4) <= VN253_sign_out(3);
    CN228_data_in(5) <= VN307_data_out(3);
    CN228_sign_in(5) <= VN307_sign_out(3);
    CN228_data_in(6) <= VN398_data_out(3);
    CN228_sign_in(6) <= VN398_sign_out(3);
    CN228_data_in(7) <= VN480_data_out(3);
    CN228_sign_in(7) <= VN480_sign_out(3);
    CN228_data_in(8) <= VN580_data_out(3);
    CN228_sign_in(8) <= VN580_sign_out(3);
    CN228_data_in(9) <= VN668_data_out(3);
    CN228_sign_in(9) <= VN668_sign_out(3);
    CN228_data_in(10) <= VN713_data_out(3);
    CN228_sign_in(10) <= VN713_sign_out(3);
    CN228_data_in(11) <= VN733_data_out(3);
    CN228_sign_in(11) <= VN733_sign_out(3);
    CN228_data_in(12) <= VN819_data_out(3);
    CN228_sign_in(12) <= VN819_sign_out(3);
    CN228_data_in(13) <= VN994_data_out(3);
    CN228_sign_in(13) <= VN994_sign_out(3);
    CN228_data_in(14) <= VN1046_data_out(3);
    CN228_sign_in(14) <= VN1046_sign_out(3);
    CN228_data_in(15) <= VN1086_data_out(3);
    CN228_sign_in(15) <= VN1086_sign_out(3);
    CN228_data_in(16) <= VN1120_data_out(3);
    CN228_sign_in(16) <= VN1120_sign_out(3);
    CN228_data_in(17) <= VN1275_data_out(3);
    CN228_sign_in(17) <= VN1275_sign_out(3);
    CN228_data_in(18) <= VN1303_data_out(3);
    CN228_sign_in(18) <= VN1303_sign_out(3);
    CN228_data_in(19) <= VN1380_data_out(3);
    CN228_sign_in(19) <= VN1380_sign_out(3);
    CN228_data_in(20) <= VN1449_data_out(3);
    CN228_sign_in(20) <= VN1449_sign_out(3);
    CN228_data_in(21) <= VN1549_data_out(3);
    CN228_sign_in(21) <= VN1549_sign_out(3);
    CN228_data_in(22) <= VN1568_data_out(3);
    CN228_sign_in(22) <= VN1568_sign_out(3);
    CN228_data_in(23) <= VN1583_data_out(3);
    CN228_sign_in(23) <= VN1583_sign_out(3);
    CN228_data_in(24) <= VN1697_data_out(3);
    CN228_sign_in(24) <= VN1697_sign_out(3);
    CN228_data_in(25) <= VN1863_data_out(3);
    CN228_sign_in(25) <= VN1863_sign_out(3);
    CN228_data_in(26) <= VN1937_data_out(3);
    CN228_sign_in(26) <= VN1937_sign_out(3);
    CN228_data_in(27) <= VN1942_data_out(3);
    CN228_sign_in(27) <= VN1942_sign_out(3);
    CN228_data_in(28) <= VN1962_data_out(3);
    CN228_sign_in(28) <= VN1962_sign_out(3);
    CN228_data_in(29) <= VN1972_data_out(3);
    CN228_sign_in(29) <= VN1972_sign_out(3);
    CN228_data_in(30) <= VN1998_data_out(3);
    CN228_sign_in(30) <= VN1998_sign_out(3);
    CN228_data_in(31) <= VN2004_data_out(3);
    CN228_sign_in(31) <= VN2004_sign_out(3);
    CN229_data_in(0) <= VN17_data_out(3);
    CN229_sign_in(0) <= VN17_sign_out(3);
    CN229_data_in(1) <= VN74_data_out(3);
    CN229_sign_in(1) <= VN74_sign_out(3);
    CN229_data_in(2) <= VN124_data_out(3);
    CN229_sign_in(2) <= VN124_sign_out(3);
    CN229_data_in(3) <= VN259_data_out(3);
    CN229_sign_in(3) <= VN259_sign_out(3);
    CN229_data_in(4) <= VN374_data_out(3);
    CN229_sign_in(4) <= VN374_sign_out(3);
    CN229_data_in(5) <= VN466_data_out(3);
    CN229_sign_in(5) <= VN466_sign_out(3);
    CN229_data_in(6) <= VN538_data_out(3);
    CN229_sign_in(6) <= VN538_sign_out(3);
    CN229_data_in(7) <= VN610_data_out(3);
    CN229_sign_in(7) <= VN610_sign_out(3);
    CN229_data_in(8) <= VN633_data_out(3);
    CN229_sign_in(8) <= VN633_sign_out(3);
    CN229_data_in(9) <= VN832_data_out(3);
    CN229_sign_in(9) <= VN832_sign_out(3);
    CN229_data_in(10) <= VN923_data_out(3);
    CN229_sign_in(10) <= VN923_sign_out(3);
    CN229_data_in(11) <= VN966_data_out(3);
    CN229_sign_in(11) <= VN966_sign_out(3);
    CN229_data_in(12) <= VN1236_data_out(3);
    CN229_sign_in(12) <= VN1236_sign_out(3);
    CN229_data_in(13) <= VN1288_data_out(3);
    CN229_sign_in(13) <= VN1288_sign_out(3);
    CN229_data_in(14) <= VN1354_data_out(3);
    CN229_sign_in(14) <= VN1354_sign_out(3);
    CN229_data_in(15) <= VN1495_data_out(3);
    CN229_sign_in(15) <= VN1495_sign_out(3);
    CN229_data_in(16) <= VN1515_data_out(3);
    CN229_sign_in(16) <= VN1515_sign_out(3);
    CN229_data_in(17) <= VN1556_data_out(3);
    CN229_sign_in(17) <= VN1556_sign_out(3);
    CN229_data_in(18) <= VN1625_data_out(3);
    CN229_sign_in(18) <= VN1625_sign_out(3);
    CN229_data_in(19) <= VN1798_data_out(3);
    CN229_sign_in(19) <= VN1798_sign_out(3);
    CN229_data_in(20) <= VN1842_data_out(3);
    CN229_sign_in(20) <= VN1842_sign_out(3);
    CN229_data_in(21) <= VN1878_data_out(3);
    CN229_sign_in(21) <= VN1878_sign_out(3);
    CN229_data_in(22) <= VN1959_data_out(3);
    CN229_sign_in(22) <= VN1959_sign_out(3);
    CN229_data_in(23) <= VN1976_data_out(3);
    CN229_sign_in(23) <= VN1976_sign_out(3);
    CN229_data_in(24) <= VN1981_data_out(3);
    CN229_sign_in(24) <= VN1981_sign_out(3);
    CN229_data_in(25) <= VN1988_data_out(3);
    CN229_sign_in(25) <= VN1988_sign_out(3);
    CN229_data_in(26) <= VN1991_data_out(3);
    CN229_sign_in(26) <= VN1991_sign_out(3);
    CN229_data_in(27) <= VN2001_data_out(3);
    CN229_sign_in(27) <= VN2001_sign_out(3);
    CN229_data_in(28) <= VN2010_data_out(3);
    CN229_sign_in(28) <= VN2010_sign_out(3);
    CN229_data_in(29) <= VN2019_data_out(3);
    CN229_sign_in(29) <= VN2019_sign_out(3);
    CN229_data_in(30) <= VN2031_data_out(3);
    CN229_sign_in(30) <= VN2031_sign_out(3);
    CN229_data_in(31) <= VN2043_data_out(3);
    CN229_sign_in(31) <= VN2043_sign_out(3);
    CN230_data_in(0) <= VN16_data_out(3);
    CN230_sign_in(0) <= VN16_sign_out(3);
    CN230_data_in(1) <= VN118_data_out(3);
    CN230_sign_in(1) <= VN118_sign_out(3);
    CN230_data_in(2) <= VN176_data_out(3);
    CN230_sign_in(2) <= VN176_sign_out(3);
    CN230_data_in(3) <= VN249_data_out(3);
    CN230_sign_in(3) <= VN249_sign_out(3);
    CN230_data_in(4) <= VN293_data_out(3);
    CN230_sign_in(4) <= VN293_sign_out(3);
    CN230_data_in(5) <= VN347_data_out(3);
    CN230_sign_in(5) <= VN347_sign_out(3);
    CN230_data_in(6) <= VN442_data_out(3);
    CN230_sign_in(6) <= VN442_sign_out(3);
    CN230_data_in(7) <= VN490_data_out(3);
    CN230_sign_in(7) <= VN490_sign_out(3);
    CN230_data_in(8) <= VN539_data_out(3);
    CN230_sign_in(8) <= VN539_sign_out(3);
    CN230_data_in(9) <= VN577_data_out(3);
    CN230_sign_in(9) <= VN577_sign_out(3);
    CN230_data_in(10) <= VN690_data_out(3);
    CN230_sign_in(10) <= VN690_sign_out(3);
    CN230_data_in(11) <= VN780_data_out(3);
    CN230_sign_in(11) <= VN780_sign_out(3);
    CN230_data_in(12) <= VN838_data_out(3);
    CN230_sign_in(12) <= VN838_sign_out(3);
    CN230_data_in(13) <= VN939_data_out(3);
    CN230_sign_in(13) <= VN939_sign_out(3);
    CN230_data_in(14) <= VN981_data_out(3);
    CN230_sign_in(14) <= VN981_sign_out(3);
    CN230_data_in(15) <= VN1048_data_out(3);
    CN230_sign_in(15) <= VN1048_sign_out(3);
    CN230_data_in(16) <= VN1069_data_out(3);
    CN230_sign_in(16) <= VN1069_sign_out(3);
    CN230_data_in(17) <= VN1161_data_out(3);
    CN230_sign_in(17) <= VN1161_sign_out(3);
    CN230_data_in(18) <= VN1218_data_out(3);
    CN230_sign_in(18) <= VN1218_sign_out(3);
    CN230_data_in(19) <= VN1240_data_out(3);
    CN230_sign_in(19) <= VN1240_sign_out(3);
    CN230_data_in(20) <= VN1300_data_out(3);
    CN230_sign_in(20) <= VN1300_sign_out(3);
    CN230_data_in(21) <= VN1519_data_out(3);
    CN230_sign_in(21) <= VN1519_sign_out(3);
    CN230_data_in(22) <= VN1600_data_out(3);
    CN230_sign_in(22) <= VN1600_sign_out(3);
    CN230_data_in(23) <= VN1626_data_out(3);
    CN230_sign_in(23) <= VN1626_sign_out(3);
    CN230_data_in(24) <= VN1700_data_out(3);
    CN230_sign_in(24) <= VN1700_sign_out(3);
    CN230_data_in(25) <= VN1809_data_out(3);
    CN230_sign_in(25) <= VN1809_sign_out(3);
    CN230_data_in(26) <= VN1819_data_out(3);
    CN230_sign_in(26) <= VN1819_sign_out(3);
    CN230_data_in(27) <= VN1831_data_out(3);
    CN230_sign_in(27) <= VN1831_sign_out(3);
    CN230_data_in(28) <= VN1949_data_out(3);
    CN230_sign_in(28) <= VN1949_sign_out(3);
    CN230_data_in(29) <= VN1978_data_out(3);
    CN230_sign_in(29) <= VN1978_sign_out(3);
    CN230_data_in(30) <= VN1996_data_out(3);
    CN230_sign_in(30) <= VN1996_sign_out(3);
    CN230_data_in(31) <= VN2005_data_out(3);
    CN230_sign_in(31) <= VN2005_sign_out(3);
    CN231_data_in(0) <= VN15_data_out(3);
    CN231_sign_in(0) <= VN15_sign_out(3);
    CN231_data_in(1) <= VN56_data_out(3);
    CN231_sign_in(1) <= VN56_sign_out(3);
    CN231_data_in(2) <= VN209_data_out(3);
    CN231_sign_in(2) <= VN209_sign_out(3);
    CN231_data_in(3) <= VN272_data_out(3);
    CN231_sign_in(3) <= VN272_sign_out(3);
    CN231_data_in(4) <= VN287_data_out(3);
    CN231_sign_in(4) <= VN287_sign_out(3);
    CN231_data_in(5) <= VN344_data_out(3);
    CN231_sign_in(5) <= VN344_sign_out(3);
    CN231_data_in(6) <= VN418_data_out(3);
    CN231_sign_in(6) <= VN418_sign_out(3);
    CN231_data_in(7) <= VN482_data_out(3);
    CN231_sign_in(7) <= VN482_sign_out(3);
    CN231_data_in(8) <= VN516_data_out(3);
    CN231_sign_in(8) <= VN516_sign_out(3);
    CN231_data_in(9) <= VN602_data_out(3);
    CN231_sign_in(9) <= VN602_sign_out(3);
    CN231_data_in(10) <= VN666_data_out(3);
    CN231_sign_in(10) <= VN666_sign_out(3);
    CN231_data_in(11) <= VN682_data_out(3);
    CN231_sign_in(11) <= VN682_sign_out(3);
    CN231_data_in(12) <= VN722_data_out(3);
    CN231_sign_in(12) <= VN722_sign_out(3);
    CN231_data_in(13) <= VN776_data_out(3);
    CN231_sign_in(13) <= VN776_sign_out(3);
    CN231_data_in(14) <= VN821_data_out(3);
    CN231_sign_in(14) <= VN821_sign_out(3);
    CN231_data_in(15) <= VN877_data_out(3);
    CN231_sign_in(15) <= VN877_sign_out(3);
    CN231_data_in(16) <= VN943_data_out(3);
    CN231_sign_in(16) <= VN943_sign_out(3);
    CN231_data_in(17) <= VN952_data_out(3);
    CN231_sign_in(17) <= VN952_sign_out(3);
    CN231_data_in(18) <= VN1006_data_out(3);
    CN231_sign_in(18) <= VN1006_sign_out(3);
    CN231_data_in(19) <= VN1162_data_out(3);
    CN231_sign_in(19) <= VN1162_sign_out(3);
    CN231_data_in(20) <= VN1217_data_out(3);
    CN231_sign_in(20) <= VN1217_sign_out(3);
    CN231_data_in(21) <= VN1308_data_out(3);
    CN231_sign_in(21) <= VN1308_sign_out(3);
    CN231_data_in(22) <= VN1355_data_out(3);
    CN231_sign_in(22) <= VN1355_sign_out(3);
    CN231_data_in(23) <= VN1414_data_out(3);
    CN231_sign_in(23) <= VN1414_sign_out(3);
    CN231_data_in(24) <= VN1470_data_out(3);
    CN231_sign_in(24) <= VN1470_sign_out(3);
    CN231_data_in(25) <= VN1507_data_out(3);
    CN231_sign_in(25) <= VN1507_sign_out(3);
    CN231_data_in(26) <= VN1525_data_out(3);
    CN231_sign_in(26) <= VN1525_sign_out(3);
    CN231_data_in(27) <= VN1578_data_out(3);
    CN231_sign_in(27) <= VN1578_sign_out(3);
    CN231_data_in(28) <= VN1647_data_out(3);
    CN231_sign_in(28) <= VN1647_sign_out(3);
    CN231_data_in(29) <= VN1672_data_out(3);
    CN231_sign_in(29) <= VN1672_sign_out(3);
    CN231_data_in(30) <= VN1804_data_out(3);
    CN231_sign_in(30) <= VN1804_sign_out(3);
    CN231_data_in(31) <= VN1852_data_out(3);
    CN231_sign_in(31) <= VN1852_sign_out(3);
    CN232_data_in(0) <= VN14_data_out(3);
    CN232_sign_in(0) <= VN14_sign_out(3);
    CN232_data_in(1) <= VN57_data_out(3);
    CN232_sign_in(1) <= VN57_sign_out(3);
    CN232_data_in(2) <= VN212_data_out(3);
    CN232_sign_in(2) <= VN212_sign_out(3);
    CN232_data_in(3) <= VN278_data_out(3);
    CN232_sign_in(3) <= VN278_sign_out(3);
    CN232_data_in(4) <= VN291_data_out(3);
    CN232_sign_in(4) <= VN291_sign_out(3);
    CN232_data_in(5) <= VN359_data_out(3);
    CN232_sign_in(5) <= VN359_sign_out(3);
    CN232_data_in(6) <= VN439_data_out(3);
    CN232_sign_in(6) <= VN439_sign_out(3);
    CN232_data_in(7) <= VN470_data_out(3);
    CN232_sign_in(7) <= VN470_sign_out(3);
    CN232_data_in(8) <= VN509_data_out(3);
    CN232_sign_in(8) <= VN509_sign_out(3);
    CN232_data_in(9) <= VN700_data_out(3);
    CN232_sign_in(9) <= VN700_sign_out(3);
    CN232_data_in(10) <= VN783_data_out(3);
    CN232_sign_in(10) <= VN783_sign_out(3);
    CN232_data_in(11) <= VN879_data_out(3);
    CN232_sign_in(11) <= VN879_sign_out(3);
    CN232_data_in(12) <= VN989_data_out(3);
    CN232_sign_in(12) <= VN989_sign_out(3);
    CN232_data_in(13) <= VN1097_data_out(3);
    CN232_sign_in(13) <= VN1097_sign_out(3);
    CN232_data_in(14) <= VN1138_data_out(3);
    CN232_sign_in(14) <= VN1138_sign_out(3);
    CN232_data_in(15) <= VN1166_data_out(3);
    CN232_sign_in(15) <= VN1166_sign_out(3);
    CN232_data_in(16) <= VN1213_data_out(3);
    CN232_sign_in(16) <= VN1213_sign_out(3);
    CN232_data_in(17) <= VN1368_data_out(3);
    CN232_sign_in(17) <= VN1368_sign_out(3);
    CN232_data_in(18) <= VN1476_data_out(3);
    CN232_sign_in(18) <= VN1476_sign_out(3);
    CN232_data_in(19) <= VN1502_data_out(3);
    CN232_sign_in(19) <= VN1502_sign_out(3);
    CN232_data_in(20) <= VN1504_data_out(3);
    CN232_sign_in(20) <= VN1504_sign_out(3);
    CN232_data_in(21) <= VN1573_data_out(3);
    CN232_sign_in(21) <= VN1573_sign_out(3);
    CN232_data_in(22) <= VN1664_data_out(3);
    CN232_sign_in(22) <= VN1664_sign_out(3);
    CN232_data_in(23) <= VN1746_data_out(3);
    CN232_sign_in(23) <= VN1746_sign_out(3);
    CN232_data_in(24) <= VN1756_data_out(3);
    CN232_sign_in(24) <= VN1756_sign_out(3);
    CN232_data_in(25) <= VN1760_data_out(3);
    CN232_sign_in(25) <= VN1760_sign_out(3);
    CN232_data_in(26) <= VN1864_data_out(3);
    CN232_sign_in(26) <= VN1864_sign_out(3);
    CN232_data_in(27) <= VN1910_data_out(3);
    CN232_sign_in(27) <= VN1910_sign_out(3);
    CN232_data_in(28) <= VN1920_data_out(3);
    CN232_sign_in(28) <= VN1920_sign_out(3);
    CN232_data_in(29) <= VN1951_data_out(3);
    CN232_sign_in(29) <= VN1951_sign_out(3);
    CN232_data_in(30) <= VN1952_data_out(3);
    CN232_sign_in(30) <= VN1952_sign_out(3);
    CN232_data_in(31) <= VN1966_data_out(3);
    CN232_sign_in(31) <= VN1966_sign_out(3);
    CN233_data_in(0) <= VN13_data_out(3);
    CN233_sign_in(0) <= VN13_sign_out(3);
    CN233_data_in(1) <= VN92_data_out(3);
    CN233_sign_in(1) <= VN92_sign_out(3);
    CN233_data_in(2) <= VN149_data_out(3);
    CN233_sign_in(2) <= VN149_sign_out(3);
    CN233_data_in(3) <= VN263_data_out(3);
    CN233_sign_in(3) <= VN263_sign_out(3);
    CN233_data_in(4) <= VN352_data_out(3);
    CN233_sign_in(4) <= VN352_sign_out(3);
    CN233_data_in(5) <= VN486_data_out(3);
    CN233_sign_in(5) <= VN486_sign_out(3);
    CN233_data_in(6) <= VN612_data_out(3);
    CN233_sign_in(6) <= VN612_sign_out(3);
    CN233_data_in(7) <= VN640_data_out(3);
    CN233_sign_in(7) <= VN640_sign_out(3);
    CN233_data_in(8) <= VN723_data_out(3);
    CN233_sign_in(8) <= VN723_sign_out(3);
    CN233_data_in(9) <= VN850_data_out(3);
    CN233_sign_in(9) <= VN850_sign_out(3);
    CN233_data_in(10) <= VN954_data_out(3);
    CN233_sign_in(10) <= VN954_sign_out(3);
    CN233_data_in(11) <= VN1195_data_out(3);
    CN233_sign_in(11) <= VN1195_sign_out(3);
    CN233_data_in(12) <= VN1276_data_out(3);
    CN233_sign_in(12) <= VN1276_sign_out(3);
    CN233_data_in(13) <= VN1324_data_out(3);
    CN233_sign_in(13) <= VN1324_sign_out(3);
    CN233_data_in(14) <= VN1364_data_out(3);
    CN233_sign_in(14) <= VN1364_sign_out(3);
    CN233_data_in(15) <= VN1494_data_out(3);
    CN233_sign_in(15) <= VN1494_sign_out(3);
    CN233_data_in(16) <= VN1537_data_out(3);
    CN233_sign_in(16) <= VN1537_sign_out(3);
    CN233_data_in(17) <= VN1640_data_out(3);
    CN233_sign_in(17) <= VN1640_sign_out(3);
    CN233_data_in(18) <= VN1711_data_out(3);
    CN233_sign_in(18) <= VN1711_sign_out(3);
    CN233_data_in(19) <= VN1832_data_out(3);
    CN233_sign_in(19) <= VN1832_sign_out(3);
    CN233_data_in(20) <= VN1834_data_out(3);
    CN233_sign_in(20) <= VN1834_sign_out(3);
    CN233_data_in(21) <= VN1892_data_out(3);
    CN233_sign_in(21) <= VN1892_sign_out(3);
    CN233_data_in(22) <= VN1909_data_out(3);
    CN233_sign_in(22) <= VN1909_sign_out(3);
    CN233_data_in(23) <= VN1960_data_out(3);
    CN233_sign_in(23) <= VN1960_sign_out(3);
    CN233_data_in(24) <= VN1983_data_out(3);
    CN233_sign_in(24) <= VN1983_sign_out(3);
    CN233_data_in(25) <= VN1995_data_out(3);
    CN233_sign_in(25) <= VN1995_sign_out(3);
    CN233_data_in(26) <= VN2008_data_out(3);
    CN233_sign_in(26) <= VN2008_sign_out(3);
    CN233_data_in(27) <= VN2013_data_out(3);
    CN233_sign_in(27) <= VN2013_sign_out(3);
    CN233_data_in(28) <= VN2020_data_out(3);
    CN233_sign_in(28) <= VN2020_sign_out(3);
    CN233_data_in(29) <= VN2028_data_out(3);
    CN233_sign_in(29) <= VN2028_sign_out(3);
    CN233_data_in(30) <= VN2039_data_out(3);
    CN233_sign_in(30) <= VN2039_sign_out(3);
    CN233_data_in(31) <= VN2047_data_out(3);
    CN233_sign_in(31) <= VN2047_sign_out(3);
    CN234_data_in(0) <= VN12_data_out(3);
    CN234_sign_in(0) <= VN12_sign_out(3);
    CN234_data_in(1) <= VN84_data_out(3);
    CN234_sign_in(1) <= VN84_sign_out(3);
    CN234_data_in(2) <= VN131_data_out(3);
    CN234_sign_in(2) <= VN131_sign_out(3);
    CN234_data_in(3) <= VN177_data_out(3);
    CN234_sign_in(3) <= VN177_sign_out(3);
    CN234_data_in(4) <= VN265_data_out(3);
    CN234_sign_in(4) <= VN265_sign_out(3);
    CN234_data_in(5) <= VN315_data_out(3);
    CN234_sign_in(5) <= VN315_sign_out(3);
    CN234_data_in(6) <= VN386_data_out(3);
    CN234_sign_in(6) <= VN386_sign_out(3);
    CN234_data_in(7) <= VN394_data_out(3);
    CN234_sign_in(7) <= VN394_sign_out(3);
    CN234_data_in(8) <= VN463_data_out(3);
    CN234_sign_in(8) <= VN463_sign_out(3);
    CN234_data_in(9) <= VN528_data_out(3);
    CN234_sign_in(9) <= VN528_sign_out(3);
    CN234_data_in(10) <= VN603_data_out(3);
    CN234_sign_in(10) <= VN603_sign_out(3);
    CN234_data_in(11) <= VN638_data_out(3);
    CN234_sign_in(11) <= VN638_sign_out(3);
    CN234_data_in(12) <= VN768_data_out(3);
    CN234_sign_in(12) <= VN768_sign_out(3);
    CN234_data_in(13) <= VN809_data_out(3);
    CN234_sign_in(13) <= VN809_sign_out(3);
    CN234_data_in(14) <= VN886_data_out(3);
    CN234_sign_in(14) <= VN886_sign_out(3);
    CN234_data_in(15) <= VN937_data_out(3);
    CN234_sign_in(15) <= VN937_sign_out(3);
    CN234_data_in(16) <= VN968_data_out(3);
    CN234_sign_in(16) <= VN968_sign_out(3);
    CN234_data_in(17) <= VN1041_data_out(3);
    CN234_sign_in(17) <= VN1041_sign_out(3);
    CN234_data_in(18) <= VN1147_data_out(3);
    CN234_sign_in(18) <= VN1147_sign_out(3);
    CN234_data_in(19) <= VN1202_data_out(3);
    CN234_sign_in(19) <= VN1202_sign_out(3);
    CN234_data_in(20) <= VN1272_data_out(3);
    CN234_sign_in(20) <= VN1272_sign_out(3);
    CN234_data_in(21) <= VN1310_data_out(3);
    CN234_sign_in(21) <= VN1310_sign_out(3);
    CN234_data_in(22) <= VN1383_data_out(3);
    CN234_sign_in(22) <= VN1383_sign_out(3);
    CN234_data_in(23) <= VN1452_data_out(3);
    CN234_sign_in(23) <= VN1452_sign_out(3);
    CN234_data_in(24) <= VN1468_data_out(3);
    CN234_sign_in(24) <= VN1468_sign_out(3);
    CN234_data_in(25) <= VN1478_data_out(3);
    CN234_sign_in(25) <= VN1478_sign_out(3);
    CN234_data_in(26) <= VN1498_data_out(3);
    CN234_sign_in(26) <= VN1498_sign_out(3);
    CN234_data_in(27) <= VN1662_data_out(3);
    CN234_sign_in(27) <= VN1662_sign_out(3);
    CN234_data_in(28) <= VN1753_data_out(3);
    CN234_sign_in(28) <= VN1753_sign_out(3);
    CN234_data_in(29) <= VN1791_data_out(3);
    CN234_sign_in(29) <= VN1791_sign_out(3);
    CN234_data_in(30) <= VN1808_data_out(3);
    CN234_sign_in(30) <= VN1808_sign_out(3);
    CN234_data_in(31) <= VN1853_data_out(3);
    CN234_sign_in(31) <= VN1853_sign_out(3);
    CN235_data_in(0) <= VN100_data_out(3);
    CN235_sign_in(0) <= VN100_sign_out(3);
    CN235_data_in(1) <= VN144_data_out(3);
    CN235_sign_in(1) <= VN144_sign_out(3);
    CN235_data_in(2) <= VN196_data_out(3);
    CN235_sign_in(2) <= VN196_sign_out(3);
    CN235_data_in(3) <= VN235_data_out(3);
    CN235_sign_in(3) <= VN235_sign_out(3);
    CN235_data_in(4) <= VN336_data_out(3);
    CN235_sign_in(4) <= VN336_sign_out(3);
    CN235_data_in(5) <= VN420_data_out(3);
    CN235_sign_in(5) <= VN420_sign_out(3);
    CN235_data_in(6) <= VN460_data_out(3);
    CN235_sign_in(6) <= VN460_sign_out(3);
    CN235_data_in(7) <= VN619_data_out(3);
    CN235_sign_in(7) <= VN619_sign_out(3);
    CN235_data_in(8) <= VN704_data_out(3);
    CN235_sign_in(8) <= VN704_sign_out(3);
    CN235_data_in(9) <= VN736_data_out(3);
    CN235_sign_in(9) <= VN736_sign_out(3);
    CN235_data_in(10) <= VN805_data_out(3);
    CN235_sign_in(10) <= VN805_sign_out(3);
    CN235_data_in(11) <= VN842_data_out(3);
    CN235_sign_in(11) <= VN842_sign_out(3);
    CN235_data_in(12) <= VN921_data_out(3);
    CN235_sign_in(12) <= VN921_sign_out(3);
    CN235_data_in(13) <= VN964_data_out(3);
    CN235_sign_in(13) <= VN964_sign_out(3);
    CN235_data_in(14) <= VN1042_data_out(3);
    CN235_sign_in(14) <= VN1042_sign_out(3);
    CN235_data_in(15) <= VN1152_data_out(3);
    CN235_sign_in(15) <= VN1152_sign_out(3);
    CN235_data_in(16) <= VN1170_data_out(3);
    CN235_sign_in(16) <= VN1170_sign_out(3);
    CN235_data_in(17) <= VN1327_data_out(3);
    CN235_sign_in(17) <= VN1327_sign_out(3);
    CN235_data_in(18) <= VN1349_data_out(3);
    CN235_sign_in(18) <= VN1349_sign_out(3);
    CN235_data_in(19) <= VN1416_data_out(3);
    CN235_sign_in(19) <= VN1416_sign_out(3);
    CN235_data_in(20) <= VN1427_data_out(3);
    CN235_sign_in(20) <= VN1427_sign_out(3);
    CN235_data_in(21) <= VN1497_data_out(3);
    CN235_sign_in(21) <= VN1497_sign_out(3);
    CN235_data_in(22) <= VN1523_data_out(3);
    CN235_sign_in(22) <= VN1523_sign_out(3);
    CN235_data_in(23) <= VN1558_data_out(3);
    CN235_sign_in(23) <= VN1558_sign_out(3);
    CN235_data_in(24) <= VN1799_data_out(3);
    CN235_sign_in(24) <= VN1799_sign_out(3);
    CN235_data_in(25) <= VN1818_data_out(3);
    CN235_sign_in(25) <= VN1818_sign_out(3);
    CN235_data_in(26) <= VN1826_data_out(3);
    CN235_sign_in(26) <= VN1826_sign_out(3);
    CN235_data_in(27) <= VN1830_data_out(3);
    CN235_sign_in(27) <= VN1830_sign_out(3);
    CN235_data_in(28) <= VN1837_data_out(3);
    CN235_sign_in(28) <= VN1837_sign_out(3);
    CN235_data_in(29) <= VN1838_data_out(3);
    CN235_sign_in(29) <= VN1838_sign_out(3);
    CN235_data_in(30) <= VN1867_data_out(3);
    CN235_sign_in(30) <= VN1867_sign_out(3);
    CN235_data_in(31) <= VN1889_data_out(3);
    CN235_sign_in(31) <= VN1889_sign_out(3);
    CN236_data_in(0) <= VN11_data_out(3);
    CN236_sign_in(0) <= VN11_sign_out(3);
    CN236_data_in(1) <= VN104_data_out(3);
    CN236_sign_in(1) <= VN104_sign_out(3);
    CN236_data_in(2) <= VN155_data_out(3);
    CN236_sign_in(2) <= VN155_sign_out(3);
    CN236_data_in(3) <= VN221_data_out(3);
    CN236_sign_in(3) <= VN221_sign_out(3);
    CN236_data_in(4) <= VN271_data_out(3);
    CN236_sign_in(4) <= VN271_sign_out(3);
    CN236_data_in(5) <= VN310_data_out(3);
    CN236_sign_in(5) <= VN310_sign_out(3);
    CN236_data_in(6) <= VN390_data_out(3);
    CN236_sign_in(6) <= VN390_sign_out(3);
    CN236_data_in(7) <= VN410_data_out(3);
    CN236_sign_in(7) <= VN410_sign_out(3);
    CN236_data_in(8) <= VN475_data_out(3);
    CN236_sign_in(8) <= VN475_sign_out(3);
    CN236_data_in(9) <= VN527_data_out(3);
    CN236_sign_in(9) <= VN527_sign_out(3);
    CN236_data_in(10) <= VN608_data_out(3);
    CN236_sign_in(10) <= VN608_sign_out(3);
    CN236_data_in(11) <= VN653_data_out(3);
    CN236_sign_in(11) <= VN653_sign_out(3);
    CN236_data_in(12) <= VN698_data_out(3);
    CN236_sign_in(12) <= VN698_sign_out(3);
    CN236_data_in(13) <= VN742_data_out(3);
    CN236_sign_in(13) <= VN742_sign_out(3);
    CN236_data_in(14) <= VN810_data_out(3);
    CN236_sign_in(14) <= VN810_sign_out(3);
    CN236_data_in(15) <= VN851_data_out(3);
    CN236_sign_in(15) <= VN851_sign_out(3);
    CN236_data_in(16) <= VN927_data_out(3);
    CN236_sign_in(16) <= VN927_sign_out(3);
    CN236_data_in(17) <= VN984_data_out(3);
    CN236_sign_in(17) <= VN984_sign_out(3);
    CN236_data_in(18) <= VN1020_data_out(3);
    CN236_sign_in(18) <= VN1020_sign_out(3);
    CN236_data_in(19) <= VN1083_data_out(3);
    CN236_sign_in(19) <= VN1083_sign_out(3);
    CN236_data_in(20) <= VN1244_data_out(3);
    CN236_sign_in(20) <= VN1244_sign_out(3);
    CN236_data_in(21) <= VN1278_data_out(3);
    CN236_sign_in(21) <= VN1278_sign_out(3);
    CN236_data_in(22) <= VN1293_data_out(3);
    CN236_sign_in(22) <= VN1293_sign_out(3);
    CN236_data_in(23) <= VN1350_data_out(3);
    CN236_sign_in(23) <= VN1350_sign_out(3);
    CN236_data_in(24) <= VN1393_data_out(3);
    CN236_sign_in(24) <= VN1393_sign_out(3);
    CN236_data_in(25) <= VN1429_data_out(3);
    CN236_sign_in(25) <= VN1429_sign_out(3);
    CN236_data_in(26) <= VN1514_data_out(3);
    CN236_sign_in(26) <= VN1514_sign_out(3);
    CN236_data_in(27) <= VN1517_data_out(3);
    CN236_sign_in(27) <= VN1517_sign_out(3);
    CN236_data_in(28) <= VN1592_data_out(3);
    CN236_sign_in(28) <= VN1592_sign_out(3);
    CN236_data_in(29) <= VN1636_data_out(3);
    CN236_sign_in(29) <= VN1636_sign_out(3);
    CN236_data_in(30) <= VN1669_data_out(3);
    CN236_sign_in(30) <= VN1669_sign_out(3);
    CN236_data_in(31) <= VN1782_data_out(3);
    CN236_sign_in(31) <= VN1782_sign_out(3);
    CN237_data_in(0) <= VN10_data_out(3);
    CN237_sign_in(0) <= VN10_sign_out(3);
    CN237_data_in(1) <= VN110_data_out(3);
    CN237_sign_in(1) <= VN110_sign_out(3);
    CN237_data_in(2) <= VN125_data_out(3);
    CN237_sign_in(2) <= VN125_sign_out(3);
    CN237_data_in(3) <= VN228_data_out(3);
    CN237_sign_in(3) <= VN228_sign_out(3);
    CN237_data_in(4) <= VN322_data_out(3);
    CN237_sign_in(4) <= VN322_sign_out(3);
    CN237_data_in(5) <= VN334_data_out(3);
    CN237_sign_in(5) <= VN334_sign_out(3);
    CN237_data_in(6) <= VN399_data_out(3);
    CN237_sign_in(6) <= VN399_sign_out(3);
    CN237_data_in(7) <= VN467_data_out(3);
    CN237_sign_in(7) <= VN467_sign_out(3);
    CN237_data_in(8) <= VN522_data_out(3);
    CN237_sign_in(8) <= VN522_sign_out(3);
    CN237_data_in(9) <= VN584_data_out(3);
    CN237_sign_in(9) <= VN584_sign_out(3);
    CN237_data_in(10) <= VN654_data_out(3);
    CN237_sign_in(10) <= VN654_sign_out(3);
    CN237_data_in(11) <= VN680_data_out(3);
    CN237_sign_in(11) <= VN680_sign_out(3);
    CN237_data_in(12) <= VN726_data_out(3);
    CN237_sign_in(12) <= VN726_sign_out(3);
    CN237_data_in(13) <= VN800_data_out(3);
    CN237_sign_in(13) <= VN800_sign_out(3);
    CN237_data_in(14) <= VN878_data_out(3);
    CN237_sign_in(14) <= VN878_sign_out(3);
    CN237_data_in(15) <= VN893_data_out(3);
    CN237_sign_in(15) <= VN893_sign_out(3);
    CN237_data_in(16) <= VN947_data_out(3);
    CN237_sign_in(16) <= VN947_sign_out(3);
    CN237_data_in(17) <= VN1012_data_out(3);
    CN237_sign_in(17) <= VN1012_sign_out(3);
    CN237_data_in(18) <= VN1088_data_out(3);
    CN237_sign_in(18) <= VN1088_sign_out(3);
    CN237_data_in(19) <= VN1151_data_out(3);
    CN237_sign_in(19) <= VN1151_sign_out(3);
    CN237_data_in(20) <= VN1200_data_out(3);
    CN237_sign_in(20) <= VN1200_sign_out(3);
    CN237_data_in(21) <= VN1242_data_out(3);
    CN237_sign_in(21) <= VN1242_sign_out(3);
    CN237_data_in(22) <= VN1301_data_out(3);
    CN237_sign_in(22) <= VN1301_sign_out(3);
    CN237_data_in(23) <= VN1382_data_out(3);
    CN237_sign_in(23) <= VN1382_sign_out(3);
    CN237_data_in(24) <= VN1413_data_out(3);
    CN237_sign_in(24) <= VN1413_sign_out(3);
    CN237_data_in(25) <= VN1444_data_out(3);
    CN237_sign_in(25) <= VN1444_sign_out(3);
    CN237_data_in(26) <= VN1574_data_out(3);
    CN237_sign_in(26) <= VN1574_sign_out(3);
    CN237_data_in(27) <= VN1612_data_out(3);
    CN237_sign_in(27) <= VN1612_sign_out(3);
    CN237_data_in(28) <= VN1650_data_out(3);
    CN237_sign_in(28) <= VN1650_sign_out(3);
    CN237_data_in(29) <= VN1695_data_out(3);
    CN237_sign_in(29) <= VN1695_sign_out(3);
    CN237_data_in(30) <= VN1789_data_out(3);
    CN237_sign_in(30) <= VN1789_sign_out(3);
    CN237_data_in(31) <= VN1854_data_out(3);
    CN237_sign_in(31) <= VN1854_sign_out(3);
    CN238_data_in(0) <= VN9_data_out(3);
    CN238_sign_in(0) <= VN9_sign_out(3);
    CN238_data_in(1) <= VN103_data_out(3);
    CN238_sign_in(1) <= VN103_sign_out(3);
    CN238_data_in(2) <= VN113_data_out(3);
    CN238_sign_in(2) <= VN113_sign_out(3);
    CN238_data_in(3) <= VN179_data_out(3);
    CN238_sign_in(3) <= VN179_sign_out(3);
    CN238_data_in(4) <= VN236_data_out(3);
    CN238_sign_in(4) <= VN236_sign_out(3);
    CN238_data_in(5) <= VN294_data_out(3);
    CN238_sign_in(5) <= VN294_sign_out(3);
    CN238_data_in(6) <= VN383_data_out(3);
    CN238_sign_in(6) <= VN383_sign_out(3);
    CN238_data_in(7) <= VN416_data_out(3);
    CN238_sign_in(7) <= VN416_sign_out(3);
    CN238_data_in(8) <= VN498_data_out(3);
    CN238_sign_in(8) <= VN498_sign_out(3);
    CN238_data_in(9) <= VN507_data_out(3);
    CN238_sign_in(9) <= VN507_sign_out(3);
    CN238_data_in(10) <= VN582_data_out(3);
    CN238_sign_in(10) <= VN582_sign_out(3);
    CN238_data_in(11) <= VN641_data_out(3);
    CN238_sign_in(11) <= VN641_sign_out(3);
    CN238_data_in(12) <= VN687_data_out(3);
    CN238_sign_in(12) <= VN687_sign_out(3);
    CN238_data_in(13) <= VN728_data_out(3);
    CN238_sign_in(13) <= VN728_sign_out(3);
    CN238_data_in(14) <= VN824_data_out(3);
    CN238_sign_in(14) <= VN824_sign_out(3);
    CN238_data_in(15) <= VN837_data_out(3);
    CN238_sign_in(15) <= VN837_sign_out(3);
    CN238_data_in(16) <= VN891_data_out(3);
    CN238_sign_in(16) <= VN891_sign_out(3);
    CN238_data_in(17) <= VN948_data_out(3);
    CN238_sign_in(17) <= VN948_sign_out(3);
    CN238_data_in(18) <= VN1028_data_out(3);
    CN238_sign_in(18) <= VN1028_sign_out(3);
    CN238_data_in(19) <= VN1059_data_out(3);
    CN238_sign_in(19) <= VN1059_sign_out(3);
    CN238_data_in(20) <= VN1079_data_out(3);
    CN238_sign_in(20) <= VN1079_sign_out(3);
    CN238_data_in(21) <= VN1145_data_out(3);
    CN238_sign_in(21) <= VN1145_sign_out(3);
    CN238_data_in(22) <= VN1182_data_out(3);
    CN238_sign_in(22) <= VN1182_sign_out(3);
    CN238_data_in(23) <= VN1297_data_out(3);
    CN238_sign_in(23) <= VN1297_sign_out(3);
    CN238_data_in(24) <= VN1374_data_out(3);
    CN238_sign_in(24) <= VN1374_sign_out(3);
    CN238_data_in(25) <= VN1469_data_out(3);
    CN238_sign_in(25) <= VN1469_sign_out(3);
    CN238_data_in(26) <= VN1521_data_out(3);
    CN238_sign_in(26) <= VN1521_sign_out(3);
    CN238_data_in(27) <= VN1547_data_out(3);
    CN238_sign_in(27) <= VN1547_sign_out(3);
    CN238_data_in(28) <= VN1593_data_out(3);
    CN238_sign_in(28) <= VN1593_sign_out(3);
    CN238_data_in(29) <= VN1643_data_out(3);
    CN238_sign_in(29) <= VN1643_sign_out(3);
    CN238_data_in(30) <= VN1715_data_out(3);
    CN238_sign_in(30) <= VN1715_sign_out(3);
    CN238_data_in(31) <= VN1783_data_out(3);
    CN238_sign_in(31) <= VN1783_sign_out(3);
    CN239_data_in(0) <= VN8_data_out(3);
    CN239_sign_in(0) <= VN8_sign_out(3);
    CN239_data_in(1) <= VN98_data_out(3);
    CN239_sign_in(1) <= VN98_sign_out(3);
    CN239_data_in(2) <= VN158_data_out(3);
    CN239_sign_in(2) <= VN158_sign_out(3);
    CN239_data_in(3) <= VN223_data_out(3);
    CN239_sign_in(3) <= VN223_sign_out(3);
    CN239_data_in(4) <= VN264_data_out(3);
    CN239_sign_in(4) <= VN264_sign_out(3);
    CN239_data_in(5) <= VN284_data_out(3);
    CN239_sign_in(5) <= VN284_sign_out(3);
    CN239_data_in(6) <= VN360_data_out(3);
    CN239_sign_in(6) <= VN360_sign_out(3);
    CN239_data_in(7) <= VN392_data_out(3);
    CN239_sign_in(7) <= VN392_sign_out(3);
    CN239_data_in(8) <= VN452_data_out(3);
    CN239_sign_in(8) <= VN452_sign_out(3);
    CN239_data_in(9) <= VN513_data_out(3);
    CN239_sign_in(9) <= VN513_sign_out(3);
    CN239_data_in(10) <= VN596_data_out(3);
    CN239_sign_in(10) <= VN596_sign_out(3);
    CN239_data_in(11) <= VN620_data_out(3);
    CN239_sign_in(11) <= VN620_sign_out(3);
    CN239_data_in(12) <= VN710_data_out(3);
    CN239_sign_in(12) <= VN710_sign_out(3);
    CN239_data_in(13) <= VN752_data_out(3);
    CN239_sign_in(13) <= VN752_sign_out(3);
    CN239_data_in(14) <= VN829_data_out(3);
    CN239_sign_in(14) <= VN829_sign_out(3);
    CN239_data_in(15) <= VN866_data_out(3);
    CN239_sign_in(15) <= VN866_sign_out(3);
    CN239_data_in(16) <= VN926_data_out(3);
    CN239_sign_in(16) <= VN926_sign_out(3);
    CN239_data_in(17) <= VN983_data_out(3);
    CN239_sign_in(17) <= VN983_sign_out(3);
    CN239_data_in(18) <= VN1032_data_out(3);
    CN239_sign_in(18) <= VN1032_sign_out(3);
    CN239_data_in(19) <= VN1099_data_out(3);
    CN239_sign_in(19) <= VN1099_sign_out(3);
    CN239_data_in(20) <= VN1127_data_out(3);
    CN239_sign_in(20) <= VN1127_sign_out(3);
    CN239_data_in(21) <= VN1185_data_out(3);
    CN239_sign_in(21) <= VN1185_sign_out(3);
    CN239_data_in(22) <= VN1424_data_out(3);
    CN239_sign_in(22) <= VN1424_sign_out(3);
    CN239_data_in(23) <= VN1572_data_out(3);
    CN239_sign_in(23) <= VN1572_sign_out(3);
    CN239_data_in(24) <= VN1587_data_out(3);
    CN239_sign_in(24) <= VN1587_sign_out(3);
    CN239_data_in(25) <= VN1717_data_out(3);
    CN239_sign_in(25) <= VN1717_sign_out(3);
    CN239_data_in(26) <= VN1794_data_out(3);
    CN239_sign_in(26) <= VN1794_sign_out(3);
    CN239_data_in(27) <= VN1811_data_out(3);
    CN239_sign_in(27) <= VN1811_sign_out(3);
    CN239_data_in(28) <= VN1814_data_out(3);
    CN239_sign_in(28) <= VN1814_sign_out(3);
    CN239_data_in(29) <= VN1817_data_out(3);
    CN239_sign_in(29) <= VN1817_sign_out(3);
    CN239_data_in(30) <= VN1866_data_out(3);
    CN239_sign_in(30) <= VN1866_sign_out(3);
    CN239_data_in(31) <= VN1890_data_out(3);
    CN239_sign_in(31) <= VN1890_sign_out(3);
    CN240_data_in(0) <= VN7_data_out(3);
    CN240_sign_in(0) <= VN7_sign_out(3);
    CN240_data_in(1) <= VN81_data_out(3);
    CN240_sign_in(1) <= VN81_sign_out(3);
    CN240_data_in(2) <= VN116_data_out(3);
    CN240_sign_in(2) <= VN116_sign_out(3);
    CN240_data_in(3) <= VN210_data_out(3);
    CN240_sign_in(3) <= VN210_sign_out(3);
    CN240_data_in(4) <= VN277_data_out(3);
    CN240_sign_in(4) <= VN277_sign_out(3);
    CN240_data_in(5) <= VN324_data_out(3);
    CN240_sign_in(5) <= VN324_sign_out(3);
    CN240_data_in(6) <= VN343_data_out(3);
    CN240_sign_in(6) <= VN343_sign_out(3);
    CN240_data_in(7) <= VN444_data_out(3);
    CN240_sign_in(7) <= VN444_sign_out(3);
    CN240_data_in(8) <= VN502_data_out(3);
    CN240_sign_in(8) <= VN502_sign_out(3);
    CN240_data_in(9) <= VN534_data_out(3);
    CN240_sign_in(9) <= VN534_sign_out(3);
    CN240_data_in(10) <= VN589_data_out(3);
    CN240_sign_in(10) <= VN589_sign_out(3);
    CN240_data_in(11) <= VN637_data_out(3);
    CN240_sign_in(11) <= VN637_sign_out(3);
    CN240_data_in(12) <= VN708_data_out(3);
    CN240_sign_in(12) <= VN708_sign_out(3);
    CN240_data_in(13) <= VN734_data_out(3);
    CN240_sign_in(13) <= VN734_sign_out(3);
    CN240_data_in(14) <= VN814_data_out(3);
    CN240_sign_in(14) <= VN814_sign_out(3);
    CN240_data_in(15) <= VN845_data_out(3);
    CN240_sign_in(15) <= VN845_sign_out(3);
    CN240_data_in(16) <= VN907_data_out(3);
    CN240_sign_in(16) <= VN907_sign_out(3);
    CN240_data_in(17) <= VN975_data_out(3);
    CN240_sign_in(17) <= VN975_sign_out(3);
    CN240_data_in(18) <= VN1105_data_out(3);
    CN240_sign_in(18) <= VN1105_sign_out(3);
    CN240_data_in(19) <= VN1113_data_out(3);
    CN240_sign_in(19) <= VN1113_sign_out(3);
    CN240_data_in(20) <= VN1134_data_out(3);
    CN240_sign_in(20) <= VN1134_sign_out(3);
    CN240_data_in(21) <= VN1171_data_out(3);
    CN240_sign_in(21) <= VN1171_sign_out(3);
    CN240_data_in(22) <= VN1259_data_out(3);
    CN240_sign_in(22) <= VN1259_sign_out(3);
    CN240_data_in(23) <= VN1339_data_out(3);
    CN240_sign_in(23) <= VN1339_sign_out(3);
    CN240_data_in(24) <= VN1394_data_out(3);
    CN240_sign_in(24) <= VN1394_sign_out(3);
    CN240_data_in(25) <= VN1437_data_out(3);
    CN240_sign_in(25) <= VN1437_sign_out(3);
    CN240_data_in(26) <= VN1505_data_out(3);
    CN240_sign_in(26) <= VN1505_sign_out(3);
    CN240_data_in(27) <= VN1605_data_out(3);
    CN240_sign_in(27) <= VN1605_sign_out(3);
    CN240_data_in(28) <= VN1686_data_out(3);
    CN240_sign_in(28) <= VN1686_sign_out(3);
    CN240_data_in(29) <= VN1703_data_out(3);
    CN240_sign_in(29) <= VN1703_sign_out(3);
    CN240_data_in(30) <= VN1806_data_out(3);
    CN240_sign_in(30) <= VN1806_sign_out(3);
    CN240_data_in(31) <= VN1855_data_out(3);
    CN240_sign_in(31) <= VN1855_sign_out(3);
    CN241_data_in(0) <= VN6_data_out(3);
    CN241_sign_in(0) <= VN6_sign_out(3);
    CN241_data_in(1) <= VN88_data_out(3);
    CN241_sign_in(1) <= VN88_sign_out(3);
    CN241_data_in(2) <= VN175_data_out(3);
    CN241_sign_in(2) <= VN175_sign_out(3);
    CN241_data_in(3) <= VN250_data_out(3);
    CN241_sign_in(3) <= VN250_sign_out(3);
    CN241_data_in(4) <= VN285_data_out(3);
    CN241_sign_in(4) <= VN285_sign_out(3);
    CN241_data_in(5) <= VN355_data_out(3);
    CN241_sign_in(5) <= VN355_sign_out(3);
    CN241_data_in(6) <= VN403_data_out(3);
    CN241_sign_in(6) <= VN403_sign_out(3);
    CN241_data_in(7) <= VN449_data_out(3);
    CN241_sign_in(7) <= VN449_sign_out(3);
    CN241_data_in(8) <= VN532_data_out(3);
    CN241_sign_in(8) <= VN532_sign_out(3);
    CN241_data_in(9) <= VN565_data_out(3);
    CN241_sign_in(9) <= VN565_sign_out(3);
    CN241_data_in(10) <= VN685_data_out(3);
    CN241_sign_in(10) <= VN685_sign_out(3);
    CN241_data_in(11) <= VN745_data_out(3);
    CN241_sign_in(11) <= VN745_sign_out(3);
    CN241_data_in(12) <= VN816_data_out(3);
    CN241_sign_in(12) <= VN816_sign_out(3);
    CN241_data_in(13) <= VN992_data_out(3);
    CN241_sign_in(13) <= VN992_sign_out(3);
    CN241_data_in(14) <= VN1031_data_out(3);
    CN241_sign_in(14) <= VN1031_sign_out(3);
    CN241_data_in(15) <= VN1090_data_out(3);
    CN241_sign_in(15) <= VN1090_sign_out(3);
    CN241_data_in(16) <= VN1157_data_out(3);
    CN241_sign_in(16) <= VN1157_sign_out(3);
    CN241_data_in(17) <= VN1168_data_out(3);
    CN241_sign_in(17) <= VN1168_sign_out(3);
    CN241_data_in(18) <= VN1201_data_out(3);
    CN241_sign_in(18) <= VN1201_sign_out(3);
    CN241_data_in(19) <= VN1245_data_out(3);
    CN241_sign_in(19) <= VN1245_sign_out(3);
    CN241_data_in(20) <= VN1388_data_out(3);
    CN241_sign_in(20) <= VN1388_sign_out(3);
    CN241_data_in(21) <= VN1463_data_out(3);
    CN241_sign_in(21) <= VN1463_sign_out(3);
    CN241_data_in(22) <= VN1536_data_out(3);
    CN241_sign_in(22) <= VN1536_sign_out(3);
    CN241_data_in(23) <= VN1548_data_out(3);
    CN241_sign_in(23) <= VN1548_sign_out(3);
    CN241_data_in(24) <= VN1624_data_out(3);
    CN241_sign_in(24) <= VN1624_sign_out(3);
    CN241_data_in(25) <= VN1690_data_out(3);
    CN241_sign_in(25) <= VN1690_sign_out(3);
    CN241_data_in(26) <= VN1802_data_out(3);
    CN241_sign_in(26) <= VN1802_sign_out(3);
    CN241_data_in(27) <= VN1891_data_out(3);
    CN241_sign_in(27) <= VN1891_sign_out(3);
    CN241_data_in(28) <= VN1893_data_out(3);
    CN241_sign_in(28) <= VN1893_sign_out(3);
    CN241_data_in(29) <= VN1901_data_out(3);
    CN241_sign_in(29) <= VN1901_sign_out(3);
    CN241_data_in(30) <= VN1941_data_out(3);
    CN241_sign_in(30) <= VN1941_sign_out(3);
    CN241_data_in(31) <= VN1947_data_out(3);
    CN241_sign_in(31) <= VN1947_sign_out(3);
    CN242_data_in(0) <= VN5_data_out(3);
    CN242_sign_in(0) <= VN5_sign_out(3);
    CN242_data_in(1) <= VN108_data_out(3);
    CN242_sign_in(1) <= VN108_sign_out(3);
    CN242_data_in(2) <= VN146_data_out(3);
    CN242_sign_in(2) <= VN146_sign_out(3);
    CN242_data_in(3) <= VN203_data_out(3);
    CN242_sign_in(3) <= VN203_sign_out(3);
    CN242_data_in(4) <= VN231_data_out(3);
    CN242_sign_in(4) <= VN231_sign_out(3);
    CN242_data_in(5) <= VN303_data_out(3);
    CN242_sign_in(5) <= VN303_sign_out(3);
    CN242_data_in(6) <= VN367_data_out(3);
    CN242_sign_in(6) <= VN367_sign_out(3);
    CN242_data_in(7) <= VN396_data_out(3);
    CN242_sign_in(7) <= VN396_sign_out(3);
    CN242_data_in(8) <= VN495_data_out(3);
    CN242_sign_in(8) <= VN495_sign_out(3);
    CN242_data_in(9) <= VN511_data_out(3);
    CN242_sign_in(9) <= VN511_sign_out(3);
    CN242_data_in(10) <= VN575_data_out(3);
    CN242_sign_in(10) <= VN575_sign_out(3);
    CN242_data_in(11) <= VN650_data_out(3);
    CN242_sign_in(11) <= VN650_sign_out(3);
    CN242_data_in(12) <= VN720_data_out(3);
    CN242_sign_in(12) <= VN720_sign_out(3);
    CN242_data_in(13) <= VN753_data_out(3);
    CN242_sign_in(13) <= VN753_sign_out(3);
    CN242_data_in(14) <= VN786_data_out(3);
    CN242_sign_in(14) <= VN786_sign_out(3);
    CN242_data_in(15) <= VN880_data_out(3);
    CN242_sign_in(15) <= VN880_sign_out(3);
    CN242_data_in(16) <= VN894_data_out(3);
    CN242_sign_in(16) <= VN894_sign_out(3);
    CN242_data_in(17) <= VN997_data_out(3);
    CN242_sign_in(17) <= VN997_sign_out(3);
    CN242_data_in(18) <= VN1003_data_out(3);
    CN242_sign_in(18) <= VN1003_sign_out(3);
    CN242_data_in(19) <= VN1026_data_out(3);
    CN242_sign_in(19) <= VN1026_sign_out(3);
    CN242_data_in(20) <= VN1092_data_out(3);
    CN242_sign_in(20) <= VN1092_sign_out(3);
    CN242_data_in(21) <= VN1155_data_out(3);
    CN242_sign_in(21) <= VN1155_sign_out(3);
    CN242_data_in(22) <= VN1319_data_out(3);
    CN242_sign_in(22) <= VN1319_sign_out(3);
    CN242_data_in(23) <= VN1338_data_out(3);
    CN242_sign_in(23) <= VN1338_sign_out(3);
    CN242_data_in(24) <= VN1471_data_out(3);
    CN242_sign_in(24) <= VN1471_sign_out(3);
    CN242_data_in(25) <= VN1522_data_out(3);
    CN242_sign_in(25) <= VN1522_sign_out(3);
    CN242_data_in(26) <= VN1596_data_out(3);
    CN242_sign_in(26) <= VN1596_sign_out(3);
    CN242_data_in(27) <= VN1638_data_out(3);
    CN242_sign_in(27) <= VN1638_sign_out(3);
    CN242_data_in(28) <= VN1666_data_out(3);
    CN242_sign_in(28) <= VN1666_sign_out(3);
    CN242_data_in(29) <= VN1696_data_out(3);
    CN242_sign_in(29) <= VN1696_sign_out(3);
    CN242_data_in(30) <= VN1786_data_out(3);
    CN242_sign_in(30) <= VN1786_sign_out(3);
    CN242_data_in(31) <= VN1856_data_out(3);
    CN242_sign_in(31) <= VN1856_sign_out(3);
    CN243_data_in(0) <= VN4_data_out(3);
    CN243_sign_in(0) <= VN4_sign_out(3);
    CN243_data_in(1) <= VN106_data_out(3);
    CN243_sign_in(1) <= VN106_sign_out(3);
    CN243_data_in(2) <= VN141_data_out(3);
    CN243_sign_in(2) <= VN141_sign_out(3);
    CN243_data_in(3) <= VN200_data_out(3);
    CN243_sign_in(3) <= VN200_sign_out(3);
    CN243_data_in(4) <= VN252_data_out(3);
    CN243_sign_in(4) <= VN252_sign_out(3);
    CN243_data_in(5) <= VN312_data_out(3);
    CN243_sign_in(5) <= VN312_sign_out(3);
    CN243_data_in(6) <= VN337_data_out(3);
    CN243_sign_in(6) <= VN337_sign_out(3);
    CN243_data_in(7) <= VN427_data_out(3);
    CN243_sign_in(7) <= VN427_sign_out(3);
    CN243_data_in(8) <= VN476_data_out(3);
    CN243_sign_in(8) <= VN476_sign_out(3);
    CN243_data_in(9) <= VN548_data_out(3);
    CN243_sign_in(9) <= VN548_sign_out(3);
    CN243_data_in(10) <= VN569_data_out(3);
    CN243_sign_in(10) <= VN569_sign_out(3);
    CN243_data_in(11) <= VN670_data_out(3);
    CN243_sign_in(11) <= VN670_sign_out(3);
    CN243_data_in(12) <= VN727_data_out(3);
    CN243_sign_in(12) <= VN727_sign_out(3);
    CN243_data_in(13) <= VN822_data_out(3);
    CN243_sign_in(13) <= VN822_sign_out(3);
    CN243_data_in(14) <= VN1009_data_out(3);
    CN243_sign_in(14) <= VN1009_sign_out(3);
    CN243_data_in(15) <= VN1064_data_out(3);
    CN243_sign_in(15) <= VN1064_sign_out(3);
    CN243_data_in(16) <= VN1132_data_out(3);
    CN243_sign_in(16) <= VN1132_sign_out(3);
    CN243_data_in(17) <= VN1281_data_out(3);
    CN243_sign_in(17) <= VN1281_sign_out(3);
    CN243_data_in(18) <= VN1335_data_out(3);
    CN243_sign_in(18) <= VN1335_sign_out(3);
    CN243_data_in(19) <= VN1439_data_out(3);
    CN243_sign_in(19) <= VN1439_sign_out(3);
    CN243_data_in(20) <= VN1503_data_out(3);
    CN243_sign_in(20) <= VN1503_sign_out(3);
    CN243_data_in(21) <= VN1598_data_out(3);
    CN243_sign_in(21) <= VN1598_sign_out(3);
    CN243_data_in(22) <= VN1675_data_out(3);
    CN243_sign_in(22) <= VN1675_sign_out(3);
    CN243_data_in(23) <= VN1744_data_out(3);
    CN243_sign_in(23) <= VN1744_sign_out(3);
    CN243_data_in(24) <= VN1764_data_out(3);
    CN243_sign_in(24) <= VN1764_sign_out(3);
    CN243_data_in(25) <= VN1816_data_out(3);
    CN243_sign_in(25) <= VN1816_sign_out(3);
    CN243_data_in(26) <= VN1872_data_out(3);
    CN243_sign_in(26) <= VN1872_sign_out(3);
    CN243_data_in(27) <= VN1904_data_out(3);
    CN243_sign_in(27) <= VN1904_sign_out(3);
    CN243_data_in(28) <= VN1927_data_out(3);
    CN243_sign_in(28) <= VN1927_sign_out(3);
    CN243_data_in(29) <= VN1950_data_out(3);
    CN243_sign_in(29) <= VN1950_sign_out(3);
    CN243_data_in(30) <= VN1968_data_out(3);
    CN243_sign_in(30) <= VN1968_sign_out(3);
    CN243_data_in(31) <= VN1971_data_out(3);
    CN243_sign_in(31) <= VN1971_sign_out(3);
    CN244_data_in(0) <= VN147_data_out(3);
    CN244_sign_in(0) <= VN147_sign_out(3);
    CN244_data_in(1) <= VN266_data_out(3);
    CN244_sign_in(1) <= VN266_sign_out(3);
    CN244_data_in(2) <= VN385_data_out(3);
    CN244_sign_in(2) <= VN385_sign_out(3);
    CN244_data_in(3) <= VN459_data_out(3);
    CN244_sign_in(3) <= VN459_sign_out(3);
    CN244_data_in(4) <= VN551_data_out(3);
    CN244_sign_in(4) <= VN551_sign_out(3);
    CN244_data_in(5) <= VN572_data_out(3);
    CN244_sign_in(5) <= VN572_sign_out(3);
    CN244_data_in(6) <= VN665_data_out(3);
    CN244_sign_in(6) <= VN665_sign_out(3);
    CN244_data_in(7) <= VN741_data_out(3);
    CN244_sign_in(7) <= VN741_sign_out(3);
    CN244_data_in(8) <= VN840_data_out(3);
    CN244_sign_in(8) <= VN840_sign_out(3);
    CN244_data_in(9) <= VN890_data_out(3);
    CN244_sign_in(9) <= VN890_sign_out(3);
    CN244_data_in(10) <= VN996_data_out(3);
    CN244_sign_in(10) <= VN996_sign_out(3);
    CN244_data_in(11) <= VN1016_data_out(3);
    CN244_sign_in(11) <= VN1016_sign_out(3);
    CN244_data_in(12) <= VN1178_data_out(3);
    CN244_sign_in(12) <= VN1178_sign_out(3);
    CN244_data_in(13) <= VN1269_data_out(3);
    CN244_sign_in(13) <= VN1269_sign_out(3);
    CN244_data_in(14) <= VN1305_data_out(3);
    CN244_sign_in(14) <= VN1305_sign_out(3);
    CN244_data_in(15) <= VN1371_data_out(3);
    CN244_sign_in(15) <= VN1371_sign_out(3);
    CN244_data_in(16) <= VN1421_data_out(3);
    CN244_sign_in(16) <= VN1421_sign_out(3);
    CN244_data_in(17) <= VN1482_data_out(3);
    CN244_sign_in(17) <= VN1482_sign_out(3);
    CN244_data_in(18) <= VN1554_data_out(3);
    CN244_sign_in(18) <= VN1554_sign_out(3);
    CN244_data_in(19) <= VN1609_data_out(3);
    CN244_sign_in(19) <= VN1609_sign_out(3);
    CN244_data_in(20) <= VN1716_data_out(3);
    CN244_sign_in(20) <= VN1716_sign_out(3);
    CN244_data_in(21) <= VN1807_data_out(3);
    CN244_sign_in(21) <= VN1807_sign_out(3);
    CN244_data_in(22) <= VN1980_data_out(3);
    CN244_sign_in(22) <= VN1980_sign_out(3);
    CN244_data_in(23) <= VN1986_data_out(3);
    CN244_sign_in(23) <= VN1986_sign_out(3);
    CN244_data_in(24) <= VN1987_data_out(3);
    CN244_sign_in(24) <= VN1987_sign_out(3);
    CN244_data_in(25) <= VN1992_data_out(3);
    CN244_sign_in(25) <= VN1992_sign_out(3);
    CN244_data_in(26) <= VN1999_data_out(3);
    CN244_sign_in(26) <= VN1999_sign_out(3);
    CN244_data_in(27) <= VN2011_data_out(3);
    CN244_sign_in(27) <= VN2011_sign_out(3);
    CN244_data_in(28) <= VN2014_data_out(3);
    CN244_sign_in(28) <= VN2014_sign_out(3);
    CN244_data_in(29) <= VN2024_data_out(3);
    CN244_sign_in(29) <= VN2024_sign_out(3);
    CN244_data_in(30) <= VN2030_data_out(3);
    CN244_sign_in(30) <= VN2030_sign_out(3);
    CN244_data_in(31) <= VN2038_data_out(3);
    CN244_sign_in(31) <= VN2038_sign_out(3);
    CN245_data_in(0) <= VN3_data_out(3);
    CN245_sign_in(0) <= VN3_sign_out(3);
    CN245_data_in(1) <= VN66_data_out(3);
    CN245_sign_in(1) <= VN66_sign_out(3);
    CN245_data_in(2) <= VN136_data_out(3);
    CN245_sign_in(2) <= VN136_sign_out(3);
    CN245_data_in(3) <= VN207_data_out(3);
    CN245_sign_in(3) <= VN207_sign_out(3);
    CN245_data_in(4) <= VN262_data_out(3);
    CN245_sign_in(4) <= VN262_sign_out(3);
    CN245_data_in(5) <= VN313_data_out(3);
    CN245_sign_in(5) <= VN313_sign_out(3);
    CN245_data_in(6) <= VN370_data_out(3);
    CN245_sign_in(6) <= VN370_sign_out(3);
    CN245_data_in(7) <= VN431_data_out(3);
    CN245_sign_in(7) <= VN431_sign_out(3);
    CN245_data_in(8) <= VN471_data_out(3);
    CN245_sign_in(8) <= VN471_sign_out(3);
    CN245_data_in(9) <= VN535_data_out(3);
    CN245_sign_in(9) <= VN535_sign_out(3);
    CN245_data_in(10) <= VN562_data_out(3);
    CN245_sign_in(10) <= VN562_sign_out(3);
    CN245_data_in(11) <= VN686_data_out(3);
    CN245_sign_in(11) <= VN686_sign_out(3);
    CN245_data_in(12) <= VN769_data_out(3);
    CN245_sign_in(12) <= VN769_sign_out(3);
    CN245_data_in(13) <= VN787_data_out(3);
    CN245_sign_in(13) <= VN787_sign_out(3);
    CN245_data_in(14) <= VN862_data_out(3);
    CN245_sign_in(14) <= VN862_sign_out(3);
    CN245_data_in(15) <= VN918_data_out(3);
    CN245_sign_in(15) <= VN918_sign_out(3);
    CN245_data_in(16) <= VN991_data_out(3);
    CN245_sign_in(16) <= VN991_sign_out(3);
    CN245_data_in(17) <= VN1037_data_out(3);
    CN245_sign_in(17) <= VN1037_sign_out(3);
    CN245_data_in(18) <= VN1109_data_out(3);
    CN245_sign_in(18) <= VN1109_sign_out(3);
    CN245_data_in(19) <= VN1115_data_out(3);
    CN245_sign_in(19) <= VN1115_sign_out(3);
    CN245_data_in(20) <= VN1203_data_out(3);
    CN245_sign_in(20) <= VN1203_sign_out(3);
    CN245_data_in(21) <= VN1220_data_out(3);
    CN245_sign_in(21) <= VN1220_sign_out(3);
    CN245_data_in(22) <= VN1254_data_out(3);
    CN245_sign_in(22) <= VN1254_sign_out(3);
    CN245_data_in(23) <= VN1378_data_out(3);
    CN245_sign_in(23) <= VN1378_sign_out(3);
    CN245_data_in(24) <= VN1418_data_out(3);
    CN245_sign_in(24) <= VN1418_sign_out(3);
    CN245_data_in(25) <= VN1467_data_out(3);
    CN245_sign_in(25) <= VN1467_sign_out(3);
    CN245_data_in(26) <= VN1528_data_out(3);
    CN245_sign_in(26) <= VN1528_sign_out(3);
    CN245_data_in(27) <= VN1603_data_out(3);
    CN245_sign_in(27) <= VN1603_sign_out(3);
    CN245_data_in(28) <= VN1637_data_out(3);
    CN245_sign_in(28) <= VN1637_sign_out(3);
    CN245_data_in(29) <= VN1653_data_out(3);
    CN245_sign_in(29) <= VN1653_sign_out(3);
    CN245_data_in(30) <= VN1759_data_out(3);
    CN245_sign_in(30) <= VN1759_sign_out(3);
    CN245_data_in(31) <= VN1857_data_out(3);
    CN245_sign_in(31) <= VN1857_sign_out(3);
    CN246_data_in(0) <= VN2_data_out(3);
    CN246_sign_in(0) <= VN2_sign_out(3);
    CN246_data_in(1) <= VN69_data_out(3);
    CN246_sign_in(1) <= VN69_sign_out(3);
    CN246_data_in(2) <= VN161_data_out(3);
    CN246_sign_in(2) <= VN161_sign_out(3);
    CN246_data_in(3) <= VN185_data_out(3);
    CN246_sign_in(3) <= VN185_sign_out(3);
    CN246_data_in(4) <= VN226_data_out(3);
    CN246_sign_in(4) <= VN226_sign_out(3);
    CN246_data_in(5) <= VN302_data_out(3);
    CN246_sign_in(5) <= VN302_sign_out(3);
    CN246_data_in(6) <= VN388_data_out(3);
    CN246_sign_in(6) <= VN388_sign_out(3);
    CN246_data_in(7) <= VN435_data_out(3);
    CN246_sign_in(7) <= VN435_sign_out(3);
    CN246_data_in(8) <= VN481_data_out(3);
    CN246_sign_in(8) <= VN481_sign_out(3);
    CN246_data_in(9) <= VN512_data_out(3);
    CN246_sign_in(9) <= VN512_sign_out(3);
    CN246_data_in(10) <= VN597_data_out(3);
    CN246_sign_in(10) <= VN597_sign_out(3);
    CN246_data_in(11) <= VN618_data_out(3);
    CN246_sign_in(11) <= VN618_sign_out(3);
    CN246_data_in(12) <= VN707_data_out(3);
    CN246_sign_in(12) <= VN707_sign_out(3);
    CN246_data_in(13) <= VN748_data_out(3);
    CN246_sign_in(13) <= VN748_sign_out(3);
    CN246_data_in(14) <= VN815_data_out(3);
    CN246_sign_in(14) <= VN815_sign_out(3);
    CN246_data_in(15) <= VN863_data_out(3);
    CN246_sign_in(15) <= VN863_sign_out(3);
    CN246_data_in(16) <= VN903_data_out(3);
    CN246_sign_in(16) <= VN903_sign_out(3);
    CN246_data_in(17) <= VN972_data_out(3);
    CN246_sign_in(17) <= VN972_sign_out(3);
    CN246_data_in(18) <= VN1035_data_out(3);
    CN246_sign_in(18) <= VN1035_sign_out(3);
    CN246_data_in(19) <= VN1065_data_out(3);
    CN246_sign_in(19) <= VN1065_sign_out(3);
    CN246_data_in(20) <= VN1158_data_out(3);
    CN246_sign_in(20) <= VN1158_sign_out(3);
    CN246_data_in(21) <= VN1194_data_out(3);
    CN246_sign_in(21) <= VN1194_sign_out(3);
    CN246_data_in(22) <= VN1222_data_out(3);
    CN246_sign_in(22) <= VN1222_sign_out(3);
    CN246_data_in(23) <= VN1311_data_out(3);
    CN246_sign_in(23) <= VN1311_sign_out(3);
    CN246_data_in(24) <= VN1345_data_out(3);
    CN246_sign_in(24) <= VN1345_sign_out(3);
    CN246_data_in(25) <= VN1384_data_out(3);
    CN246_sign_in(25) <= VN1384_sign_out(3);
    CN246_data_in(26) <= VN1524_data_out(3);
    CN246_sign_in(26) <= VN1524_sign_out(3);
    CN246_data_in(27) <= VN1540_data_out(3);
    CN246_sign_in(27) <= VN1540_sign_out(3);
    CN246_data_in(28) <= VN1630_data_out(3);
    CN246_sign_in(28) <= VN1630_sign_out(3);
    CN246_data_in(29) <= VN1661_data_out(3);
    CN246_sign_in(29) <= VN1661_sign_out(3);
    CN246_data_in(30) <= VN1709_data_out(3);
    CN246_sign_in(30) <= VN1709_sign_out(3);
    CN246_data_in(31) <= VN1784_data_out(3);
    CN246_sign_in(31) <= VN1784_sign_out(3);
    CN247_data_in(0) <= VN1_data_out(3);
    CN247_sign_in(0) <= VN1_sign_out(3);
    CN247_data_in(1) <= VN109_data_out(3);
    CN247_sign_in(1) <= VN109_sign_out(3);
    CN247_data_in(2) <= VN168_data_out(3);
    CN247_sign_in(2) <= VN168_sign_out(3);
    CN247_data_in(3) <= VN194_data_out(3);
    CN247_sign_in(3) <= VN194_sign_out(3);
    CN247_data_in(4) <= VN247_data_out(3);
    CN247_sign_in(4) <= VN247_sign_out(3);
    CN247_data_in(5) <= VN327_data_out(3);
    CN247_sign_in(5) <= VN327_sign_out(3);
    CN247_data_in(6) <= VN349_data_out(3);
    CN247_sign_in(6) <= VN349_sign_out(3);
    CN247_data_in(7) <= VN424_data_out(3);
    CN247_sign_in(7) <= VN424_sign_out(3);
    CN247_data_in(8) <= VN453_data_out(3);
    CN247_sign_in(8) <= VN453_sign_out(3);
    CN247_data_in(9) <= VN531_data_out(3);
    CN247_sign_in(9) <= VN531_sign_out(3);
    CN247_data_in(10) <= VN581_data_out(3);
    CN247_sign_in(10) <= VN581_sign_out(3);
    CN247_data_in(11) <= VN646_data_out(3);
    CN247_sign_in(11) <= VN646_sign_out(3);
    CN247_data_in(12) <= VN677_data_out(3);
    CN247_sign_in(12) <= VN677_sign_out(3);
    CN247_data_in(13) <= VN771_data_out(3);
    CN247_sign_in(13) <= VN771_sign_out(3);
    CN247_data_in(14) <= VN828_data_out(3);
    CN247_sign_in(14) <= VN828_sign_out(3);
    CN247_data_in(15) <= VN839_data_out(3);
    CN247_sign_in(15) <= VN839_sign_out(3);
    CN247_data_in(16) <= VN928_data_out(3);
    CN247_sign_in(16) <= VN928_sign_out(3);
    CN247_data_in(17) <= VN980_data_out(3);
    CN247_sign_in(17) <= VN980_sign_out(3);
    CN247_data_in(18) <= VN1014_data_out(3);
    CN247_sign_in(18) <= VN1014_sign_out(3);
    CN247_data_in(19) <= VN1091_data_out(3);
    CN247_sign_in(19) <= VN1091_sign_out(3);
    CN247_data_in(20) <= VN1133_data_out(3);
    CN247_sign_in(20) <= VN1133_sign_out(3);
    CN247_data_in(21) <= VN1183_data_out(3);
    CN247_sign_in(21) <= VN1183_sign_out(3);
    CN247_data_in(22) <= VN1271_data_out(3);
    CN247_sign_in(22) <= VN1271_sign_out(3);
    CN247_data_in(23) <= VN1323_data_out(3);
    CN247_sign_in(23) <= VN1323_sign_out(3);
    CN247_data_in(24) <= VN1333_data_out(3);
    CN247_sign_in(24) <= VN1333_sign_out(3);
    CN247_data_in(25) <= VN1343_data_out(3);
    CN247_sign_in(25) <= VN1343_sign_out(3);
    CN247_data_in(26) <= VN1447_data_out(3);
    CN247_sign_in(26) <= VN1447_sign_out(3);
    CN247_data_in(27) <= VN1483_data_out(3);
    CN247_sign_in(27) <= VN1483_sign_out(3);
    CN247_data_in(28) <= VN1646_data_out(3);
    CN247_sign_in(28) <= VN1646_sign_out(3);
    CN247_data_in(29) <= VN1699_data_out(3);
    CN247_sign_in(29) <= VN1699_sign_out(3);
    CN247_data_in(30) <= VN1755_data_out(3);
    CN247_sign_in(30) <= VN1755_sign_out(3);
    CN247_data_in(31) <= VN1858_data_out(3);
    CN247_sign_in(31) <= VN1858_sign_out(3);
    CN248_data_in(0) <= VN0_data_out(3);
    CN248_sign_in(0) <= VN0_sign_out(3);
    CN248_data_in(1) <= VN87_data_out(3);
    CN248_sign_in(1) <= VN87_sign_out(3);
    CN248_data_in(2) <= VN151_data_out(3);
    CN248_sign_in(2) <= VN151_sign_out(3);
    CN248_data_in(3) <= VN189_data_out(3);
    CN248_sign_in(3) <= VN189_sign_out(3);
    CN248_data_in(4) <= VN248_data_out(3);
    CN248_sign_in(4) <= VN248_sign_out(3);
    CN248_data_in(5) <= VN280_data_out(3);
    CN248_sign_in(5) <= VN280_sign_out(3);
    CN248_data_in(6) <= VN357_data_out(3);
    CN248_sign_in(6) <= VN357_sign_out(3);
    CN248_data_in(7) <= VN404_data_out(3);
    CN248_sign_in(7) <= VN404_sign_out(3);
    CN248_data_in(8) <= VN497_data_out(3);
    CN248_sign_in(8) <= VN497_sign_out(3);
    CN248_data_in(9) <= VN559_data_out(3);
    CN248_sign_in(9) <= VN559_sign_out(3);
    CN248_data_in(10) <= VN592_data_out(3);
    CN248_sign_in(10) <= VN592_sign_out(3);
    CN248_data_in(11) <= VN643_data_out(3);
    CN248_sign_in(11) <= VN643_sign_out(3);
    CN248_data_in(12) <= VN717_data_out(3);
    CN248_sign_in(12) <= VN717_sign_out(3);
    CN248_data_in(13) <= VN729_data_out(3);
    CN248_sign_in(13) <= VN729_sign_out(3);
    CN248_data_in(14) <= VN801_data_out(3);
    CN248_sign_in(14) <= VN801_sign_out(3);
    CN248_data_in(15) <= VN831_data_out(3);
    CN248_sign_in(15) <= VN831_sign_out(3);
    CN248_data_in(16) <= VN920_data_out(3);
    CN248_sign_in(16) <= VN920_sign_out(3);
    CN248_data_in(17) <= VN1002_data_out(3);
    CN248_sign_in(17) <= VN1002_sign_out(3);
    CN248_data_in(18) <= VN1051_data_out(3);
    CN248_sign_in(18) <= VN1051_sign_out(3);
    CN248_data_in(19) <= VN1104_data_out(3);
    CN248_sign_in(19) <= VN1104_sign_out(3);
    CN248_data_in(20) <= VN1154_data_out(3);
    CN248_sign_in(20) <= VN1154_sign_out(3);
    CN248_data_in(21) <= VN1199_data_out(3);
    CN248_sign_in(21) <= VN1199_sign_out(3);
    CN248_data_in(22) <= VN1257_data_out(3);
    CN248_sign_in(22) <= VN1257_sign_out(3);
    CN248_data_in(23) <= VN1279_data_out(3);
    CN248_sign_in(23) <= VN1279_sign_out(3);
    CN248_data_in(24) <= VN1377_data_out(3);
    CN248_sign_in(24) <= VN1377_sign_out(3);
    CN248_data_in(25) <= VN1401_data_out(3);
    CN248_sign_in(25) <= VN1401_sign_out(3);
    CN248_data_in(26) <= VN1431_data_out(3);
    CN248_sign_in(26) <= VN1431_sign_out(3);
    CN248_data_in(27) <= VN1490_data_out(3);
    CN248_sign_in(27) <= VN1490_sign_out(3);
    CN248_data_in(28) <= VN1529_data_out(3);
    CN248_sign_in(28) <= VN1529_sign_out(3);
    CN248_data_in(29) <= VN1597_data_out(3);
    CN248_sign_in(29) <= VN1597_sign_out(3);
    CN248_data_in(30) <= VN1658_data_out(3);
    CN248_sign_in(30) <= VN1658_sign_out(3);
    CN248_data_in(31) <= VN1785_data_out(3);
    CN248_sign_in(31) <= VN1785_sign_out(3);
    CN249_data_in(0) <= VN152_data_out(3);
    CN249_sign_in(0) <= VN152_sign_out(3);
    CN249_data_in(1) <= VN192_data_out(3);
    CN249_sign_in(1) <= VN192_sign_out(3);
    CN249_data_in(2) <= VN225_data_out(3);
    CN249_sign_in(2) <= VN225_sign_out(3);
    CN249_data_in(3) <= VN317_data_out(3);
    CN249_sign_in(3) <= VN317_sign_out(3);
    CN249_data_in(4) <= VN353_data_out(3);
    CN249_sign_in(4) <= VN353_sign_out(3);
    CN249_data_in(5) <= VN443_data_out(3);
    CN249_sign_in(5) <= VN443_sign_out(3);
    CN249_data_in(6) <= VN544_data_out(3);
    CN249_sign_in(6) <= VN544_sign_out(3);
    CN249_data_in(7) <= VN657_data_out(3);
    CN249_sign_in(7) <= VN657_sign_out(3);
    CN249_data_in(8) <= VN688_data_out(3);
    CN249_sign_in(8) <= VN688_sign_out(3);
    CN249_data_in(9) <= VN725_data_out(3);
    CN249_sign_in(9) <= VN725_sign_out(3);
    CN249_data_in(10) <= VN782_data_out(3);
    CN249_sign_in(10) <= VN782_sign_out(3);
    CN249_data_in(11) <= VN849_data_out(3);
    CN249_sign_in(11) <= VN849_sign_out(3);
    CN249_data_in(12) <= VN908_data_out(3);
    CN249_sign_in(12) <= VN908_sign_out(3);
    CN249_data_in(13) <= VN1000_data_out(3);
    CN249_sign_in(13) <= VN1000_sign_out(3);
    CN249_data_in(14) <= VN1054_data_out(3);
    CN249_sign_in(14) <= VN1054_sign_out(3);
    CN249_data_in(15) <= VN1124_data_out(3);
    CN249_sign_in(15) <= VN1124_sign_out(3);
    CN249_data_in(16) <= VN1175_data_out(3);
    CN249_sign_in(16) <= VN1175_sign_out(3);
    CN249_data_in(17) <= VN1304_data_out(3);
    CN249_sign_in(17) <= VN1304_sign_out(3);
    CN249_data_in(18) <= VN1390_data_out(3);
    CN249_sign_in(18) <= VN1390_sign_out(3);
    CN249_data_in(19) <= VN1462_data_out(3);
    CN249_sign_in(19) <= VN1462_sign_out(3);
    CN249_data_in(20) <= VN1520_data_out(3);
    CN249_sign_in(20) <= VN1520_sign_out(3);
    CN249_data_in(21) <= VN1557_data_out(3);
    CN249_sign_in(21) <= VN1557_sign_out(3);
    CN249_data_in(22) <= VN1648_data_out(3);
    CN249_sign_in(22) <= VN1648_sign_out(3);
    CN249_data_in(23) <= VN1723_data_out(3);
    CN249_sign_in(23) <= VN1723_sign_out(3);
    CN249_data_in(24) <= VN1735_data_out(3);
    CN249_sign_in(24) <= VN1735_sign_out(3);
    CN249_data_in(25) <= VN1736_data_out(3);
    CN249_sign_in(25) <= VN1736_sign_out(3);
    CN249_data_in(26) <= VN1741_data_out(3);
    CN249_sign_in(26) <= VN1741_sign_out(3);
    CN249_data_in(27) <= VN1751_data_out(3);
    CN249_sign_in(27) <= VN1751_sign_out(3);
    CN249_data_in(28) <= VN1822_data_out(3);
    CN249_sign_in(28) <= VN1822_sign_out(3);
    CN249_data_in(29) <= VN1840_data_out(3);
    CN249_sign_in(29) <= VN1840_sign_out(3);
    CN249_data_in(30) <= VN1883_data_out(3);
    CN249_sign_in(30) <= VN1883_sign_out(3);
    CN249_data_in(31) <= VN1911_data_out(3);
    CN249_sign_in(31) <= VN1911_sign_out(3);
    CN250_data_in(0) <= VN79_data_out(3);
    CN250_sign_in(0) <= VN79_sign_out(3);
    CN250_data_in(1) <= VN120_data_out(3);
    CN250_sign_in(1) <= VN120_sign_out(3);
    CN250_data_in(2) <= VN184_data_out(3);
    CN250_sign_in(2) <= VN184_sign_out(3);
    CN250_data_in(3) <= VN319_data_out(3);
    CN250_sign_in(3) <= VN319_sign_out(3);
    CN250_data_in(4) <= VN358_data_out(3);
    CN250_sign_in(4) <= VN358_sign_out(3);
    CN250_data_in(5) <= VN400_data_out(3);
    CN250_sign_in(5) <= VN400_sign_out(3);
    CN250_data_in(6) <= VN500_data_out(3);
    CN250_sign_in(6) <= VN500_sign_out(3);
    CN250_data_in(7) <= VN514_data_out(3);
    CN250_sign_in(7) <= VN514_sign_out(3);
    CN250_data_in(8) <= VN576_data_out(3);
    CN250_sign_in(8) <= VN576_sign_out(3);
    CN250_data_in(9) <= VN652_data_out(3);
    CN250_sign_in(9) <= VN652_sign_out(3);
    CN250_data_in(10) <= VN679_data_out(3);
    CN250_sign_in(10) <= VN679_sign_out(3);
    CN250_data_in(11) <= VN744_data_out(3);
    CN250_sign_in(11) <= VN744_sign_out(3);
    CN250_data_in(12) <= VN803_data_out(3);
    CN250_sign_in(12) <= VN803_sign_out(3);
    CN250_data_in(13) <= VN854_data_out(3);
    CN250_sign_in(13) <= VN854_sign_out(3);
    CN250_data_in(14) <= VN925_data_out(3);
    CN250_sign_in(14) <= VN925_sign_out(3);
    CN250_data_in(15) <= VN978_data_out(3);
    CN250_sign_in(15) <= VN978_sign_out(3);
    CN250_data_in(16) <= VN1038_data_out(3);
    CN250_sign_in(16) <= VN1038_sign_out(3);
    CN250_data_in(17) <= VN1173_data_out(3);
    CN250_sign_in(17) <= VN1173_sign_out(3);
    CN250_data_in(18) <= VN1250_data_out(3);
    CN250_sign_in(18) <= VN1250_sign_out(3);
    CN250_data_in(19) <= VN1318_data_out(3);
    CN250_sign_in(19) <= VN1318_sign_out(3);
    CN250_data_in(20) <= VN1360_data_out(3);
    CN250_sign_in(20) <= VN1360_sign_out(3);
    CN250_data_in(21) <= VN1405_data_out(3);
    CN250_sign_in(21) <= VN1405_sign_out(3);
    CN250_data_in(22) <= VN1448_data_out(3);
    CN250_sign_in(22) <= VN1448_sign_out(3);
    CN250_data_in(23) <= VN1489_data_out(3);
    CN250_sign_in(23) <= VN1489_sign_out(3);
    CN250_data_in(24) <= VN1508_data_out(3);
    CN250_sign_in(24) <= VN1508_sign_out(3);
    CN250_data_in(25) <= VN1512_data_out(3);
    CN250_sign_in(25) <= VN1512_sign_out(3);
    CN250_data_in(26) <= VN1560_data_out(3);
    CN250_sign_in(26) <= VN1560_sign_out(3);
    CN250_data_in(27) <= VN1588_data_out(3);
    CN250_sign_in(27) <= VN1588_sign_out(3);
    CN250_data_in(28) <= VN1676_data_out(3);
    CN250_sign_in(28) <= VN1676_sign_out(3);
    CN250_data_in(29) <= VN1762_data_out(3);
    CN250_sign_in(29) <= VN1762_sign_out(3);
    CN250_data_in(30) <= VN1928_data_out(3);
    CN250_sign_in(30) <= VN1928_sign_out(3);
    CN250_data_in(31) <= VN1933_data_out(3);
    CN250_sign_in(31) <= VN1933_sign_out(3);
    CN251_data_in(0) <= VN62_data_out(3);
    CN251_sign_in(0) <= VN62_sign_out(3);
    CN251_data_in(1) <= VN159_data_out(3);
    CN251_sign_in(1) <= VN159_sign_out(3);
    CN251_data_in(2) <= VN215_data_out(3);
    CN251_sign_in(2) <= VN215_sign_out(3);
    CN251_data_in(3) <= VN289_data_out(3);
    CN251_sign_in(3) <= VN289_sign_out(3);
    CN251_data_in(4) <= VN348_data_out(3);
    CN251_sign_in(4) <= VN348_sign_out(3);
    CN251_data_in(5) <= VN409_data_out(3);
    CN251_sign_in(5) <= VN409_sign_out(3);
    CN251_data_in(6) <= VN464_data_out(3);
    CN251_sign_in(6) <= VN464_sign_out(3);
    CN251_data_in(7) <= VN506_data_out(3);
    CN251_sign_in(7) <= VN506_sign_out(3);
    CN251_data_in(8) <= VN564_data_out(3);
    CN251_sign_in(8) <= VN564_sign_out(3);
    CN251_data_in(9) <= VN626_data_out(3);
    CN251_sign_in(9) <= VN626_sign_out(3);
    CN251_data_in(10) <= VN721_data_out(3);
    CN251_sign_in(10) <= VN721_sign_out(3);
    CN251_data_in(11) <= VN765_data_out(3);
    CN251_sign_in(11) <= VN765_sign_out(3);
    CN251_data_in(12) <= VN817_data_out(3);
    CN251_sign_in(12) <= VN817_sign_out(3);
    CN251_data_in(13) <= VN899_data_out(3);
    CN251_sign_in(13) <= VN899_sign_out(3);
    CN251_data_in(14) <= VN957_data_out(3);
    CN251_sign_in(14) <= VN957_sign_out(3);
    CN251_data_in(15) <= VN1015_data_out(3);
    CN251_sign_in(15) <= VN1015_sign_out(3);
    CN251_data_in(16) <= VN1081_data_out(3);
    CN251_sign_in(16) <= VN1081_sign_out(3);
    CN251_data_in(17) <= VN1135_data_out(3);
    CN251_sign_in(17) <= VN1135_sign_out(3);
    CN251_data_in(18) <= VN1187_data_out(3);
    CN251_sign_in(18) <= VN1187_sign_out(3);
    CN251_data_in(19) <= VN1221_data_out(3);
    CN251_sign_in(19) <= VN1221_sign_out(3);
    CN251_data_in(20) <= VN1247_data_out(3);
    CN251_sign_in(20) <= VN1247_sign_out(3);
    CN251_data_in(21) <= VN1294_data_out(3);
    CN251_sign_in(21) <= VN1294_sign_out(3);
    CN251_data_in(22) <= VN1346_data_out(3);
    CN251_sign_in(22) <= VN1346_sign_out(3);
    CN251_data_in(23) <= VN1409_data_out(3);
    CN251_sign_in(23) <= VN1409_sign_out(3);
    CN251_data_in(24) <= VN1477_data_out(3);
    CN251_sign_in(24) <= VN1477_sign_out(3);
    CN251_data_in(25) <= VN1501_data_out(3);
    CN251_sign_in(25) <= VN1501_sign_out(3);
    CN251_data_in(26) <= VN1570_data_out(3);
    CN251_sign_in(26) <= VN1570_sign_out(3);
    CN251_data_in(27) <= VN1644_data_out(3);
    CN251_sign_in(27) <= VN1644_sign_out(3);
    CN251_data_in(28) <= VN1665_data_out(3);
    CN251_sign_in(28) <= VN1665_sign_out(3);
    CN251_data_in(29) <= VN1722_data_out(3);
    CN251_sign_in(29) <= VN1722_sign_out(3);
    CN251_data_in(30) <= VN1793_data_out(3);
    CN251_sign_in(30) <= VN1793_sign_out(3);
    CN251_data_in(31) <= VN1859_data_out(3);
    CN251_sign_in(31) <= VN1859_sign_out(3);
    CN252_data_in(0) <= VN89_data_out(3);
    CN252_sign_in(0) <= VN89_sign_out(3);
    CN252_data_in(1) <= VN112_data_out(3);
    CN252_sign_in(1) <= VN112_sign_out(3);
    CN252_data_in(2) <= VN199_data_out(3);
    CN252_sign_in(2) <= VN199_sign_out(3);
    CN252_data_in(3) <= VN239_data_out(3);
    CN252_sign_in(3) <= VN239_sign_out(3);
    CN252_data_in(4) <= VN325_data_out(3);
    CN252_sign_in(4) <= VN325_sign_out(3);
    CN252_data_in(5) <= VN373_data_out(3);
    CN252_sign_in(5) <= VN373_sign_out(3);
    CN252_data_in(6) <= VN438_data_out(3);
    CN252_sign_in(6) <= VN438_sign_out(3);
    CN252_data_in(7) <= VN473_data_out(3);
    CN252_sign_in(7) <= VN473_sign_out(3);
    CN252_data_in(8) <= VN549_data_out(3);
    CN252_sign_in(8) <= VN549_sign_out(3);
    CN252_data_in(9) <= VN605_data_out(3);
    CN252_sign_in(9) <= VN605_sign_out(3);
    CN252_data_in(10) <= VN635_data_out(3);
    CN252_sign_in(10) <= VN635_sign_out(3);
    CN252_data_in(11) <= VN684_data_out(3);
    CN252_sign_in(11) <= VN684_sign_out(3);
    CN252_data_in(12) <= VN766_data_out(3);
    CN252_sign_in(12) <= VN766_sign_out(3);
    CN252_data_in(13) <= VN813_data_out(3);
    CN252_sign_in(13) <= VN813_sign_out(3);
    CN252_data_in(14) <= VN853_data_out(3);
    CN252_sign_in(14) <= VN853_sign_out(3);
    CN252_data_in(15) <= VN896_data_out(3);
    CN252_sign_in(15) <= VN896_sign_out(3);
    CN252_data_in(16) <= VN960_data_out(3);
    CN252_sign_in(16) <= VN960_sign_out(3);
    CN252_data_in(17) <= VN1034_data_out(3);
    CN252_sign_in(17) <= VN1034_sign_out(3);
    CN252_data_in(18) <= VN1093_data_out(3);
    CN252_sign_in(18) <= VN1093_sign_out(3);
    CN252_data_in(19) <= VN1126_data_out(3);
    CN252_sign_in(19) <= VN1126_sign_out(3);
    CN252_data_in(20) <= VN1180_data_out(3);
    CN252_sign_in(20) <= VN1180_sign_out(3);
    CN252_data_in(21) <= VN1262_data_out(3);
    CN252_sign_in(21) <= VN1262_sign_out(3);
    CN252_data_in(22) <= VN1326_data_out(3);
    CN252_sign_in(22) <= VN1326_sign_out(3);
    CN252_data_in(23) <= VN1398_data_out(3);
    CN252_sign_in(23) <= VN1398_sign_out(3);
    CN252_data_in(24) <= VN1563_data_out(3);
    CN252_sign_in(24) <= VN1563_sign_out(3);
    CN252_data_in(25) <= VN1589_data_out(3);
    CN252_sign_in(25) <= VN1589_sign_out(3);
    CN252_data_in(26) <= VN1671_data_out(3);
    CN252_sign_in(26) <= VN1671_sign_out(3);
    CN252_data_in(27) <= VN1721_data_out(3);
    CN252_sign_in(27) <= VN1721_sign_out(3);
    CN252_data_in(28) <= VN1731_data_out(3);
    CN252_sign_in(28) <= VN1731_sign_out(3);
    CN252_data_in(29) <= VN1742_data_out(3);
    CN252_sign_in(29) <= VN1742_sign_out(3);
    CN252_data_in(30) <= VN1805_data_out(3);
    CN252_sign_in(30) <= VN1805_sign_out(3);
    CN252_data_in(31) <= VN1860_data_out(3);
    CN252_sign_in(31) <= VN1860_sign_out(3);
    CN253_data_in(0) <= VN80_data_out(3);
    CN253_sign_in(0) <= VN80_sign_out(3);
    CN253_data_in(1) <= VN121_data_out(3);
    CN253_sign_in(1) <= VN121_sign_out(3);
    CN253_data_in(2) <= VN211_data_out(3);
    CN253_sign_in(2) <= VN211_sign_out(3);
    CN253_data_in(3) <= VN279_data_out(3);
    CN253_sign_in(3) <= VN279_sign_out(3);
    CN253_data_in(4) <= VN283_data_out(3);
    CN253_sign_in(4) <= VN283_sign_out(3);
    CN253_data_in(5) <= VN380_data_out(3);
    CN253_sign_in(5) <= VN380_sign_out(3);
    CN253_data_in(6) <= VN426_data_out(3);
    CN253_sign_in(6) <= VN426_sign_out(3);
    CN253_data_in(7) <= VN468_data_out(3);
    CN253_sign_in(7) <= VN468_sign_out(3);
    CN253_data_in(8) <= VN510_data_out(3);
    CN253_sign_in(8) <= VN510_sign_out(3);
    CN253_data_in(9) <= VN567_data_out(3);
    CN253_sign_in(9) <= VN567_sign_out(3);
    CN253_data_in(10) <= VN629_data_out(3);
    CN253_sign_in(10) <= VN629_sign_out(3);
    CN253_data_in(11) <= VN714_data_out(3);
    CN253_sign_in(11) <= VN714_sign_out(3);
    CN253_data_in(12) <= VN743_data_out(3);
    CN253_sign_in(12) <= VN743_sign_out(3);
    CN253_data_in(13) <= VN778_data_out(3);
    CN253_sign_in(13) <= VN778_sign_out(3);
    CN253_data_in(14) <= VN847_data_out(3);
    CN253_sign_in(14) <= VN847_sign_out(3);
    CN253_data_in(15) <= VN912_data_out(3);
    CN253_sign_in(15) <= VN912_sign_out(3);
    CN253_data_in(16) <= VN944_data_out(3);
    CN253_sign_in(16) <= VN944_sign_out(3);
    CN253_data_in(17) <= VN1007_data_out(3);
    CN253_sign_in(17) <= VN1007_sign_out(3);
    CN253_data_in(18) <= VN1060_data_out(3);
    CN253_sign_in(18) <= VN1060_sign_out(3);
    CN253_data_in(19) <= VN1114_data_out(3);
    CN253_sign_in(19) <= VN1114_sign_out(3);
    CN253_data_in(20) <= VN1211_data_out(3);
    CN253_sign_in(20) <= VN1211_sign_out(3);
    CN253_data_in(21) <= VN1255_data_out(3);
    CN253_sign_in(21) <= VN1255_sign_out(3);
    CN253_data_in(22) <= VN1296_data_out(3);
    CN253_sign_in(22) <= VN1296_sign_out(3);
    CN253_data_in(23) <= VN1342_data_out(3);
    CN253_sign_in(23) <= VN1342_sign_out(3);
    CN253_data_in(24) <= VN1541_data_out(3);
    CN253_sign_in(24) <= VN1541_sign_out(3);
    CN253_data_in(25) <= VN1567_data_out(3);
    CN253_sign_in(25) <= VN1567_sign_out(3);
    CN253_data_in(26) <= VN1599_data_out(3);
    CN253_sign_in(26) <= VN1599_sign_out(3);
    CN253_data_in(27) <= VN1635_data_out(3);
    CN253_sign_in(27) <= VN1635_sign_out(3);
    CN253_data_in(28) <= VN1681_data_out(3);
    CN253_sign_in(28) <= VN1681_sign_out(3);
    CN253_data_in(29) <= VN1719_data_out(3);
    CN253_sign_in(29) <= VN1719_sign_out(3);
    CN253_data_in(30) <= VN1768_data_out(3);
    CN253_sign_in(30) <= VN1768_sign_out(3);
    CN253_data_in(31) <= VN1861_data_out(3);
    CN253_sign_in(31) <= VN1861_sign_out(3);
    CN254_data_in(0) <= VN67_data_out(3);
    CN254_sign_in(0) <= VN67_sign_out(3);
    CN254_data_in(1) <= VN222_data_out(3);
    CN254_sign_in(1) <= VN222_sign_out(3);
    CN254_data_in(2) <= VN238_data_out(3);
    CN254_sign_in(2) <= VN238_sign_out(3);
    CN254_data_in(3) <= VN290_data_out(3);
    CN254_sign_in(3) <= VN290_sign_out(3);
    CN254_data_in(4) <= VN362_data_out(3);
    CN254_sign_in(4) <= VN362_sign_out(3);
    CN254_data_in(5) <= VN412_data_out(3);
    CN254_sign_in(5) <= VN412_sign_out(3);
    CN254_data_in(6) <= VN474_data_out(3);
    CN254_sign_in(6) <= VN474_sign_out(3);
    CN254_data_in(7) <= VN540_data_out(3);
    CN254_sign_in(7) <= VN540_sign_out(3);
    CN254_data_in(8) <= VN586_data_out(3);
    CN254_sign_in(8) <= VN586_sign_out(3);
    CN254_data_in(9) <= VN632_data_out(3);
    CN254_sign_in(9) <= VN632_sign_out(3);
    CN254_data_in(10) <= VN712_data_out(3);
    CN254_sign_in(10) <= VN712_sign_out(3);
    CN254_data_in(11) <= VN735_data_out(3);
    CN254_sign_in(11) <= VN735_sign_out(3);
    CN254_data_in(12) <= VN798_data_out(3);
    CN254_sign_in(12) <= VN798_sign_out(3);
    CN254_data_in(13) <= VN884_data_out(3);
    CN254_sign_in(13) <= VN884_sign_out(3);
    CN254_data_in(14) <= VN905_data_out(3);
    CN254_sign_in(14) <= VN905_sign_out(3);
    CN254_data_in(15) <= VN979_data_out(3);
    CN254_sign_in(15) <= VN979_sign_out(3);
    CN254_data_in(16) <= VN1047_data_out(3);
    CN254_sign_in(16) <= VN1047_sign_out(3);
    CN254_data_in(17) <= VN1107_data_out(3);
    CN254_sign_in(17) <= VN1107_sign_out(3);
    CN254_data_in(18) <= VN1131_data_out(3);
    CN254_sign_in(18) <= VN1131_sign_out(3);
    CN254_data_in(19) <= VN1232_data_out(3);
    CN254_sign_in(19) <= VN1232_sign_out(3);
    CN254_data_in(20) <= VN1306_data_out(3);
    CN254_sign_in(20) <= VN1306_sign_out(3);
    CN254_data_in(21) <= VN1369_data_out(3);
    CN254_sign_in(21) <= VN1369_sign_out(3);
    CN254_data_in(22) <= VN1417_data_out(3);
    CN254_sign_in(22) <= VN1417_sign_out(3);
    CN254_data_in(23) <= VN1443_data_out(3);
    CN254_sign_in(23) <= VN1443_sign_out(3);
    CN254_data_in(24) <= VN1456_data_out(3);
    CN254_sign_in(24) <= VN1456_sign_out(3);
    CN254_data_in(25) <= VN1493_data_out(3);
    CN254_sign_in(25) <= VN1493_sign_out(3);
    CN254_data_in(26) <= VN1516_data_out(3);
    CN254_sign_in(26) <= VN1516_sign_out(3);
    CN254_data_in(27) <= VN1720_data_out(3);
    CN254_sign_in(27) <= VN1720_sign_out(3);
    CN254_data_in(28) <= VN1733_data_out(3);
    CN254_sign_in(28) <= VN1733_sign_out(3);
    CN254_data_in(29) <= VN1754_data_out(3);
    CN254_sign_in(29) <= VN1754_sign_out(3);
    CN254_data_in(30) <= VN1923_data_out(3);
    CN254_sign_in(30) <= VN1923_sign_out(3);
    CN254_data_in(31) <= VN1926_data_out(3);
    CN254_sign_in(31) <= VN1926_sign_out(3);
    CN255_data_in(0) <= VN52_data_out(3);
    CN255_sign_in(0) <= VN52_sign_out(3);
    CN255_data_in(1) <= VN86_data_out(3);
    CN255_sign_in(1) <= VN86_sign_out(3);
    CN255_data_in(2) <= VN167_data_out(3);
    CN255_sign_in(2) <= VN167_sign_out(3);
    CN255_data_in(3) <= VN195_data_out(3);
    CN255_sign_in(3) <= VN195_sign_out(3);
    CN255_data_in(4) <= VN233_data_out(3);
    CN255_sign_in(4) <= VN233_sign_out(3);
    CN255_data_in(5) <= VN318_data_out(3);
    CN255_sign_in(5) <= VN318_sign_out(3);
    CN255_data_in(6) <= VN364_data_out(3);
    CN255_sign_in(6) <= VN364_sign_out(3);
    CN255_data_in(7) <= VN429_data_out(3);
    CN255_sign_in(7) <= VN429_sign_out(3);
    CN255_data_in(8) <= VN537_data_out(3);
    CN255_sign_in(8) <= VN537_sign_out(3);
    CN255_data_in(9) <= VN594_data_out(3);
    CN255_sign_in(9) <= VN594_sign_out(3);
    CN255_data_in(10) <= VN672_data_out(3);
    CN255_sign_in(10) <= VN672_sign_out(3);
    CN255_data_in(11) <= VN751_data_out(3);
    CN255_sign_in(11) <= VN751_sign_out(3);
    CN255_data_in(12) <= VN799_data_out(3);
    CN255_sign_in(12) <= VN799_sign_out(3);
    CN255_data_in(13) <= VN934_data_out(3);
    CN255_sign_in(13) <= VN934_sign_out(3);
    CN255_data_in(14) <= VN1017_data_out(3);
    CN255_sign_in(14) <= VN1017_sign_out(3);
    CN255_data_in(15) <= VN1077_data_out(3);
    CN255_sign_in(15) <= VN1077_sign_out(3);
    CN255_data_in(16) <= VN1110_data_out(3);
    CN255_sign_in(16) <= VN1110_sign_out(3);
    CN255_data_in(17) <= VN1163_data_out(3);
    CN255_sign_in(17) <= VN1163_sign_out(3);
    CN255_data_in(18) <= VN1214_data_out(3);
    CN255_sign_in(18) <= VN1214_sign_out(3);
    CN255_data_in(19) <= VN1432_data_out(3);
    CN255_sign_in(19) <= VN1432_sign_out(3);
    CN255_data_in(20) <= VN1465_data_out(3);
    CN255_sign_in(20) <= VN1465_sign_out(3);
    CN255_data_in(21) <= VN1538_data_out(3);
    CN255_sign_in(21) <= VN1538_sign_out(3);
    CN255_data_in(22) <= VN1691_data_out(3);
    CN255_sign_in(22) <= VN1691_sign_out(3);
    CN255_data_in(23) <= VN1787_data_out(3);
    CN255_sign_in(23) <= VN1787_sign_out(3);
    CN255_data_in(24) <= VN1836_data_out(3);
    CN255_sign_in(24) <= VN1836_sign_out(3);
    CN255_data_in(25) <= VN1879_data_out(3);
    CN255_sign_in(25) <= VN1879_sign_out(3);
    CN255_data_in(26) <= VN1897_data_out(3);
    CN255_sign_in(26) <= VN1897_sign_out(3);
    CN255_data_in(27) <= VN1906_data_out(3);
    CN255_sign_in(27) <= VN1906_sign_out(3);
    CN255_data_in(28) <= VN1929_data_out(3);
    CN255_sign_in(28) <= VN1929_sign_out(3);
    CN255_data_in(29) <= VN1936_data_out(3);
    CN255_sign_in(29) <= VN1936_sign_out(3);
    CN255_data_in(30) <= VN1961_data_out(3);
    CN255_sign_in(30) <= VN1961_sign_out(3);
    CN255_data_in(31) <= VN1979_data_out(3);
    CN255_sign_in(31) <= VN1979_sign_out(3);
    CN256_data_in(0) <= VN53_data_out(4);
    CN256_sign_in(0) <= VN53_sign_out(4);
    CN256_data_in(1) <= VN106_data_out(4);
    CN256_sign_in(1) <= VN106_sign_out(4);
    CN256_data_in(2) <= VN127_data_out(4);
    CN256_sign_in(2) <= VN127_sign_out(4);
    CN256_data_in(3) <= VN242_data_out(4);
    CN256_sign_in(3) <= VN242_sign_out(4);
    CN256_data_in(4) <= VN296_data_out(4);
    CN256_sign_in(4) <= VN296_sign_out(4);
    CN256_data_in(5) <= VN339_data_out(4);
    CN256_sign_in(5) <= VN339_sign_out(4);
    CN256_data_in(6) <= VN455_data_out(4);
    CN256_sign_in(6) <= VN455_sign_out(4);
    CN256_data_in(7) <= VN532_data_out(4);
    CN256_sign_in(7) <= VN532_sign_out(4);
    CN256_data_in(8) <= VN638_data_out(4);
    CN256_sign_in(8) <= VN638_sign_out(4);
    CN256_data_in(9) <= VN708_data_out(4);
    CN256_sign_in(9) <= VN708_sign_out(4);
    CN256_data_in(10) <= VN760_data_out(4);
    CN256_sign_in(10) <= VN760_sign_out(4);
    CN256_data_in(11) <= VN793_data_out(4);
    CN256_sign_in(11) <= VN793_sign_out(4);
    CN256_data_in(12) <= VN891_data_out(4);
    CN256_sign_in(12) <= VN891_sign_out(4);
    CN256_data_in(13) <= VN1000_data_out(4);
    CN256_sign_in(13) <= VN1000_sign_out(4);
    CN256_data_in(14) <= VN1035_data_out(4);
    CN256_sign_in(14) <= VN1035_sign_out(4);
    CN256_data_in(15) <= VN1071_data_out(4);
    CN256_sign_in(15) <= VN1071_sign_out(4);
    CN256_data_in(16) <= VN1155_data_out(4);
    CN256_sign_in(16) <= VN1155_sign_out(4);
    CN256_data_in(17) <= VN1242_data_out(4);
    CN256_sign_in(17) <= VN1242_sign_out(4);
    CN256_data_in(18) <= VN1285_data_out(4);
    CN256_sign_in(18) <= VN1285_sign_out(4);
    CN256_data_in(19) <= VN1343_data_out(4);
    CN256_sign_in(19) <= VN1343_sign_out(4);
    CN256_data_in(20) <= VN1414_data_out(4);
    CN256_sign_in(20) <= VN1414_sign_out(4);
    CN256_data_in(21) <= VN1454_data_out(4);
    CN256_sign_in(21) <= VN1454_sign_out(4);
    CN256_data_in(22) <= VN1517_data_out(4);
    CN256_sign_in(22) <= VN1517_sign_out(4);
    CN256_data_in(23) <= VN1747_data_out(4);
    CN256_sign_in(23) <= VN1747_sign_out(4);
    CN256_data_in(24) <= VN1780_data_out(4);
    CN256_sign_in(24) <= VN1780_sign_out(4);
    CN256_data_in(25) <= VN1846_data_out(4);
    CN256_sign_in(25) <= VN1846_sign_out(4);
    CN256_data_in(26) <= VN1929_data_out(4);
    CN256_sign_in(26) <= VN1929_sign_out(4);
    CN256_data_in(27) <= VN1959_data_out(4);
    CN256_sign_in(27) <= VN1959_sign_out(4);
    CN256_data_in(28) <= VN1962_data_out(4);
    CN256_sign_in(28) <= VN1962_sign_out(4);
    CN256_data_in(29) <= VN1990_data_out(4);
    CN256_sign_in(29) <= VN1990_sign_out(4);
    CN256_data_in(30) <= VN1995_data_out(4);
    CN256_sign_in(30) <= VN1995_sign_out(4);
    CN256_data_in(31) <= VN1997_data_out(4);
    CN256_sign_in(31) <= VN1997_sign_out(4);
    CN257_data_in(0) <= VN51_data_out(4);
    CN257_sign_in(0) <= VN51_sign_out(4);
    CN257_data_in(1) <= VN85_data_out(4);
    CN257_sign_in(1) <= VN85_sign_out(4);
    CN257_data_in(2) <= VN166_data_out(4);
    CN257_sign_in(2) <= VN166_sign_out(4);
    CN257_data_in(3) <= VN194_data_out(4);
    CN257_sign_in(3) <= VN194_sign_out(4);
    CN257_data_in(4) <= VN232_data_out(4);
    CN257_sign_in(4) <= VN232_sign_out(4);
    CN257_data_in(5) <= VN317_data_out(4);
    CN257_sign_in(5) <= VN317_sign_out(4);
    CN257_data_in(6) <= VN363_data_out(4);
    CN257_sign_in(6) <= VN363_sign_out(4);
    CN257_data_in(7) <= VN428_data_out(4);
    CN257_sign_in(7) <= VN428_sign_out(4);
    CN257_data_in(8) <= VN463_data_out(4);
    CN257_sign_in(8) <= VN463_sign_out(4);
    CN257_data_in(9) <= VN536_data_out(4);
    CN257_sign_in(9) <= VN536_sign_out(4);
    CN257_data_in(10) <= VN593_data_out(4);
    CN257_sign_in(10) <= VN593_sign_out(4);
    CN257_data_in(11) <= VN624_data_out(4);
    CN257_sign_in(11) <= VN624_sign_out(4);
    CN257_data_in(12) <= VN671_data_out(4);
    CN257_sign_in(12) <= VN671_sign_out(4);
    CN257_data_in(13) <= VN750_data_out(4);
    CN257_sign_in(13) <= VN750_sign_out(4);
    CN257_data_in(14) <= VN798_data_out(4);
    CN257_sign_in(14) <= VN798_sign_out(4);
    CN257_data_in(15) <= VN835_data_out(4);
    CN257_sign_in(15) <= VN835_sign_out(4);
    CN257_data_in(16) <= VN933_data_out(4);
    CN257_sign_in(16) <= VN933_sign_out(4);
    CN257_data_in(17) <= VN999_data_out(4);
    CN257_sign_in(17) <= VN999_sign_out(4);
    CN257_data_in(18) <= VN1016_data_out(4);
    CN257_sign_in(18) <= VN1016_sign_out(4);
    CN257_data_in(19) <= VN1076_data_out(4);
    CN257_sign_in(19) <= VN1076_sign_out(4);
    CN257_data_in(20) <= VN1108_data_out(4);
    CN257_sign_in(20) <= VN1108_sign_out(4);
    CN257_data_in(21) <= VN1162_data_out(4);
    CN257_sign_in(21) <= VN1162_sign_out(4);
    CN257_data_in(22) <= VN1213_data_out(4);
    CN257_sign_in(22) <= VN1213_sign_out(4);
    CN257_data_in(23) <= VN1240_data_out(4);
    CN257_sign_in(23) <= VN1240_sign_out(4);
    CN257_data_in(24) <= VN1303_data_out(4);
    CN257_sign_in(24) <= VN1303_sign_out(4);
    CN257_data_in(25) <= VN1354_data_out(4);
    CN257_sign_in(25) <= VN1354_sign_out(4);
    CN257_data_in(26) <= VN1431_data_out(4);
    CN257_sign_in(26) <= VN1431_sign_out(4);
    CN257_data_in(27) <= VN1464_data_out(4);
    CN257_sign_in(27) <= VN1464_sign_out(4);
    CN257_data_in(28) <= VN1484_data_out(4);
    CN257_sign_in(28) <= VN1484_sign_out(4);
    CN257_data_in(29) <= VN1652_data_out(4);
    CN257_sign_in(29) <= VN1652_sign_out(4);
    CN257_data_in(30) <= VN1690_data_out(4);
    CN257_sign_in(30) <= VN1690_sign_out(4);
    CN257_data_in(31) <= VN1786_data_out(4);
    CN257_sign_in(31) <= VN1786_sign_out(4);
    CN258_data_in(0) <= VN50_data_out(4);
    CN258_sign_in(0) <= VN50_sign_out(4);
    CN258_data_in(1) <= VN57_data_out(4);
    CN258_sign_in(1) <= VN57_sign_out(4);
    CN258_data_in(2) <= VN331_data_out(4);
    CN258_sign_in(2) <= VN331_sign_out(4);
    CN258_data_in(3) <= VN553_data_out(4);
    CN258_sign_in(3) <= VN553_sign_out(4);
    CN258_data_in(4) <= VN589_data_out(4);
    CN258_sign_in(4) <= VN589_sign_out(4);
    CN258_data_in(5) <= VN657_data_out(4);
    CN258_sign_in(5) <= VN657_sign_out(4);
    CN258_data_in(6) <= VN718_data_out(4);
    CN258_sign_in(6) <= VN718_sign_out(4);
    CN258_data_in(7) <= VN755_data_out(4);
    CN258_sign_in(7) <= VN755_sign_out(4);
    CN258_data_in(8) <= VN829_data_out(4);
    CN258_sign_in(8) <= VN829_sign_out(4);
    CN258_data_in(9) <= VN857_data_out(4);
    CN258_sign_in(9) <= VN857_sign_out(4);
    CN258_data_in(10) <= VN943_data_out(4);
    CN258_sign_in(10) <= VN943_sign_out(4);
    CN258_data_in(11) <= VN968_data_out(4);
    CN258_sign_in(11) <= VN968_sign_out(4);
    CN258_data_in(12) <= VN1077_data_out(4);
    CN258_sign_in(12) <= VN1077_sign_out(4);
    CN258_data_in(13) <= VN1159_data_out(4);
    CN258_sign_in(13) <= VN1159_sign_out(4);
    CN258_data_in(14) <= VN1215_data_out(4);
    CN258_sign_in(14) <= VN1215_sign_out(4);
    CN258_data_in(15) <= VN1222_data_out(4);
    CN258_sign_in(15) <= VN1222_sign_out(4);
    CN258_data_in(16) <= VN1320_data_out(4);
    CN258_sign_in(16) <= VN1320_sign_out(4);
    CN258_data_in(17) <= VN1378_data_out(4);
    CN258_sign_in(17) <= VN1378_sign_out(4);
    CN258_data_in(18) <= VN1547_data_out(4);
    CN258_sign_in(18) <= VN1547_sign_out(4);
    CN258_data_in(19) <= VN1574_data_out(4);
    CN258_sign_in(19) <= VN1574_sign_out(4);
    CN258_data_in(20) <= VN1632_data_out(4);
    CN258_sign_in(20) <= VN1632_sign_out(4);
    CN258_data_in(21) <= VN1682_data_out(4);
    CN258_sign_in(21) <= VN1682_sign_out(4);
    CN258_data_in(22) <= VN1770_data_out(4);
    CN258_sign_in(22) <= VN1770_sign_out(4);
    CN258_data_in(23) <= VN1778_data_out(4);
    CN258_sign_in(23) <= VN1778_sign_out(4);
    CN258_data_in(24) <= VN1801_data_out(4);
    CN258_sign_in(24) <= VN1801_sign_out(4);
    CN258_data_in(25) <= VN1834_data_out(4);
    CN258_sign_in(25) <= VN1834_sign_out(4);
    CN258_data_in(26) <= VN1884_data_out(4);
    CN258_sign_in(26) <= VN1884_sign_out(4);
    CN258_data_in(27) <= VN1901_data_out(4);
    CN258_sign_in(27) <= VN1901_sign_out(4);
    CN258_data_in(28) <= VN1921_data_out(4);
    CN258_sign_in(28) <= VN1921_sign_out(4);
    CN258_data_in(29) <= VN1922_data_out(4);
    CN258_sign_in(29) <= VN1922_sign_out(4);
    CN258_data_in(30) <= VN1945_data_out(4);
    CN258_sign_in(30) <= VN1945_sign_out(4);
    CN258_data_in(31) <= VN1954_data_out(4);
    CN258_sign_in(31) <= VN1954_sign_out(4);
    CN259_data_in(0) <= VN54_data_out(4);
    CN259_sign_in(0) <= VN54_sign_out(4);
    CN259_data_in(1) <= VN114_data_out(4);
    CN259_sign_in(1) <= VN114_sign_out(4);
    CN259_data_in(2) <= VN274_data_out(4);
    CN259_sign_in(2) <= VN274_sign_out(4);
    CN259_data_in(3) <= VN303_data_out(4);
    CN259_sign_in(3) <= VN303_sign_out(4);
    CN259_data_in(4) <= VN370_data_out(4);
    CN259_sign_in(4) <= VN370_sign_out(4);
    CN259_data_in(5) <= VN491_data_out(4);
    CN259_sign_in(5) <= VN491_sign_out(4);
    CN259_data_in(6) <= VN545_data_out(4);
    CN259_sign_in(6) <= VN545_sign_out(4);
    CN259_data_in(7) <= VN594_data_out(4);
    CN259_sign_in(7) <= VN594_sign_out(4);
    CN259_data_in(8) <= VN641_data_out(4);
    CN259_sign_in(8) <= VN641_sign_out(4);
    CN259_data_in(9) <= VN694_data_out(4);
    CN259_sign_in(9) <= VN694_sign_out(4);
    CN259_data_in(10) <= VN822_data_out(4);
    CN259_sign_in(10) <= VN822_sign_out(4);
    CN259_data_in(11) <= VN856_data_out(4);
    CN259_sign_in(11) <= VN856_sign_out(4);
    CN259_data_in(12) <= VN937_data_out(4);
    CN259_sign_in(12) <= VN937_sign_out(4);
    CN259_data_in(13) <= VN952_data_out(4);
    CN259_sign_in(13) <= VN952_sign_out(4);
    CN259_data_in(14) <= VN1051_data_out(4);
    CN259_sign_in(14) <= VN1051_sign_out(4);
    CN259_data_in(15) <= VN1105_data_out(4);
    CN259_sign_in(15) <= VN1105_sign_out(4);
    CN259_data_in(16) <= VN1117_data_out(4);
    CN259_sign_in(16) <= VN1117_sign_out(4);
    CN259_data_in(17) <= VN1207_data_out(4);
    CN259_sign_in(17) <= VN1207_sign_out(4);
    CN259_data_in(18) <= VN1218_data_out(4);
    CN259_sign_in(18) <= VN1218_sign_out(4);
    CN259_data_in(19) <= VN1238_data_out(4);
    CN259_sign_in(19) <= VN1238_sign_out(4);
    CN259_data_in(20) <= VN1289_data_out(4);
    CN259_sign_in(20) <= VN1289_sign_out(4);
    CN259_data_in(21) <= VN1499_data_out(4);
    CN259_sign_in(21) <= VN1499_sign_out(4);
    CN259_data_in(22) <= VN1584_data_out(4);
    CN259_sign_in(22) <= VN1584_sign_out(4);
    CN259_data_in(23) <= VN1615_data_out(4);
    CN259_sign_in(23) <= VN1615_sign_out(4);
    CN259_data_in(24) <= VN1728_data_out(4);
    CN259_sign_in(24) <= VN1728_sign_out(4);
    CN259_data_in(25) <= VN1735_data_out(4);
    CN259_sign_in(25) <= VN1735_sign_out(4);
    CN259_data_in(26) <= VN1738_data_out(4);
    CN259_sign_in(26) <= VN1738_sign_out(4);
    CN259_data_in(27) <= VN1833_data_out(4);
    CN259_sign_in(27) <= VN1833_sign_out(4);
    CN259_data_in(28) <= VN1844_data_out(4);
    CN259_sign_in(28) <= VN1844_sign_out(4);
    CN259_data_in(29) <= VN1970_data_out(4);
    CN259_sign_in(29) <= VN1970_sign_out(4);
    CN259_data_in(30) <= VN1981_data_out(4);
    CN259_sign_in(30) <= VN1981_sign_out(4);
    CN259_data_in(31) <= VN1986_data_out(4);
    CN259_sign_in(31) <= VN1986_sign_out(4);
    CN260_data_in(0) <= VN49_data_out(4);
    CN260_sign_in(0) <= VN49_sign_out(4);
    CN260_data_in(1) <= VN71_data_out(4);
    CN260_sign_in(1) <= VN71_sign_out(4);
    CN260_data_in(2) <= VN138_data_out(4);
    CN260_sign_in(2) <= VN138_sign_out(4);
    CN260_data_in(3) <= VN186_data_out(4);
    CN260_sign_in(3) <= VN186_sign_out(4);
    CN260_data_in(4) <= VN243_data_out(4);
    CN260_sign_in(4) <= VN243_sign_out(4);
    CN260_data_in(5) <= VN383_data_out(4);
    CN260_sign_in(5) <= VN383_sign_out(4);
    CN260_data_in(6) <= VN396_data_out(4);
    CN260_sign_in(6) <= VN396_sign_out(4);
    CN260_data_in(7) <= VN584_data_out(4);
    CN260_sign_in(7) <= VN584_sign_out(4);
    CN260_data_in(8) <= VN754_data_out(4);
    CN260_sign_in(8) <= VN754_sign_out(4);
    CN260_data_in(9) <= VN833_data_out(4);
    CN260_sign_in(9) <= VN833_sign_out(4);
    CN260_data_in(10) <= VN941_data_out(4);
    CN260_sign_in(10) <= VN941_sign_out(4);
    CN260_data_in(11) <= VN980_data_out(4);
    CN260_sign_in(11) <= VN980_sign_out(4);
    CN260_data_in(12) <= VN1013_data_out(4);
    CN260_sign_in(12) <= VN1013_sign_out(4);
    CN260_data_in(13) <= VN1187_data_out(4);
    CN260_sign_in(13) <= VN1187_sign_out(4);
    CN260_data_in(14) <= VN1228_data_out(4);
    CN260_sign_in(14) <= VN1228_sign_out(4);
    CN260_data_in(15) <= VN1290_data_out(4);
    CN260_sign_in(15) <= VN1290_sign_out(4);
    CN260_data_in(16) <= VN1399_data_out(4);
    CN260_sign_in(16) <= VN1399_sign_out(4);
    CN260_data_in(17) <= VN1437_data_out(4);
    CN260_sign_in(17) <= VN1437_sign_out(4);
    CN260_data_in(18) <= VN1463_data_out(4);
    CN260_sign_in(18) <= VN1463_sign_out(4);
    CN260_data_in(19) <= VN1618_data_out(4);
    CN260_sign_in(19) <= VN1618_sign_out(4);
    CN260_data_in(20) <= VN1718_data_out(4);
    CN260_sign_in(20) <= VN1718_sign_out(4);
    CN260_data_in(21) <= VN1765_data_out(4);
    CN260_sign_in(21) <= VN1765_sign_out(4);
    CN260_data_in(22) <= VN1771_data_out(4);
    CN260_sign_in(22) <= VN1771_sign_out(4);
    CN260_data_in(23) <= VN1822_data_out(4);
    CN260_sign_in(23) <= VN1822_sign_out(4);
    CN260_data_in(24) <= VN1857_data_out(4);
    CN260_sign_in(24) <= VN1857_sign_out(4);
    CN260_data_in(25) <= VN1943_data_out(4);
    CN260_sign_in(25) <= VN1943_sign_out(4);
    CN260_data_in(26) <= VN1963_data_out(4);
    CN260_sign_in(26) <= VN1963_sign_out(4);
    CN260_data_in(27) <= VN1988_data_out(4);
    CN260_sign_in(27) <= VN1988_sign_out(4);
    CN260_data_in(28) <= VN2015_data_out(4);
    CN260_sign_in(28) <= VN2015_sign_out(4);
    CN260_data_in(29) <= VN2020_data_out(4);
    CN260_sign_in(29) <= VN2020_sign_out(4);
    CN260_data_in(30) <= VN2023_data_out(4);
    CN260_sign_in(30) <= VN2023_sign_out(4);
    CN260_data_in(31) <= VN2030_data_out(4);
    CN260_sign_in(31) <= VN2030_sign_out(4);
    CN261_data_in(0) <= VN48_data_out(4);
    CN261_sign_in(0) <= VN48_sign_out(4);
    CN261_data_in(1) <= VN63_data_out(4);
    CN261_sign_in(1) <= VN63_sign_out(4);
    CN261_data_in(2) <= VN152_data_out(4);
    CN261_sign_in(2) <= VN152_sign_out(4);
    CN261_data_in(3) <= VN204_data_out(4);
    CN261_sign_in(3) <= VN204_sign_out(4);
    CN261_data_in(4) <= VN305_data_out(4);
    CN261_sign_in(4) <= VN305_sign_out(4);
    CN261_data_in(5) <= VN333_data_out(4);
    CN261_sign_in(5) <= VN333_sign_out(4);
    CN261_data_in(6) <= VN401_data_out(4);
    CN261_sign_in(6) <= VN401_sign_out(4);
    CN261_data_in(7) <= VN477_data_out(4);
    CN261_sign_in(7) <= VN477_sign_out(4);
    CN261_data_in(8) <= VN528_data_out(4);
    CN261_sign_in(8) <= VN528_sign_out(4);
    CN261_data_in(9) <= VN607_data_out(4);
    CN261_sign_in(9) <= VN607_sign_out(4);
    CN261_data_in(10) <= VN698_data_out(4);
    CN261_sign_in(10) <= VN698_sign_out(4);
    CN261_data_in(11) <= VN777_data_out(4);
    CN261_sign_in(11) <= VN777_sign_out(4);
    CN261_data_in(12) <= VN789_data_out(4);
    CN261_sign_in(12) <= VN789_sign_out(4);
    CN261_data_in(13) <= VN868_data_out(4);
    CN261_sign_in(13) <= VN868_sign_out(4);
    CN261_data_in(14) <= VN970_data_out(4);
    CN261_sign_in(14) <= VN970_sign_out(4);
    CN261_data_in(15) <= VN1042_data_out(4);
    CN261_sign_in(15) <= VN1042_sign_out(4);
    CN261_data_in(16) <= VN1062_data_out(4);
    CN261_sign_in(16) <= VN1062_sign_out(4);
    CN261_data_in(17) <= VN1141_data_out(4);
    CN261_sign_in(17) <= VN1141_sign_out(4);
    CN261_data_in(18) <= VN1171_data_out(4);
    CN261_sign_in(18) <= VN1171_sign_out(4);
    CN261_data_in(19) <= VN1262_data_out(4);
    CN261_sign_in(19) <= VN1262_sign_out(4);
    CN261_data_in(20) <= VN1319_data_out(4);
    CN261_sign_in(20) <= VN1319_sign_out(4);
    CN261_data_in(21) <= VN1375_data_out(4);
    CN261_sign_in(21) <= VN1375_sign_out(4);
    CN261_data_in(22) <= VN1493_data_out(4);
    CN261_sign_in(22) <= VN1493_sign_out(4);
    CN261_data_in(23) <= VN1549_data_out(4);
    CN261_sign_in(23) <= VN1549_sign_out(4);
    CN261_data_in(24) <= VN1570_data_out(4);
    CN261_sign_in(24) <= VN1570_sign_out(4);
    CN261_data_in(25) <= VN1603_data_out(4);
    CN261_sign_in(25) <= VN1603_sign_out(4);
    CN261_data_in(26) <= VN1672_data_out(4);
    CN261_sign_in(26) <= VN1672_sign_out(4);
    CN261_data_in(27) <= VN1704_data_out(4);
    CN261_sign_in(27) <= VN1704_sign_out(4);
    CN261_data_in(28) <= VN1761_data_out(4);
    CN261_sign_in(28) <= VN1761_sign_out(4);
    CN261_data_in(29) <= VN1842_data_out(4);
    CN261_sign_in(29) <= VN1842_sign_out(4);
    CN261_data_in(30) <= VN1874_data_out(4);
    CN261_sign_in(30) <= VN1874_sign_out(4);
    CN261_data_in(31) <= VN1891_data_out(4);
    CN261_sign_in(31) <= VN1891_sign_out(4);
    CN262_data_in(0) <= VN47_data_out(4);
    CN262_sign_in(0) <= VN47_sign_out(4);
    CN262_data_in(1) <= VN95_data_out(4);
    CN262_sign_in(1) <= VN95_sign_out(4);
    CN262_data_in(2) <= VN149_data_out(4);
    CN262_sign_in(2) <= VN149_sign_out(4);
    CN262_data_in(3) <= VN212_data_out(4);
    CN262_sign_in(3) <= VN212_sign_out(4);
    CN262_data_in(4) <= VN319_data_out(4);
    CN262_sign_in(4) <= VN319_sign_out(4);
    CN262_data_in(5) <= VN362_data_out(4);
    CN262_sign_in(5) <= VN362_sign_out(4);
    CN262_data_in(6) <= VN392_data_out(4);
    CN262_sign_in(6) <= VN392_sign_out(4);
    CN262_data_in(7) <= VN503_data_out(4);
    CN262_sign_in(7) <= VN503_sign_out(4);
    CN262_data_in(8) <= VN522_data_out(4);
    CN262_sign_in(8) <= VN522_sign_out(4);
    CN262_data_in(9) <= VN613_data_out(4);
    CN262_sign_in(9) <= VN613_sign_out(4);
    CN262_data_in(10) <= VN635_data_out(4);
    CN262_sign_in(10) <= VN635_sign_out(4);
    CN262_data_in(11) <= VN702_data_out(4);
    CN262_sign_in(11) <= VN702_sign_out(4);
    CN262_data_in(12) <= VN731_data_out(4);
    CN262_sign_in(12) <= VN731_sign_out(4);
    CN262_data_in(13) <= VN830_data_out(4);
    CN262_sign_in(13) <= VN830_sign_out(4);
    CN262_data_in(14) <= VN871_data_out(4);
    CN262_sign_in(14) <= VN871_sign_out(4);
    CN262_data_in(15) <= VN912_data_out(4);
    CN262_sign_in(15) <= VN912_sign_out(4);
    CN262_data_in(16) <= VN957_data_out(4);
    CN262_sign_in(16) <= VN957_sign_out(4);
    CN262_data_in(17) <= VN1039_data_out(4);
    CN262_sign_in(17) <= VN1039_sign_out(4);
    CN262_data_in(18) <= VN1067_data_out(4);
    CN262_sign_in(18) <= VN1067_sign_out(4);
    CN262_data_in(19) <= VN1152_data_out(4);
    CN262_sign_in(19) <= VN1152_sign_out(4);
    CN262_data_in(20) <= VN1183_data_out(4);
    CN262_sign_in(20) <= VN1183_sign_out(4);
    CN262_data_in(21) <= VN1245_data_out(4);
    CN262_sign_in(21) <= VN1245_sign_out(4);
    CN262_data_in(22) <= VN1311_data_out(4);
    CN262_sign_in(22) <= VN1311_sign_out(4);
    CN262_data_in(23) <= VN1350_data_out(4);
    CN262_sign_in(23) <= VN1350_sign_out(4);
    CN262_data_in(24) <= VN1402_data_out(4);
    CN262_sign_in(24) <= VN1402_sign_out(4);
    CN262_data_in(25) <= VN1480_data_out(4);
    CN262_sign_in(25) <= VN1480_sign_out(4);
    CN262_data_in(26) <= VN1500_data_out(4);
    CN262_sign_in(26) <= VN1500_sign_out(4);
    CN262_data_in(27) <= VN1559_data_out(4);
    CN262_sign_in(27) <= VN1559_sign_out(4);
    CN262_data_in(28) <= VN1633_data_out(4);
    CN262_sign_in(28) <= VN1633_sign_out(4);
    CN262_data_in(29) <= VN1700_data_out(4);
    CN262_sign_in(29) <= VN1700_sign_out(4);
    CN262_data_in(30) <= VN1807_data_out(4);
    CN262_sign_in(30) <= VN1807_sign_out(4);
    CN262_data_in(31) <= VN1862_data_out(4);
    CN262_sign_in(31) <= VN1862_sign_out(4);
    CN263_data_in(0) <= VN46_data_out(4);
    CN263_sign_in(0) <= VN46_sign_out(4);
    CN263_data_in(1) <= VN104_data_out(4);
    CN263_sign_in(1) <= VN104_sign_out(4);
    CN263_data_in(2) <= VN169_data_out(4);
    CN263_sign_in(2) <= VN169_sign_out(4);
    CN263_data_in(3) <= VN207_data_out(4);
    CN263_sign_in(3) <= VN207_sign_out(4);
    CN263_data_in(4) <= VN253_data_out(4);
    CN263_sign_in(4) <= VN253_sign_out(4);
    CN263_data_in(5) <= VN315_data_out(4);
    CN263_sign_in(5) <= VN315_sign_out(4);
    CN263_data_in(6) <= VN378_data_out(4);
    CN263_sign_in(6) <= VN378_sign_out(4);
    CN263_data_in(7) <= VN414_data_out(4);
    CN263_sign_in(7) <= VN414_sign_out(4);
    CN263_data_in(8) <= VN525_data_out(4);
    CN263_sign_in(8) <= VN525_sign_out(4);
    CN263_data_in(9) <= VN598_data_out(4);
    CN263_sign_in(9) <= VN598_sign_out(4);
    CN263_data_in(10) <= VN691_data_out(4);
    CN263_sign_in(10) <= VN691_sign_out(4);
    CN263_data_in(11) <= VN738_data_out(4);
    CN263_sign_in(11) <= VN738_sign_out(4);
    CN263_data_in(12) <= VN788_data_out(4);
    CN263_sign_in(12) <= VN788_sign_out(4);
    CN263_data_in(13) <= VN858_data_out(4);
    CN263_sign_in(13) <= VN858_sign_out(4);
    CN263_data_in(14) <= VN894_data_out(4);
    CN263_sign_in(14) <= VN894_sign_out(4);
    CN263_data_in(15) <= VN976_data_out(4);
    CN263_sign_in(15) <= VN976_sign_out(4);
    CN263_data_in(16) <= VN1056_data_out(4);
    CN263_sign_in(16) <= VN1056_sign_out(4);
    CN263_data_in(17) <= VN1145_data_out(4);
    CN263_sign_in(17) <= VN1145_sign_out(4);
    CN263_data_in(18) <= VN1257_data_out(4);
    CN263_sign_in(18) <= VN1257_sign_out(4);
    CN263_data_in(19) <= VN1347_data_out(4);
    CN263_sign_in(19) <= VN1347_sign_out(4);
    CN263_data_in(20) <= VN1492_data_out(4);
    CN263_sign_in(20) <= VN1492_sign_out(4);
    CN263_data_in(21) <= VN1509_data_out(4);
    CN263_sign_in(21) <= VN1509_sign_out(4);
    CN263_data_in(22) <= VN1526_data_out(4);
    CN263_sign_in(22) <= VN1526_sign_out(4);
    CN263_data_in(23) <= VN1554_data_out(4);
    CN263_sign_in(23) <= VN1554_sign_out(4);
    CN263_data_in(24) <= VN1576_data_out(4);
    CN263_sign_in(24) <= VN1576_sign_out(4);
    CN263_data_in(25) <= VN1673_data_out(4);
    CN263_sign_in(25) <= VN1673_sign_out(4);
    CN263_data_in(26) <= VN1743_data_out(4);
    CN263_sign_in(26) <= VN1743_sign_out(4);
    CN263_data_in(27) <= VN1840_data_out(4);
    CN263_sign_in(27) <= VN1840_sign_out(4);
    CN263_data_in(28) <= VN1841_data_out(4);
    CN263_sign_in(28) <= VN1841_sign_out(4);
    CN263_data_in(29) <= VN1905_data_out(4);
    CN263_sign_in(29) <= VN1905_sign_out(4);
    CN263_data_in(30) <= VN1971_data_out(4);
    CN263_sign_in(30) <= VN1971_sign_out(4);
    CN263_data_in(31) <= VN1978_data_out(4);
    CN263_sign_in(31) <= VN1978_sign_out(4);
    CN264_data_in(0) <= VN45_data_out(4);
    CN264_sign_in(0) <= VN45_sign_out(4);
    CN264_data_in(1) <= VN98_data_out(4);
    CN264_sign_in(1) <= VN98_sign_out(4);
    CN264_data_in(2) <= VN132_data_out(4);
    CN264_sign_in(2) <= VN132_sign_out(4);
    CN264_data_in(3) <= VN213_data_out(4);
    CN264_sign_in(3) <= VN213_sign_out(4);
    CN264_data_in(4) <= VN256_data_out(4);
    CN264_sign_in(4) <= VN256_sign_out(4);
    CN264_data_in(5) <= VN281_data_out(4);
    CN264_sign_in(5) <= VN281_sign_out(4);
    CN264_data_in(6) <= VN349_data_out(4);
    CN264_sign_in(6) <= VN349_sign_out(4);
    CN264_data_in(7) <= VN421_data_out(4);
    CN264_sign_in(7) <= VN421_sign_out(4);
    CN264_data_in(8) <= VN495_data_out(4);
    CN264_sign_in(8) <= VN495_sign_out(4);
    CN264_data_in(9) <= VN600_data_out(4);
    CN264_sign_in(9) <= VN600_sign_out(4);
    CN264_data_in(10) <= VN666_data_out(4);
    CN264_sign_in(10) <= VN666_sign_out(4);
    CN264_data_in(11) <= VN672_data_out(4);
    CN264_sign_in(11) <= VN672_sign_out(4);
    CN264_data_in(12) <= VN761_data_out(4);
    CN264_sign_in(12) <= VN761_sign_out(4);
    CN264_data_in(13) <= VN783_data_out(4);
    CN264_sign_in(13) <= VN783_sign_out(4);
    CN264_data_in(14) <= VN834_data_out(4);
    CN264_sign_in(14) <= VN834_sign_out(4);
    CN264_data_in(15) <= VN908_data_out(4);
    CN264_sign_in(15) <= VN908_sign_out(4);
    CN264_data_in(16) <= VN948_data_out(4);
    CN264_sign_in(16) <= VN948_sign_out(4);
    CN264_data_in(17) <= VN1048_data_out(4);
    CN264_sign_in(17) <= VN1048_sign_out(4);
    CN264_data_in(18) <= VN1066_data_out(4);
    CN264_sign_in(18) <= VN1066_sign_out(4);
    CN264_data_in(19) <= VN1149_data_out(4);
    CN264_sign_in(19) <= VN1149_sign_out(4);
    CN264_data_in(20) <= VN1269_data_out(4);
    CN264_sign_in(20) <= VN1269_sign_out(4);
    CN264_data_in(21) <= VN1279_data_out(4);
    CN264_sign_in(21) <= VN1279_sign_out(4);
    CN264_data_in(22) <= VN1362_data_out(4);
    CN264_sign_in(22) <= VN1362_sign_out(4);
    CN264_data_in(23) <= VN1516_data_out(4);
    CN264_sign_in(23) <= VN1516_sign_out(4);
    CN264_data_in(24) <= VN1531_data_out(4);
    CN264_sign_in(24) <= VN1531_sign_out(4);
    CN264_data_in(25) <= VN1561_data_out(4);
    CN264_sign_in(25) <= VN1561_sign_out(4);
    CN264_data_in(26) <= VN1607_data_out(4);
    CN264_sign_in(26) <= VN1607_sign_out(4);
    CN264_data_in(27) <= VN1693_data_out(4);
    CN264_sign_in(27) <= VN1693_sign_out(4);
    CN264_data_in(28) <= VN1753_data_out(4);
    CN264_sign_in(28) <= VN1753_sign_out(4);
    CN264_data_in(29) <= VN1802_data_out(4);
    CN264_sign_in(29) <= VN1802_sign_out(4);
    CN264_data_in(30) <= VN1806_data_out(4);
    CN264_sign_in(30) <= VN1806_sign_out(4);
    CN264_data_in(31) <= VN1863_data_out(4);
    CN264_sign_in(31) <= VN1863_sign_out(4);
    CN265_data_in(0) <= VN44_data_out(4);
    CN265_sign_in(0) <= VN44_sign_out(4);
    CN265_data_in(1) <= VN133_data_out(4);
    CN265_sign_in(1) <= VN133_sign_out(4);
    CN265_data_in(2) <= VN203_data_out(4);
    CN265_sign_in(2) <= VN203_sign_out(4);
    CN265_data_in(3) <= VN244_data_out(4);
    CN265_sign_in(3) <= VN244_sign_out(4);
    CN265_data_in(4) <= VN386_data_out(4);
    CN265_sign_in(4) <= VN386_sign_out(4);
    CN265_data_in(5) <= VN405_data_out(4);
    CN265_sign_in(5) <= VN405_sign_out(4);
    CN265_data_in(6) <= VN504_data_out(4);
    CN265_sign_in(6) <= VN504_sign_out(4);
    CN265_data_in(7) <= VN627_data_out(4);
    CN265_sign_in(7) <= VN627_sign_out(4);
    CN265_data_in(8) <= VN759_data_out(4);
    CN265_sign_in(8) <= VN759_sign_out(4);
    CN265_data_in(9) <= VN855_data_out(4);
    CN265_sign_in(9) <= VN855_sign_out(4);
    CN265_data_in(10) <= VN918_data_out(4);
    CN265_sign_in(10) <= VN918_sign_out(4);
    CN265_data_in(11) <= VN945_data_out(4);
    CN265_sign_in(11) <= VN945_sign_out(4);
    CN265_data_in(12) <= VN1023_data_out(4);
    CN265_sign_in(12) <= VN1023_sign_out(4);
    CN265_data_in(13) <= VN1209_data_out(4);
    CN265_sign_in(13) <= VN1209_sign_out(4);
    CN265_data_in(14) <= VN1355_data_out(4);
    CN265_sign_in(14) <= VN1355_sign_out(4);
    CN265_data_in(15) <= VN1385_data_out(4);
    CN265_sign_in(15) <= VN1385_sign_out(4);
    CN265_data_in(16) <= VN1445_data_out(4);
    CN265_sign_in(16) <= VN1445_sign_out(4);
    CN265_data_in(17) <= VN1486_data_out(4);
    CN265_sign_in(17) <= VN1486_sign_out(4);
    CN265_data_in(18) <= VN1532_data_out(4);
    CN265_sign_in(18) <= VN1532_sign_out(4);
    CN265_data_in(19) <= VN1612_data_out(4);
    CN265_sign_in(19) <= VN1612_sign_out(4);
    CN265_data_in(20) <= VN1757_data_out(4);
    CN265_sign_in(20) <= VN1757_sign_out(4);
    CN265_data_in(21) <= VN1845_data_out(4);
    CN265_sign_in(21) <= VN1845_sign_out(4);
    CN265_data_in(22) <= VN1858_data_out(4);
    CN265_sign_in(22) <= VN1858_sign_out(4);
    CN265_data_in(23) <= VN1888_data_out(4);
    CN265_sign_in(23) <= VN1888_sign_out(4);
    CN265_data_in(24) <= VN1906_data_out(4);
    CN265_sign_in(24) <= VN1906_sign_out(4);
    CN265_data_in(25) <= VN1915_data_out(4);
    CN265_sign_in(25) <= VN1915_sign_out(4);
    CN265_data_in(26) <= VN1992_data_out(4);
    CN265_sign_in(26) <= VN1992_sign_out(4);
    CN265_data_in(27) <= VN1993_data_out(4);
    CN265_sign_in(27) <= VN1993_sign_out(4);
    CN265_data_in(28) <= VN2028_data_out(4);
    CN265_sign_in(28) <= VN2028_sign_out(4);
    CN265_data_in(29) <= VN2032_data_out(4);
    CN265_sign_in(29) <= VN2032_sign_out(4);
    CN265_data_in(30) <= VN2043_data_out(4);
    CN265_sign_in(30) <= VN2043_sign_out(4);
    CN265_data_in(31) <= VN2046_data_out(4);
    CN265_sign_in(31) <= VN2046_sign_out(4);
    CN266_data_in(0) <= VN43_data_out(4);
    CN266_sign_in(0) <= VN43_sign_out(4);
    CN266_data_in(1) <= VN168_data_out(4);
    CN266_sign_in(1) <= VN168_sign_out(4);
    CN266_data_in(2) <= VN173_data_out(4);
    CN266_sign_in(2) <= VN173_sign_out(4);
    CN266_data_in(3) <= VN273_data_out(4);
    CN266_sign_in(3) <= VN273_sign_out(4);
    CN266_data_in(4) <= VN300_data_out(4);
    CN266_sign_in(4) <= VN300_sign_out(4);
    CN266_data_in(5) <= VN535_data_out(4);
    CN266_sign_in(5) <= VN535_sign_out(4);
    CN266_data_in(6) <= VN605_data_out(4);
    CN266_sign_in(6) <= VN605_sign_out(4);
    CN266_data_in(7) <= VN647_data_out(4);
    CN266_sign_in(7) <= VN647_sign_out(4);
    CN266_data_in(8) <= VN721_data_out(4);
    CN266_sign_in(8) <= VN721_sign_out(4);
    CN266_data_in(9) <= VN880_data_out(4);
    CN266_sign_in(9) <= VN880_sign_out(4);
    CN266_data_in(10) <= VN888_data_out(4);
    CN266_sign_in(10) <= VN888_sign_out(4);
    CN266_data_in(11) <= VN962_data_out(4);
    CN266_sign_in(11) <= VN962_sign_out(4);
    CN266_data_in(12) <= VN1032_data_out(4);
    CN266_sign_in(12) <= VN1032_sign_out(4);
    CN266_data_in(13) <= VN1095_data_out(4);
    CN266_sign_in(13) <= VN1095_sign_out(4);
    CN266_data_in(14) <= VN1118_data_out(4);
    CN266_sign_in(14) <= VN1118_sign_out(4);
    CN266_data_in(15) <= VN1195_data_out(4);
    CN266_sign_in(15) <= VN1195_sign_out(4);
    CN266_data_in(16) <= VN1230_data_out(4);
    CN266_sign_in(16) <= VN1230_sign_out(4);
    CN266_data_in(17) <= VN1429_data_out(4);
    CN266_sign_in(17) <= VN1429_sign_out(4);
    CN266_data_in(18) <= VN1478_data_out(4);
    CN266_sign_in(18) <= VN1478_sign_out(4);
    CN266_data_in(19) <= VN1530_data_out(4);
    CN266_sign_in(19) <= VN1530_sign_out(4);
    CN266_data_in(20) <= VN1534_data_out(4);
    CN266_sign_in(20) <= VN1534_sign_out(4);
    CN266_data_in(21) <= VN1539_data_out(4);
    CN266_sign_in(21) <= VN1539_sign_out(4);
    CN266_data_in(22) <= VN1635_data_out(4);
    CN266_sign_in(22) <= VN1635_sign_out(4);
    CN266_data_in(23) <= VN1725_data_out(4);
    CN266_sign_in(23) <= VN1725_sign_out(4);
    CN266_data_in(24) <= VN1815_data_out(4);
    CN266_sign_in(24) <= VN1815_sign_out(4);
    CN266_data_in(25) <= VN1824_data_out(4);
    CN266_sign_in(25) <= VN1824_sign_out(4);
    CN266_data_in(26) <= VN1827_data_out(4);
    CN266_sign_in(26) <= VN1827_sign_out(4);
    CN266_data_in(27) <= VN1898_data_out(4);
    CN266_sign_in(27) <= VN1898_sign_out(4);
    CN266_data_in(28) <= VN1908_data_out(4);
    CN266_sign_in(28) <= VN1908_sign_out(4);
    CN266_data_in(29) <= VN1965_data_out(4);
    CN266_sign_in(29) <= VN1965_sign_out(4);
    CN266_data_in(30) <= VN1996_data_out(4);
    CN266_sign_in(30) <= VN1996_sign_out(4);
    CN266_data_in(31) <= VN2006_data_out(4);
    CN266_sign_in(31) <= VN2006_sign_out(4);
    CN267_data_in(0) <= VN42_data_out(4);
    CN267_sign_in(0) <= VN42_sign_out(4);
    CN267_data_in(1) <= VN72_data_out(4);
    CN267_sign_in(1) <= VN72_sign_out(4);
    CN267_data_in(2) <= VN159_data_out(4);
    CN267_sign_in(2) <= VN159_sign_out(4);
    CN267_data_in(3) <= VN180_data_out(4);
    CN267_sign_in(3) <= VN180_sign_out(4);
    CN267_data_in(4) <= VN241_data_out(4);
    CN267_sign_in(4) <= VN241_sign_out(4);
    CN267_data_in(5) <= VN280_data_out(4);
    CN267_sign_in(5) <= VN280_sign_out(4);
    CN267_data_in(6) <= VN364_data_out(4);
    CN267_sign_in(6) <= VN364_sign_out(4);
    CN267_data_in(7) <= VN432_data_out(4);
    CN267_sign_in(7) <= VN432_sign_out(4);
    CN267_data_in(8) <= VN490_data_out(4);
    CN267_sign_in(8) <= VN490_sign_out(4);
    CN267_data_in(9) <= VN549_data_out(4);
    CN267_sign_in(9) <= VN549_sign_out(4);
    CN267_data_in(10) <= VN562_data_out(4);
    CN267_sign_in(10) <= VN562_sign_out(4);
    CN267_data_in(11) <= VN654_data_out(4);
    CN267_sign_in(11) <= VN654_sign_out(4);
    CN267_data_in(12) <= VN677_data_out(4);
    CN267_sign_in(12) <= VN677_sign_out(4);
    CN267_data_in(13) <= VN794_data_out(4);
    CN267_sign_in(13) <= VN794_sign_out(4);
    CN267_data_in(14) <= VN866_data_out(4);
    CN267_sign_in(14) <= VN866_sign_out(4);
    CN267_data_in(15) <= VN932_data_out(4);
    CN267_sign_in(15) <= VN932_sign_out(4);
    CN267_data_in(16) <= VN954_data_out(4);
    CN267_sign_in(16) <= VN954_sign_out(4);
    CN267_data_in(17) <= VN1026_data_out(4);
    CN267_sign_in(17) <= VN1026_sign_out(4);
    CN267_data_in(18) <= VN1101_data_out(4);
    CN267_sign_in(18) <= VN1101_sign_out(4);
    CN267_data_in(19) <= VN1158_data_out(4);
    CN267_sign_in(19) <= VN1158_sign_out(4);
    CN267_data_in(20) <= VN1212_data_out(4);
    CN267_sign_in(20) <= VN1212_sign_out(4);
    CN267_data_in(21) <= VN1272_data_out(4);
    CN267_sign_in(21) <= VN1272_sign_out(4);
    CN267_data_in(22) <= VN1327_data_out(4);
    CN267_sign_in(22) <= VN1327_sign_out(4);
    CN267_data_in(23) <= VN1339_data_out(4);
    CN267_sign_in(23) <= VN1339_sign_out(4);
    CN267_data_in(24) <= VN1390_data_out(4);
    CN267_sign_in(24) <= VN1390_sign_out(4);
    CN267_data_in(25) <= VN1421_data_out(4);
    CN267_sign_in(25) <= VN1421_sign_out(4);
    CN267_data_in(26) <= VN1601_data_out(4);
    CN267_sign_in(26) <= VN1601_sign_out(4);
    CN267_data_in(27) <= VN1628_data_out(4);
    CN267_sign_in(27) <= VN1628_sign_out(4);
    CN267_data_in(28) <= VN1677_data_out(4);
    CN267_sign_in(28) <= VN1677_sign_out(4);
    CN267_data_in(29) <= VN1692_data_out(4);
    CN267_sign_in(29) <= VN1692_sign_out(4);
    CN267_data_in(30) <= VN1724_data_out(4);
    CN267_sign_in(30) <= VN1724_sign_out(4);
    CN267_data_in(31) <= VN1864_data_out(4);
    CN267_sign_in(31) <= VN1864_sign_out(4);
    CN268_data_in(0) <= VN41_data_out(4);
    CN268_sign_in(0) <= VN41_sign_out(4);
    CN268_data_in(1) <= VN109_data_out(4);
    CN268_sign_in(1) <= VN109_sign_out(4);
    CN268_data_in(2) <= VN118_data_out(4);
    CN268_sign_in(2) <= VN118_sign_out(4);
    CN268_data_in(3) <= VN216_data_out(4);
    CN268_sign_in(3) <= VN216_sign_out(4);
    CN268_data_in(4) <= VN266_data_out(4);
    CN268_sign_in(4) <= VN266_sign_out(4);
    CN268_data_in(5) <= VN325_data_out(4);
    CN268_sign_in(5) <= VN325_sign_out(4);
    CN268_data_in(6) <= VN360_data_out(4);
    CN268_sign_in(6) <= VN360_sign_out(4);
    CN268_data_in(7) <= VN412_data_out(4);
    CN268_sign_in(7) <= VN412_sign_out(4);
    CN268_data_in(8) <= VN464_data_out(4);
    CN268_sign_in(8) <= VN464_sign_out(4);
    CN268_data_in(9) <= VN559_data_out(4);
    CN268_sign_in(9) <= VN559_sign_out(4);
    CN268_data_in(10) <= VN570_data_out(4);
    CN268_sign_in(10) <= VN570_sign_out(4);
    CN268_data_in(11) <= VN652_data_out(4);
    CN268_sign_in(11) <= VN652_sign_out(4);
    CN268_data_in(12) <= VN705_data_out(4);
    CN268_sign_in(12) <= VN705_sign_out(4);
    CN268_data_in(13) <= VN775_data_out(4);
    CN268_sign_in(13) <= VN775_sign_out(4);
    CN268_data_in(14) <= VN792_data_out(4);
    CN268_sign_in(14) <= VN792_sign_out(4);
    CN268_data_in(15) <= VN921_data_out(4);
    CN268_sign_in(15) <= VN921_sign_out(4);
    CN268_data_in(16) <= VN987_data_out(4);
    CN268_sign_in(16) <= VN987_sign_out(4);
    CN268_data_in(17) <= VN1029_data_out(4);
    CN268_sign_in(17) <= VN1029_sign_out(4);
    CN268_data_in(18) <= VN1072_data_out(4);
    CN268_sign_in(18) <= VN1072_sign_out(4);
    CN268_data_in(19) <= VN1114_data_out(4);
    CN268_sign_in(19) <= VN1114_sign_out(4);
    CN268_data_in(20) <= VN1176_data_out(4);
    CN268_sign_in(20) <= VN1176_sign_out(4);
    CN268_data_in(21) <= VN1233_data_out(4);
    CN268_sign_in(21) <= VN1233_sign_out(4);
    CN268_data_in(22) <= VN1309_data_out(4);
    CN268_sign_in(22) <= VN1309_sign_out(4);
    CN268_data_in(23) <= VN1335_data_out(4);
    CN268_sign_in(23) <= VN1335_sign_out(4);
    CN268_data_in(24) <= VN1391_data_out(4);
    CN268_sign_in(24) <= VN1391_sign_out(4);
    CN268_data_in(25) <= VN1430_data_out(4);
    CN268_sign_in(25) <= VN1430_sign_out(4);
    CN268_data_in(26) <= VN1449_data_out(4);
    CN268_sign_in(26) <= VN1449_sign_out(4);
    CN268_data_in(27) <= VN1459_data_out(4);
    CN268_sign_in(27) <= VN1459_sign_out(4);
    CN268_data_in(28) <= VN1616_data_out(4);
    CN268_sign_in(28) <= VN1616_sign_out(4);
    CN268_data_in(29) <= VN1678_data_out(4);
    CN268_sign_in(29) <= VN1678_sign_out(4);
    CN268_data_in(30) <= VN1711_data_out(4);
    CN268_sign_in(30) <= VN1711_sign_out(4);
    CN268_data_in(31) <= VN1787_data_out(4);
    CN268_sign_in(31) <= VN1787_sign_out(4);
    CN269_data_in(0) <= VN67_data_out(4);
    CN269_sign_in(0) <= VN67_sign_out(4);
    CN269_data_in(1) <= VN122_data_out(4);
    CN269_sign_in(1) <= VN122_sign_out(4);
    CN269_data_in(2) <= VN218_data_out(4);
    CN269_sign_in(2) <= VN218_sign_out(4);
    CN269_data_in(3) <= VN250_data_out(4);
    CN269_sign_in(3) <= VN250_sign_out(4);
    CN269_data_in(4) <= VN287_data_out(4);
    CN269_sign_in(4) <= VN287_sign_out(4);
    CN269_data_in(5) <= VN381_data_out(4);
    CN269_sign_in(5) <= VN381_sign_out(4);
    CN269_data_in(6) <= VN424_data_out(4);
    CN269_sign_in(6) <= VN424_sign_out(4);
    CN269_data_in(7) <= VN498_data_out(4);
    CN269_sign_in(7) <= VN498_sign_out(4);
    CN269_data_in(8) <= VN529_data_out(4);
    CN269_sign_in(8) <= VN529_sign_out(4);
    CN269_data_in(9) <= VN599_data_out(4);
    CN269_sign_in(9) <= VN599_sign_out(4);
    CN269_data_in(10) <= VN655_data_out(4);
    CN269_sign_in(10) <= VN655_sign_out(4);
    CN269_data_in(11) <= VN693_data_out(4);
    CN269_sign_in(11) <= VN693_sign_out(4);
    CN269_data_in(12) <= VN762_data_out(4);
    CN269_sign_in(12) <= VN762_sign_out(4);
    CN269_data_in(13) <= VN825_data_out(4);
    CN269_sign_in(13) <= VN825_sign_out(4);
    CN269_data_in(14) <= VN882_data_out(4);
    CN269_sign_in(14) <= VN882_sign_out(4);
    CN269_data_in(15) <= VN935_data_out(4);
    CN269_sign_in(15) <= VN935_sign_out(4);
    CN269_data_in(16) <= VN997_data_out(4);
    CN269_sign_in(16) <= VN997_sign_out(4);
    CN269_data_in(17) <= VN1070_data_out(4);
    CN269_sign_in(17) <= VN1070_sign_out(4);
    CN269_data_in(18) <= VN1124_data_out(4);
    CN269_sign_in(18) <= VN1124_sign_out(4);
    CN269_data_in(19) <= VN1185_data_out(4);
    CN269_sign_in(19) <= VN1185_sign_out(4);
    CN269_data_in(20) <= VN1251_data_out(4);
    CN269_sign_in(20) <= VN1251_sign_out(4);
    CN269_data_in(21) <= VN1315_data_out(4);
    CN269_sign_in(21) <= VN1315_sign_out(4);
    CN269_data_in(22) <= VN1337_data_out(4);
    CN269_sign_in(22) <= VN1337_sign_out(4);
    CN269_data_in(23) <= VN1384_data_out(4);
    CN269_sign_in(23) <= VN1384_sign_out(4);
    CN269_data_in(24) <= VN1395_data_out(4);
    CN269_sign_in(24) <= VN1395_sign_out(4);
    CN269_data_in(25) <= VN1444_data_out(4);
    CN269_sign_in(25) <= VN1444_sign_out(4);
    CN269_data_in(26) <= VN1580_data_out(4);
    CN269_sign_in(26) <= VN1580_sign_out(4);
    CN269_data_in(27) <= VN1631_data_out(4);
    CN269_sign_in(27) <= VN1631_sign_out(4);
    CN269_data_in(28) <= VN1656_data_out(4);
    CN269_sign_in(28) <= VN1656_sign_out(4);
    CN269_data_in(29) <= VN1739_data_out(4);
    CN269_sign_in(29) <= VN1739_sign_out(4);
    CN269_data_in(30) <= VN1810_data_out(4);
    CN269_sign_in(30) <= VN1810_sign_out(4);
    CN269_data_in(31) <= VN1892_data_out(4);
    CN269_sign_in(31) <= VN1892_sign_out(4);
    CN270_data_in(0) <= VN40_data_out(4);
    CN270_sign_in(0) <= VN40_sign_out(4);
    CN270_data_in(1) <= VN79_data_out(4);
    CN270_sign_in(1) <= VN79_sign_out(4);
    CN270_data_in(2) <= VN170_data_out(4);
    CN270_sign_in(2) <= VN170_sign_out(4);
    CN270_data_in(3) <= VN190_data_out(4);
    CN270_sign_in(3) <= VN190_sign_out(4);
    CN270_data_in(4) <= VN275_data_out(4);
    CN270_sign_in(4) <= VN275_sign_out(4);
    CN270_data_in(5) <= VN292_data_out(4);
    CN270_sign_in(5) <= VN292_sign_out(4);
    CN270_data_in(6) <= VN344_data_out(4);
    CN270_sign_in(6) <= VN344_sign_out(4);
    CN270_data_in(7) <= VN433_data_out(4);
    CN270_sign_in(7) <= VN433_sign_out(4);
    CN270_data_in(8) <= VN466_data_out(4);
    CN270_sign_in(8) <= VN466_sign_out(4);
    CN270_data_in(9) <= VN518_data_out(4);
    CN270_sign_in(9) <= VN518_sign_out(4);
    CN270_data_in(10) <= VN612_data_out(4);
    CN270_sign_in(10) <= VN612_sign_out(4);
    CN270_data_in(11) <= VN646_data_out(4);
    CN270_sign_in(11) <= VN646_sign_out(4);
    CN270_data_in(12) <= VN680_data_out(4);
    CN270_sign_in(12) <= VN680_sign_out(4);
    CN270_data_in(13) <= VN737_data_out(4);
    CN270_sign_in(13) <= VN737_sign_out(4);
    CN270_data_in(14) <= VN805_data_out(4);
    CN270_sign_in(14) <= VN805_sign_out(4);
    CN270_data_in(15) <= VN869_data_out(4);
    CN270_sign_in(15) <= VN869_sign_out(4);
    CN270_data_in(16) <= VN900_data_out(4);
    CN270_sign_in(16) <= VN900_sign_out(4);
    CN270_data_in(17) <= VN991_data_out(4);
    CN270_sign_in(17) <= VN991_sign_out(4);
    CN270_data_in(18) <= VN1057_data_out(4);
    CN270_sign_in(18) <= VN1057_sign_out(4);
    CN270_data_in(19) <= VN1100_data_out(4);
    CN270_sign_in(19) <= VN1100_sign_out(4);
    CN270_data_in(20) <= VN1153_data_out(4);
    CN270_sign_in(20) <= VN1153_sign_out(4);
    CN270_data_in(21) <= VN1180_data_out(4);
    CN270_sign_in(21) <= VN1180_sign_out(4);
    CN270_data_in(22) <= VN1259_data_out(4);
    CN270_sign_in(22) <= VN1259_sign_out(4);
    CN270_data_in(23) <= VN1277_data_out(4);
    CN270_sign_in(23) <= VN1277_sign_out(4);
    CN270_data_in(24) <= VN1383_data_out(4);
    CN270_sign_in(24) <= VN1383_sign_out(4);
    CN270_data_in(25) <= VN1442_data_out(4);
    CN270_sign_in(25) <= VN1442_sign_out(4);
    CN270_data_in(26) <= VN1542_data_out(4);
    CN270_sign_in(26) <= VN1542_sign_out(4);
    CN270_data_in(27) <= VN1579_data_out(4);
    CN270_sign_in(27) <= VN1579_sign_out(4);
    CN270_data_in(28) <= VN1609_data_out(4);
    CN270_sign_in(28) <= VN1609_sign_out(4);
    CN270_data_in(29) <= VN1683_data_out(4);
    CN270_sign_in(29) <= VN1683_sign_out(4);
    CN270_data_in(30) <= VN1707_data_out(4);
    CN270_sign_in(30) <= VN1707_sign_out(4);
    CN270_data_in(31) <= VN1788_data_out(4);
    CN270_sign_in(31) <= VN1788_sign_out(4);
    CN271_data_in(0) <= VN39_data_out(4);
    CN271_sign_in(0) <= VN39_sign_out(4);
    CN271_data_in(1) <= VN105_data_out(4);
    CN271_sign_in(1) <= VN105_sign_out(4);
    CN271_data_in(2) <= VN171_data_out(4);
    CN271_sign_in(2) <= VN171_sign_out(4);
    CN271_data_in(3) <= VN268_data_out(4);
    CN271_sign_in(3) <= VN268_sign_out(4);
    CN271_data_in(4) <= VN332_data_out(4);
    CN271_sign_in(4) <= VN332_sign_out(4);
    CN271_data_in(5) <= VN345_data_out(4);
    CN271_sign_in(5) <= VN345_sign_out(4);
    CN271_data_in(6) <= VN406_data_out(4);
    CN271_sign_in(6) <= VN406_sign_out(4);
    CN271_data_in(7) <= VN478_data_out(4);
    CN271_sign_in(7) <= VN478_sign_out(4);
    CN271_data_in(8) <= VN507_data_out(4);
    CN271_sign_in(8) <= VN507_sign_out(4);
    CN271_data_in(9) <= VN586_data_out(4);
    CN271_sign_in(9) <= VN586_sign_out(4);
    CN271_data_in(10) <= VN696_data_out(4);
    CN271_sign_in(10) <= VN696_sign_out(4);
    CN271_data_in(11) <= VN758_data_out(4);
    CN271_sign_in(11) <= VN758_sign_out(4);
    CN271_data_in(12) <= VN807_data_out(4);
    CN271_sign_in(12) <= VN807_sign_out(4);
    CN271_data_in(13) <= VN832_data_out(4);
    CN271_sign_in(13) <= VN832_sign_out(4);
    CN271_data_in(14) <= VN994_data_out(4);
    CN271_sign_in(14) <= VN994_sign_out(4);
    CN271_data_in(15) <= VN1038_data_out(4);
    CN271_sign_in(15) <= VN1038_sign_out(4);
    CN271_data_in(16) <= VN1083_data_out(4);
    CN271_sign_in(16) <= VN1083_sign_out(4);
    CN271_data_in(17) <= VN1140_data_out(4);
    CN271_sign_in(17) <= VN1140_sign_out(4);
    CN271_data_in(18) <= VN1255_data_out(4);
    CN271_sign_in(18) <= VN1255_sign_out(4);
    CN271_data_in(19) <= VN1330_data_out(4);
    CN271_sign_in(19) <= VN1330_sign_out(4);
    CN271_data_in(20) <= VN1363_data_out(4);
    CN271_sign_in(20) <= VN1363_sign_out(4);
    CN271_data_in(21) <= VN1472_data_out(4);
    CN271_sign_in(21) <= VN1472_sign_out(4);
    CN271_data_in(22) <= VN1544_data_out(4);
    CN271_sign_in(22) <= VN1544_sign_out(4);
    CN271_data_in(23) <= VN1606_data_out(4);
    CN271_sign_in(23) <= VN1606_sign_out(4);
    CN271_data_in(24) <= VN1608_data_out(4);
    CN271_sign_in(24) <= VN1608_sign_out(4);
    CN271_data_in(25) <= VN1803_data_out(4);
    CN271_sign_in(25) <= VN1803_sign_out(4);
    CN271_data_in(26) <= VN1849_data_out(4);
    CN271_sign_in(26) <= VN1849_sign_out(4);
    CN271_data_in(27) <= VN1852_data_out(4);
    CN271_sign_in(27) <= VN1852_sign_out(4);
    CN271_data_in(28) <= VN1895_data_out(4);
    CN271_sign_in(28) <= VN1895_sign_out(4);
    CN271_data_in(29) <= VN1911_data_out(4);
    CN271_sign_in(29) <= VN1911_sign_out(4);
    CN271_data_in(30) <= VN1941_data_out(4);
    CN271_sign_in(30) <= VN1941_sign_out(4);
    CN271_data_in(31) <= VN1948_data_out(4);
    CN271_sign_in(31) <= VN1948_sign_out(4);
    CN272_data_in(0) <= VN38_data_out(4);
    CN272_sign_in(0) <= VN38_sign_out(4);
    CN272_data_in(1) <= VN94_data_out(4);
    CN272_sign_in(1) <= VN94_sign_out(4);
    CN272_data_in(2) <= VN116_data_out(4);
    CN272_sign_in(2) <= VN116_sign_out(4);
    CN272_data_in(3) <= VN184_data_out(4);
    CN272_sign_in(3) <= VN184_sign_out(4);
    CN272_data_in(4) <= VN254_data_out(4);
    CN272_sign_in(4) <= VN254_sign_out(4);
    CN272_data_in(5) <= VN291_data_out(4);
    CN272_sign_in(5) <= VN291_sign_out(4);
    CN272_data_in(6) <= VN380_data_out(4);
    CN272_sign_in(6) <= VN380_sign_out(4);
    CN272_data_in(7) <= VN420_data_out(4);
    CN272_sign_in(7) <= VN420_sign_out(4);
    CN272_data_in(8) <= VN476_data_out(4);
    CN272_sign_in(8) <= VN476_sign_out(4);
    CN272_data_in(9) <= VN520_data_out(4);
    CN272_sign_in(9) <= VN520_sign_out(4);
    CN272_data_in(10) <= VN565_data_out(4);
    CN272_sign_in(10) <= VN565_sign_out(4);
    CN272_data_in(11) <= VN621_data_out(4);
    CN272_sign_in(11) <= VN621_sign_out(4);
    CN272_data_in(12) <= VN715_data_out(4);
    CN272_sign_in(12) <= VN715_sign_out(4);
    CN272_data_in(13) <= VN729_data_out(4);
    CN272_sign_in(13) <= VN729_sign_out(4);
    CN272_data_in(14) <= VN795_data_out(4);
    CN272_sign_in(14) <= VN795_sign_out(4);
    CN272_data_in(15) <= VN863_data_out(4);
    CN272_sign_in(15) <= VN863_sign_out(4);
    CN272_data_in(16) <= VN905_data_out(4);
    CN272_sign_in(16) <= VN905_sign_out(4);
    CN272_data_in(17) <= VN984_data_out(4);
    CN272_sign_in(17) <= VN984_sign_out(4);
    CN272_data_in(18) <= VN1052_data_out(4);
    CN272_sign_in(18) <= VN1052_sign_out(4);
    CN272_data_in(19) <= VN1086_data_out(4);
    CN272_sign_in(19) <= VN1086_sign_out(4);
    CN272_data_in(20) <= VN1127_data_out(4);
    CN272_sign_in(20) <= VN1127_sign_out(4);
    CN272_data_in(21) <= VN1175_data_out(4);
    CN272_sign_in(21) <= VN1175_sign_out(4);
    CN272_data_in(22) <= VN1260_data_out(4);
    CN272_sign_in(22) <= VN1260_sign_out(4);
    CN272_data_in(23) <= VN1313_data_out(4);
    CN272_sign_in(23) <= VN1313_sign_out(4);
    CN272_data_in(24) <= VN1346_data_out(4);
    CN272_sign_in(24) <= VN1346_sign_out(4);
    CN272_data_in(25) <= VN1406_data_out(4);
    CN272_sign_in(25) <= VN1406_sign_out(4);
    CN272_data_in(26) <= VN1433_data_out(4);
    CN272_sign_in(26) <= VN1433_sign_out(4);
    CN272_data_in(27) <= VN1455_data_out(4);
    CN272_sign_in(27) <= VN1455_sign_out(4);
    CN272_data_in(28) <= VN1621_data_out(4);
    CN272_sign_in(28) <= VN1621_sign_out(4);
    CN272_data_in(29) <= VN1657_data_out(4);
    CN272_sign_in(29) <= VN1657_sign_out(4);
    CN272_data_in(30) <= VN1706_data_out(4);
    CN272_sign_in(30) <= VN1706_sign_out(4);
    CN272_data_in(31) <= VN1789_data_out(4);
    CN272_sign_in(31) <= VN1789_sign_out(4);
    CN273_data_in(0) <= VN37_data_out(4);
    CN273_sign_in(0) <= VN37_sign_out(4);
    CN273_data_in(1) <= VN81_data_out(4);
    CN273_sign_in(1) <= VN81_sign_out(4);
    CN273_data_in(2) <= VN156_data_out(4);
    CN273_sign_in(2) <= VN156_sign_out(4);
    CN273_data_in(3) <= VN272_data_out(4);
    CN273_sign_in(3) <= VN272_sign_out(4);
    CN273_data_in(4) <= VN285_data_out(4);
    CN273_sign_in(4) <= VN285_sign_out(4);
    CN273_data_in(5) <= VN371_data_out(4);
    CN273_sign_in(5) <= VN371_sign_out(4);
    CN273_data_in(6) <= VN493_data_out(4);
    CN273_sign_in(6) <= VN493_sign_out(4);
    CN273_data_in(7) <= VN541_data_out(4);
    CN273_sign_in(7) <= VN541_sign_out(4);
    CN273_data_in(8) <= VN659_data_out(4);
    CN273_sign_in(8) <= VN659_sign_out(4);
    CN273_data_in(9) <= VN670_data_out(4);
    CN273_sign_in(9) <= VN670_sign_out(4);
    CN273_data_in(10) <= VN769_data_out(4);
    CN273_sign_in(10) <= VN769_sign_out(4);
    CN273_data_in(11) <= VN826_data_out(4);
    CN273_sign_in(11) <= VN826_sign_out(4);
    CN273_data_in(12) <= VN860_data_out(4);
    CN273_sign_in(12) <= VN860_sign_out(4);
    CN273_data_in(13) <= VN910_data_out(4);
    CN273_sign_in(13) <= VN910_sign_out(4);
    CN273_data_in(14) <= VN963_data_out(4);
    CN273_sign_in(14) <= VN963_sign_out(4);
    CN273_data_in(15) <= VN1007_data_out(4);
    CN273_sign_in(15) <= VN1007_sign_out(4);
    CN273_data_in(16) <= VN1073_data_out(4);
    CN273_sign_in(16) <= VN1073_sign_out(4);
    CN273_data_in(17) <= VN1143_data_out(4);
    CN273_sign_in(17) <= VN1143_sign_out(4);
    CN273_data_in(18) <= VN1198_data_out(4);
    CN273_sign_in(18) <= VN1198_sign_out(4);
    CN273_data_in(19) <= VN1250_data_out(4);
    CN273_sign_in(19) <= VN1250_sign_out(4);
    CN273_data_in(20) <= VN1297_data_out(4);
    CN273_sign_in(20) <= VN1297_sign_out(4);
    CN273_data_in(21) <= VN1358_data_out(4);
    CN273_sign_in(21) <= VN1358_sign_out(4);
    CN273_data_in(22) <= VN1453_data_out(4);
    CN273_sign_in(22) <= VN1453_sign_out(4);
    CN273_data_in(23) <= VN1550_data_out(4);
    CN273_sign_in(23) <= VN1550_sign_out(4);
    CN273_data_in(24) <= VN1726_data_out(4);
    CN273_sign_in(24) <= VN1726_sign_out(4);
    CN273_data_in(25) <= VN1736_data_out(4);
    CN273_sign_in(25) <= VN1736_sign_out(4);
    CN273_data_in(26) <= VN1817_data_out(4);
    CN273_sign_in(26) <= VN1817_sign_out(4);
    CN273_data_in(27) <= VN1910_data_out(4);
    CN273_sign_in(27) <= VN1910_sign_out(4);
    CN273_data_in(28) <= VN1918_data_out(4);
    CN273_sign_in(28) <= VN1918_sign_out(4);
    CN273_data_in(29) <= VN1984_data_out(4);
    CN273_sign_in(29) <= VN1984_sign_out(4);
    CN273_data_in(30) <= VN2031_data_out(4);
    CN273_sign_in(30) <= VN2031_sign_out(4);
    CN273_data_in(31) <= VN2042_data_out(4);
    CN273_sign_in(31) <= VN2042_sign_out(4);
    CN274_data_in(0) <= VN36_data_out(4);
    CN274_sign_in(0) <= VN36_sign_out(4);
    CN274_data_in(1) <= VN164_data_out(4);
    CN274_sign_in(1) <= VN164_sign_out(4);
    CN274_data_in(2) <= VN217_data_out(4);
    CN274_sign_in(2) <= VN217_sign_out(4);
    CN274_data_in(3) <= VN248_data_out(4);
    CN274_sign_in(3) <= VN248_sign_out(4);
    CN274_data_in(4) <= VN390_data_out(4);
    CN274_sign_in(4) <= VN390_sign_out(4);
    CN274_data_in(5) <= VN427_data_out(4);
    CN274_sign_in(5) <= VN427_sign_out(4);
    CN274_data_in(6) <= VN460_data_out(4);
    CN274_sign_in(6) <= VN460_sign_out(4);
    CN274_data_in(7) <= VN551_data_out(4);
    CN274_sign_in(7) <= VN551_sign_out(4);
    CN274_data_in(8) <= VN601_data_out(4);
    CN274_sign_in(8) <= VN601_sign_out(4);
    CN274_data_in(9) <= VN661_data_out(4);
    CN274_sign_in(9) <= VN661_sign_out(4);
    CN274_data_in(10) <= VN739_data_out(4);
    CN274_sign_in(10) <= VN739_sign_out(4);
    CN274_data_in(11) <= VN874_data_out(4);
    CN274_sign_in(11) <= VN874_sign_out(4);
    CN274_data_in(12) <= VN899_data_out(4);
    CN274_sign_in(12) <= VN899_sign_out(4);
    CN274_data_in(13) <= VN944_data_out(4);
    CN274_sign_in(13) <= VN944_sign_out(4);
    CN274_data_in(14) <= VN1033_data_out(4);
    CN274_sign_in(14) <= VN1033_sign_out(4);
    CN274_data_in(15) <= VN1204_data_out(4);
    CN274_sign_in(15) <= VN1204_sign_out(4);
    CN274_data_in(16) <= VN1275_data_out(4);
    CN274_sign_in(16) <= VN1275_sign_out(4);
    CN274_data_in(17) <= VN1282_data_out(4);
    CN274_sign_in(17) <= VN1282_sign_out(4);
    CN274_data_in(18) <= VN1300_data_out(4);
    CN274_sign_in(18) <= VN1300_sign_out(4);
    CN274_data_in(19) <= VN1369_data_out(4);
    CN274_sign_in(19) <= VN1369_sign_out(4);
    CN274_data_in(20) <= VN1398_data_out(4);
    CN274_sign_in(20) <= VN1398_sign_out(4);
    CN274_data_in(21) <= VN1564_data_out(4);
    CN274_sign_in(21) <= VN1564_sign_out(4);
    CN274_data_in(22) <= VN1581_data_out(4);
    CN274_sign_in(22) <= VN1581_sign_out(4);
    CN274_data_in(23) <= VN1641_data_out(4);
    CN274_sign_in(23) <= VN1641_sign_out(4);
    CN274_data_in(24) <= VN1650_data_out(4);
    CN274_sign_in(24) <= VN1650_sign_out(4);
    CN274_data_in(25) <= VN1709_data_out(4);
    CN274_sign_in(25) <= VN1709_sign_out(4);
    CN274_data_in(26) <= VN1985_data_out(4);
    CN274_sign_in(26) <= VN1985_sign_out(4);
    CN274_data_in(27) <= VN2002_data_out(4);
    CN274_sign_in(27) <= VN2002_sign_out(4);
    CN274_data_in(28) <= VN2017_data_out(4);
    CN274_sign_in(28) <= VN2017_sign_out(4);
    CN274_data_in(29) <= VN2019_data_out(4);
    CN274_sign_in(29) <= VN2019_sign_out(4);
    CN274_data_in(30) <= VN2029_data_out(4);
    CN274_sign_in(30) <= VN2029_sign_out(4);
    CN274_data_in(31) <= VN2033_data_out(4);
    CN274_sign_in(31) <= VN2033_sign_out(4);
    CN275_data_in(0) <= VN35_data_out(4);
    CN275_sign_in(0) <= VN35_sign_out(4);
    CN275_data_in(1) <= VN59_data_out(4);
    CN275_sign_in(1) <= VN59_sign_out(4);
    CN275_data_in(2) <= VN128_data_out(4);
    CN275_sign_in(2) <= VN128_sign_out(4);
    CN275_data_in(3) <= VN179_data_out(4);
    CN275_sign_in(3) <= VN179_sign_out(4);
    CN275_data_in(4) <= VN329_data_out(4);
    CN275_sign_in(4) <= VN329_sign_out(4);
    CN275_data_in(5) <= VN394_data_out(4);
    CN275_sign_in(5) <= VN394_sign_out(4);
    CN275_data_in(6) <= VN461_data_out(4);
    CN275_sign_in(6) <= VN461_sign_out(4);
    CN275_data_in(7) <= VN546_data_out(4);
    CN275_sign_in(7) <= VN546_sign_out(4);
    CN275_data_in(8) <= VN597_data_out(4);
    CN275_sign_in(8) <= VN597_sign_out(4);
    CN275_data_in(9) <= VN817_data_out(4);
    CN275_sign_in(9) <= VN817_sign_out(4);
    CN275_data_in(10) <= VN923_data_out(4);
    CN275_sign_in(10) <= VN923_sign_out(4);
    CN275_data_in(11) <= VN958_data_out(4);
    CN275_sign_in(11) <= VN958_sign_out(4);
    CN275_data_in(12) <= VN1022_data_out(4);
    CN275_sign_in(12) <= VN1022_sign_out(4);
    CN275_data_in(13) <= VN1069_data_out(4);
    CN275_sign_in(13) <= VN1069_sign_out(4);
    CN275_data_in(14) <= VN1113_data_out(4);
    CN275_sign_in(14) <= VN1113_sign_out(4);
    CN275_data_in(15) <= VN1115_data_out(4);
    CN275_sign_in(15) <= VN1115_sign_out(4);
    CN275_data_in(16) <= VN1189_data_out(4);
    CN275_sign_in(16) <= VN1189_sign_out(4);
    CN275_data_in(17) <= VN1225_data_out(4);
    CN275_sign_in(17) <= VN1225_sign_out(4);
    CN275_data_in(18) <= VN1286_data_out(4);
    CN275_sign_in(18) <= VN1286_sign_out(4);
    CN275_data_in(19) <= VN1340_data_out(4);
    CN275_sign_in(19) <= VN1340_sign_out(4);
    CN275_data_in(20) <= VN1407_data_out(4);
    CN275_sign_in(20) <= VN1407_sign_out(4);
    CN275_data_in(21) <= VN1440_data_out(4);
    CN275_sign_in(21) <= VN1440_sign_out(4);
    CN275_data_in(22) <= VN1458_data_out(4);
    CN275_sign_in(22) <= VN1458_sign_out(4);
    CN275_data_in(23) <= VN1490_data_out(4);
    CN275_sign_in(23) <= VN1490_sign_out(4);
    CN275_data_in(24) <= VN1668_data_out(4);
    CN275_sign_in(24) <= VN1668_sign_out(4);
    CN275_data_in(25) <= VN1813_data_out(4);
    CN275_sign_in(25) <= VN1813_sign_out(4);
    CN275_data_in(26) <= VN1825_data_out(4);
    CN275_sign_in(26) <= VN1825_sign_out(4);
    CN275_data_in(27) <= VN1848_data_out(4);
    CN275_sign_in(27) <= VN1848_sign_out(4);
    CN275_data_in(28) <= VN1851_data_out(4);
    CN275_sign_in(28) <= VN1851_sign_out(4);
    CN275_data_in(29) <= VN1873_data_out(4);
    CN275_sign_in(29) <= VN1873_sign_out(4);
    CN275_data_in(30) <= VN1875_data_out(4);
    CN275_sign_in(30) <= VN1875_sign_out(4);
    CN275_data_in(31) <= VN1893_data_out(4);
    CN275_sign_in(31) <= VN1893_sign_out(4);
    CN276_data_in(0) <= VN34_data_out(4);
    CN276_sign_in(0) <= VN34_sign_out(4);
    CN276_data_in(1) <= VN69_data_out(4);
    CN276_sign_in(1) <= VN69_sign_out(4);
    CN276_data_in(2) <= VN126_data_out(4);
    CN276_sign_in(2) <= VN126_sign_out(4);
    CN276_data_in(3) <= VN205_data_out(4);
    CN276_sign_in(3) <= VN205_sign_out(4);
    CN276_data_in(4) <= VN259_data_out(4);
    CN276_sign_in(4) <= VN259_sign_out(4);
    CN276_data_in(5) <= VN297_data_out(4);
    CN276_sign_in(5) <= VN297_sign_out(4);
    CN276_data_in(6) <= VN407_data_out(4);
    CN276_sign_in(6) <= VN407_sign_out(4);
    CN276_data_in(7) <= VN492_data_out(4);
    CN276_sign_in(7) <= VN492_sign_out(4);
    CN276_data_in(8) <= VN552_data_out(4);
    CN276_sign_in(8) <= VN552_sign_out(4);
    CN276_data_in(9) <= VN615_data_out(4);
    CN276_sign_in(9) <= VN615_sign_out(4);
    CN276_data_in(10) <= VN667_data_out(4);
    CN276_sign_in(10) <= VN667_sign_out(4);
    CN276_data_in(11) <= VN714_data_out(4);
    CN276_sign_in(11) <= VN714_sign_out(4);
    CN276_data_in(12) <= VN773_data_out(4);
    CN276_sign_in(12) <= VN773_sign_out(4);
    CN276_data_in(13) <= VN801_data_out(4);
    CN276_sign_in(13) <= VN801_sign_out(4);
    CN276_data_in(14) <= VN843_data_out(4);
    CN276_sign_in(14) <= VN843_sign_out(4);
    CN276_data_in(15) <= VN929_data_out(4);
    CN276_sign_in(15) <= VN929_sign_out(4);
    CN276_data_in(16) <= VN969_data_out(4);
    CN276_sign_in(16) <= VN969_sign_out(4);
    CN276_data_in(17) <= VN1009_data_out(4);
    CN276_sign_in(17) <= VN1009_sign_out(4);
    CN276_data_in(18) <= VN1093_data_out(4);
    CN276_sign_in(18) <= VN1093_sign_out(4);
    CN276_data_in(19) <= VN1166_data_out(4);
    CN276_sign_in(19) <= VN1166_sign_out(4);
    CN276_data_in(20) <= VN1191_data_out(4);
    CN276_sign_in(20) <= VN1191_sign_out(4);
    CN276_data_in(21) <= VN1264_data_out(4);
    CN276_sign_in(21) <= VN1264_sign_out(4);
    CN276_data_in(22) <= VN1314_data_out(4);
    CN276_sign_in(22) <= VN1314_sign_out(4);
    CN276_data_in(23) <= VN1456_data_out(4);
    CN276_sign_in(23) <= VN1456_sign_out(4);
    CN276_data_in(24) <= VN1496_data_out(4);
    CN276_sign_in(24) <= VN1496_sign_out(4);
    CN276_data_in(25) <= VN1533_data_out(4);
    CN276_sign_in(25) <= VN1533_sign_out(4);
    CN276_data_in(26) <= VN1543_data_out(4);
    CN276_sign_in(26) <= VN1543_sign_out(4);
    CN276_data_in(27) <= VN1578_data_out(4);
    CN276_sign_in(27) <= VN1578_sign_out(4);
    CN276_data_in(28) <= VN1644_data_out(4);
    CN276_sign_in(28) <= VN1644_sign_out(4);
    CN276_data_in(29) <= VN1653_data_out(4);
    CN276_sign_in(29) <= VN1653_sign_out(4);
    CN276_data_in(30) <= VN1688_data_out(4);
    CN276_sign_in(30) <= VN1688_sign_out(4);
    CN276_data_in(31) <= VN1790_data_out(4);
    CN276_sign_in(31) <= VN1790_sign_out(4);
    CN277_data_in(0) <= VN33_data_out(4);
    CN277_sign_in(0) <= VN33_sign_out(4);
    CN277_data_in(1) <= VN64_data_out(4);
    CN277_sign_in(1) <= VN64_sign_out(4);
    CN277_data_in(2) <= VN162_data_out(4);
    CN277_sign_in(2) <= VN162_sign_out(4);
    CN277_data_in(3) <= VN185_data_out(4);
    CN277_sign_in(3) <= VN185_sign_out(4);
    CN277_data_in(4) <= VN252_data_out(4);
    CN277_sign_in(4) <= VN252_sign_out(4);
    CN277_data_in(5) <= VN295_data_out(4);
    CN277_sign_in(5) <= VN295_sign_out(4);
    CN277_data_in(6) <= VN334_data_out(4);
    CN277_sign_in(6) <= VN334_sign_out(4);
    CN277_data_in(7) <= VN391_data_out(4);
    CN277_sign_in(7) <= VN391_sign_out(4);
    CN277_data_in(8) <= VN404_data_out(4);
    CN277_sign_in(8) <= VN404_sign_out(4);
    CN277_data_in(9) <= VN484_data_out(4);
    CN277_sign_in(9) <= VN484_sign_out(4);
    CN277_data_in(10) <= VN540_data_out(4);
    CN277_sign_in(10) <= VN540_sign_out(4);
    CN277_data_in(11) <= VN582_data_out(4);
    CN277_sign_in(11) <= VN582_sign_out(4);
    CN277_data_in(12) <= VN682_data_out(4);
    CN277_sign_in(12) <= VN682_sign_out(4);
    CN277_data_in(13) <= VN736_data_out(4);
    CN277_sign_in(13) <= VN736_sign_out(4);
    CN277_data_in(14) <= VN854_data_out(4);
    CN277_sign_in(14) <= VN854_sign_out(4);
    CN277_data_in(15) <= VN914_data_out(4);
    CN277_sign_in(15) <= VN914_sign_out(4);
    CN277_data_in(16) <= VN998_data_out(4);
    CN277_sign_in(16) <= VN998_sign_out(4);
    CN277_data_in(17) <= VN1116_data_out(4);
    CN277_sign_in(17) <= VN1116_sign_out(4);
    CN277_data_in(18) <= VN1266_data_out(4);
    CN277_sign_in(18) <= VN1266_sign_out(4);
    CN277_data_in(19) <= VN1371_data_out(4);
    CN277_sign_in(19) <= VN1371_sign_out(4);
    CN277_data_in(20) <= VN1394_data_out(4);
    CN277_sign_in(20) <= VN1394_sign_out(4);
    CN277_data_in(21) <= VN1565_data_out(4);
    CN277_sign_in(21) <= VN1565_sign_out(4);
    CN277_data_in(22) <= VN1599_data_out(4);
    CN277_sign_in(22) <= VN1599_sign_out(4);
    CN277_data_in(23) <= VN1669_data_out(4);
    CN277_sign_in(23) <= VN1669_sign_out(4);
    CN277_data_in(24) <= VN1751_data_out(4);
    CN277_sign_in(24) <= VN1751_sign_out(4);
    CN277_data_in(25) <= VN1758_data_out(4);
    CN277_sign_in(25) <= VN1758_sign_out(4);
    CN277_data_in(26) <= VN1808_data_out(4);
    CN277_sign_in(26) <= VN1808_sign_out(4);
    CN277_data_in(27) <= VN1936_data_out(4);
    CN277_sign_in(27) <= VN1936_sign_out(4);
    CN277_data_in(28) <= VN1951_data_out(4);
    CN277_sign_in(28) <= VN1951_sign_out(4);
    CN277_data_in(29) <= VN2000_data_out(4);
    CN277_sign_in(29) <= VN2000_sign_out(4);
    CN277_data_in(30) <= VN2004_data_out(4);
    CN277_sign_in(30) <= VN2004_sign_out(4);
    CN277_data_in(31) <= VN2010_data_out(4);
    CN277_sign_in(31) <= VN2010_sign_out(4);
    CN278_data_in(0) <= VN32_data_out(4);
    CN278_sign_in(0) <= VN32_sign_out(4);
    CN278_data_in(1) <= VN70_data_out(4);
    CN278_sign_in(1) <= VN70_sign_out(4);
    CN278_data_in(2) <= VN141_data_out(4);
    CN278_sign_in(2) <= VN141_sign_out(4);
    CN278_data_in(3) <= VN229_data_out(4);
    CN278_sign_in(3) <= VN229_sign_out(4);
    CN278_data_in(4) <= VN328_data_out(4);
    CN278_sign_in(4) <= VN328_sign_out(4);
    CN278_data_in(5) <= VN388_data_out(4);
    CN278_sign_in(5) <= VN388_sign_out(4);
    CN278_data_in(6) <= VN423_data_out(4);
    CN278_sign_in(6) <= VN423_sign_out(4);
    CN278_data_in(7) <= VN502_data_out(4);
    CN278_sign_in(7) <= VN502_sign_out(4);
    CN278_data_in(8) <= VN509_data_out(4);
    CN278_sign_in(8) <= VN509_sign_out(4);
    CN278_data_in(9) <= VN630_data_out(4);
    CN278_sign_in(9) <= VN630_sign_out(4);
    CN278_data_in(10) <= VN689_data_out(4);
    CN278_sign_in(10) <= VN689_sign_out(4);
    CN278_data_in(11) <= VN766_data_out(4);
    CN278_sign_in(11) <= VN766_sign_out(4);
    CN278_data_in(12) <= VN819_data_out(4);
    CN278_sign_in(12) <= VN819_sign_out(4);
    CN278_data_in(13) <= VN847_data_out(4);
    CN278_sign_in(13) <= VN847_sign_out(4);
    CN278_data_in(14) <= VN915_data_out(4);
    CN278_sign_in(14) <= VN915_sign_out(4);
    CN278_data_in(15) <= VN986_data_out(4);
    CN278_sign_in(15) <= VN986_sign_out(4);
    CN278_data_in(16) <= VN1044_data_out(4);
    CN278_sign_in(16) <= VN1044_sign_out(4);
    CN278_data_in(17) <= VN1102_data_out(4);
    CN278_sign_in(17) <= VN1102_sign_out(4);
    CN278_data_in(18) <= VN1163_data_out(4);
    CN278_sign_in(18) <= VN1163_sign_out(4);
    CN278_data_in(19) <= VN1196_data_out(4);
    CN278_sign_in(19) <= VN1196_sign_out(4);
    CN278_data_in(20) <= VN1236_data_out(4);
    CN278_sign_in(20) <= VN1236_sign_out(4);
    CN278_data_in(21) <= VN1306_data_out(4);
    CN278_sign_in(21) <= VN1306_sign_out(4);
    CN278_data_in(22) <= VN1329_data_out(4);
    CN278_sign_in(22) <= VN1329_sign_out(4);
    CN278_data_in(23) <= VN1422_data_out(4);
    CN278_sign_in(23) <= VN1422_sign_out(4);
    CN278_data_in(24) <= VN1434_data_out(4);
    CN278_sign_in(24) <= VN1434_sign_out(4);
    CN278_data_in(25) <= VN1588_data_out(4);
    CN278_sign_in(25) <= VN1588_sign_out(4);
    CN278_data_in(26) <= VN1638_data_out(4);
    CN278_sign_in(26) <= VN1638_sign_out(4);
    CN278_data_in(27) <= VN1679_data_out(4);
    CN278_sign_in(27) <= VN1679_sign_out(4);
    CN278_data_in(28) <= VN1782_data_out(4);
    CN278_sign_in(28) <= VN1782_sign_out(4);
    CN278_data_in(29) <= VN1854_data_out(4);
    CN278_sign_in(29) <= VN1854_sign_out(4);
    CN278_data_in(30) <= VN1934_data_out(4);
    CN278_sign_in(30) <= VN1934_sign_out(4);
    CN278_data_in(31) <= VN1949_data_out(4);
    CN278_sign_in(31) <= VN1949_sign_out(4);
    CN279_data_in(0) <= VN31_data_out(4);
    CN279_sign_in(0) <= VN31_sign_out(4);
    CN279_data_in(1) <= VN58_data_out(4);
    CN279_sign_in(1) <= VN58_sign_out(4);
    CN279_data_in(2) <= VN144_data_out(4);
    CN279_sign_in(2) <= VN144_sign_out(4);
    CN279_data_in(3) <= VN219_data_out(4);
    CN279_sign_in(3) <= VN219_sign_out(4);
    CN279_data_in(4) <= VN239_data_out(4);
    CN279_sign_in(4) <= VN239_sign_out(4);
    CN279_data_in(5) <= VN368_data_out(4);
    CN279_sign_in(5) <= VN368_sign_out(4);
    CN279_data_in(6) <= VN444_data_out(4);
    CN279_sign_in(6) <= VN444_sign_out(4);
    CN279_data_in(7) <= VN450_data_out(4);
    CN279_sign_in(7) <= VN450_sign_out(4);
    CN279_data_in(8) <= VN614_data_out(4);
    CN279_sign_in(8) <= VN614_sign_out(4);
    CN279_data_in(9) <= VN660_data_out(4);
    CN279_sign_in(9) <= VN660_sign_out(4);
    CN279_data_in(10) <= VN851_data_out(4);
    CN279_sign_in(10) <= VN851_sign_out(4);
    CN279_data_in(11) <= VN939_data_out(4);
    CN279_sign_in(11) <= VN939_sign_out(4);
    CN279_data_in(12) <= VN972_data_out(4);
    CN279_sign_in(12) <= VN972_sign_out(4);
    CN279_data_in(13) <= VN1054_data_out(4);
    CN279_sign_in(13) <= VN1054_sign_out(4);
    CN279_data_in(14) <= VN1208_data_out(4);
    CN279_sign_in(14) <= VN1208_sign_out(4);
    CN279_data_in(15) <= VN1273_data_out(4);
    CN279_sign_in(15) <= VN1273_sign_out(4);
    CN279_data_in(16) <= VN1294_data_out(4);
    CN279_sign_in(16) <= VN1294_sign_out(4);
    CN279_data_in(17) <= VN1352_data_out(4);
    CN279_sign_in(17) <= VN1352_sign_out(4);
    CN279_data_in(18) <= VN1401_data_out(4);
    CN279_sign_in(18) <= VN1401_sign_out(4);
    CN279_data_in(19) <= VN1452_data_out(4);
    CN279_sign_in(19) <= VN1452_sign_out(4);
    CN279_data_in(20) <= VN1460_data_out(4);
    CN279_sign_in(20) <= VN1460_sign_out(4);
    CN279_data_in(21) <= VN1471_data_out(4);
    CN279_sign_in(21) <= VN1471_sign_out(4);
    CN279_data_in(22) <= VN1622_data_out(4);
    CN279_sign_in(22) <= VN1622_sign_out(4);
    CN279_data_in(23) <= VN1676_data_out(4);
    CN279_sign_in(23) <= VN1676_sign_out(4);
    CN279_data_in(24) <= VN1768_data_out(4);
    CN279_sign_in(24) <= VN1768_sign_out(4);
    CN279_data_in(25) <= VN1779_data_out(4);
    CN279_sign_in(25) <= VN1779_sign_out(4);
    CN279_data_in(26) <= VN1964_data_out(4);
    CN279_sign_in(26) <= VN1964_sign_out(4);
    CN279_data_in(27) <= VN1991_data_out(4);
    CN279_sign_in(27) <= VN1991_sign_out(4);
    CN279_data_in(28) <= VN2007_data_out(4);
    CN279_sign_in(28) <= VN2007_sign_out(4);
    CN279_data_in(29) <= VN2011_data_out(4);
    CN279_sign_in(29) <= VN2011_sign_out(4);
    CN279_data_in(30) <= VN2013_data_out(4);
    CN279_sign_in(30) <= VN2013_sign_out(4);
    CN279_data_in(31) <= VN2025_data_out(4);
    CN279_sign_in(31) <= VN2025_sign_out(4);
    CN280_data_in(0) <= VN30_data_out(4);
    CN280_sign_in(0) <= VN30_sign_out(4);
    CN280_data_in(1) <= VN84_data_out(4);
    CN280_sign_in(1) <= VN84_sign_out(4);
    CN280_data_in(2) <= VN129_data_out(4);
    CN280_sign_in(2) <= VN129_sign_out(4);
    CN280_data_in(3) <= VN215_data_out(4);
    CN280_sign_in(3) <= VN215_sign_out(4);
    CN280_data_in(4) <= VN233_data_out(4);
    CN280_sign_in(4) <= VN233_sign_out(4);
    CN280_data_in(5) <= VN310_data_out(4);
    CN280_sign_in(5) <= VN310_sign_out(4);
    CN280_data_in(6) <= VN376_data_out(4);
    CN280_sign_in(6) <= VN376_sign_out(4);
    CN280_data_in(7) <= VN445_data_out(4);
    CN280_sign_in(7) <= VN445_sign_out(4);
    CN280_data_in(8) <= VN505_data_out(4);
    CN280_sign_in(8) <= VN505_sign_out(4);
    CN280_data_in(9) <= VN555_data_out(4);
    CN280_sign_in(9) <= VN555_sign_out(4);
    CN280_data_in(10) <= VN606_data_out(4);
    CN280_sign_in(10) <= VN606_sign_out(4);
    CN280_data_in(11) <= VN675_data_out(4);
    CN280_sign_in(11) <= VN675_sign_out(4);
    CN280_data_in(12) <= VN723_data_out(4);
    CN280_sign_in(12) <= VN723_sign_out(4);
    CN280_data_in(13) <= VN824_data_out(4);
    CN280_sign_in(13) <= VN824_sign_out(4);
    CN280_data_in(14) <= VN840_data_out(4);
    CN280_sign_in(14) <= VN840_sign_out(4);
    CN280_data_in(15) <= VN989_data_out(4);
    CN280_sign_in(15) <= VN989_sign_out(4);
    CN280_data_in(16) <= VN1049_data_out(4);
    CN280_sign_in(16) <= VN1049_sign_out(4);
    CN280_data_in(17) <= VN1084_data_out(4);
    CN280_sign_in(17) <= VN1084_sign_out(4);
    CN280_data_in(18) <= VN1136_data_out(4);
    CN280_sign_in(18) <= VN1136_sign_out(4);
    CN280_data_in(19) <= VN1223_data_out(4);
    CN280_sign_in(19) <= VN1223_sign_out(4);
    CN280_data_in(20) <= VN1229_data_out(4);
    CN280_sign_in(20) <= VN1229_sign_out(4);
    CN280_data_in(21) <= VN1316_data_out(4);
    CN280_sign_in(21) <= VN1316_sign_out(4);
    CN280_data_in(22) <= VN1360_data_out(4);
    CN280_sign_in(22) <= VN1360_sign_out(4);
    CN280_data_in(23) <= VN1386_data_out(4);
    CN280_sign_in(23) <= VN1386_sign_out(4);
    CN280_data_in(24) <= VN1424_data_out(4);
    CN280_sign_in(24) <= VN1424_sign_out(4);
    CN280_data_in(25) <= VN1600_data_out(4);
    CN280_sign_in(25) <= VN1600_sign_out(4);
    CN280_data_in(26) <= VN1708_data_out(4);
    CN280_sign_in(26) <= VN1708_sign_out(4);
    CN280_data_in(27) <= VN1740_data_out(4);
    CN280_sign_in(27) <= VN1740_sign_out(4);
    CN280_data_in(28) <= VN1777_data_out(4);
    CN280_sign_in(28) <= VN1777_sign_out(4);
    CN280_data_in(29) <= VN1896_data_out(4);
    CN280_sign_in(29) <= VN1896_sign_out(4);
    CN280_data_in(30) <= VN1924_data_out(4);
    CN280_sign_in(30) <= VN1924_sign_out(4);
    CN280_data_in(31) <= VN1927_data_out(4);
    CN280_sign_in(31) <= VN1927_sign_out(4);
    CN281_data_in(0) <= VN29_data_out(4);
    CN281_sign_in(0) <= VN29_sign_out(4);
    CN281_data_in(1) <= VN90_data_out(4);
    CN281_sign_in(1) <= VN90_sign_out(4);
    CN281_data_in(2) <= VN163_data_out(4);
    CN281_sign_in(2) <= VN163_sign_out(4);
    CN281_data_in(3) <= VN182_data_out(4);
    CN281_sign_in(3) <= VN182_sign_out(4);
    CN281_data_in(4) <= VN236_data_out(4);
    CN281_sign_in(4) <= VN236_sign_out(4);
    CN281_data_in(5) <= VN298_data_out(4);
    CN281_sign_in(5) <= VN298_sign_out(4);
    CN281_data_in(6) <= VN340_data_out(4);
    CN281_sign_in(6) <= VN340_sign_out(4);
    CN281_data_in(7) <= VN422_data_out(4);
    CN281_sign_in(7) <= VN422_sign_out(4);
    CN281_data_in(8) <= VN449_data_out(4);
    CN281_sign_in(8) <= VN449_sign_out(4);
    CN281_data_in(9) <= VN557_data_out(4);
    CN281_sign_in(9) <= VN557_sign_out(4);
    CN281_data_in(10) <= VN569_data_out(4);
    CN281_sign_in(10) <= VN569_sign_out(4);
    CN281_data_in(11) <= VN648_data_out(4);
    CN281_sign_in(11) <= VN648_sign_out(4);
    CN281_data_in(12) <= VN700_data_out(4);
    CN281_sign_in(12) <= VN700_sign_out(4);
    CN281_data_in(13) <= VN771_data_out(4);
    CN281_sign_in(13) <= VN771_sign_out(4);
    CN281_data_in(14) <= VN799_data_out(4);
    CN281_sign_in(14) <= VN799_sign_out(4);
    CN281_data_in(15) <= VN875_data_out(4);
    CN281_sign_in(15) <= VN875_sign_out(4);
    CN281_data_in(16) <= VN931_data_out(4);
    CN281_sign_in(16) <= VN931_sign_out(4);
    CN281_data_in(17) <= VN950_data_out(4);
    CN281_sign_in(17) <= VN950_sign_out(4);
    CN281_data_in(18) <= VN1055_data_out(4);
    CN281_sign_in(18) <= VN1055_sign_out(4);
    CN281_data_in(19) <= VN1060_data_out(4);
    CN281_sign_in(19) <= VN1060_sign_out(4);
    CN281_data_in(20) <= VN1099_data_out(4);
    CN281_sign_in(20) <= VN1099_sign_out(4);
    CN281_data_in(21) <= VN1120_data_out(4);
    CN281_sign_in(21) <= VN1120_sign_out(4);
    CN281_data_in(22) <= VN1190_data_out(4);
    CN281_sign_in(22) <= VN1190_sign_out(4);
    CN281_data_in(23) <= VN1237_data_out(4);
    CN281_sign_in(23) <= VN1237_sign_out(4);
    CN281_data_in(24) <= VN1308_data_out(4);
    CN281_sign_in(24) <= VN1308_sign_out(4);
    CN281_data_in(25) <= VN1356_data_out(4);
    CN281_sign_in(25) <= VN1356_sign_out(4);
    CN281_data_in(26) <= VN1545_data_out(4);
    CN281_sign_in(26) <= VN1545_sign_out(4);
    CN281_data_in(27) <= VN1560_data_out(4);
    CN281_sign_in(27) <= VN1560_sign_out(4);
    CN281_data_in(28) <= VN1591_data_out(4);
    CN281_sign_in(28) <= VN1591_sign_out(4);
    CN281_data_in(29) <= VN1617_data_out(4);
    CN281_sign_in(29) <= VN1617_sign_out(4);
    CN281_data_in(30) <= VN1666_data_out(4);
    CN281_sign_in(30) <= VN1666_sign_out(4);
    CN281_data_in(31) <= VN1791_data_out(4);
    CN281_sign_in(31) <= VN1791_sign_out(4);
    CN282_data_in(0) <= VN28_data_out(4);
    CN282_sign_in(0) <= VN28_sign_out(4);
    CN282_data_in(1) <= VN74_data_out(4);
    CN282_sign_in(1) <= VN74_sign_out(4);
    CN282_data_in(2) <= VN125_data_out(4);
    CN282_sign_in(2) <= VN125_sign_out(4);
    CN282_data_in(3) <= VN200_data_out(4);
    CN282_sign_in(3) <= VN200_sign_out(4);
    CN282_data_in(4) <= VN226_data_out(4);
    CN282_sign_in(4) <= VN226_sign_out(4);
    CN282_data_in(5) <= VN338_data_out(4);
    CN282_sign_in(5) <= VN338_sign_out(4);
    CN282_data_in(6) <= VN413_data_out(4);
    CN282_sign_in(6) <= VN413_sign_out(4);
    CN282_data_in(7) <= VN500_data_out(4);
    CN282_sign_in(7) <= VN500_sign_out(4);
    CN282_data_in(8) <= VN573_data_out(4);
    CN282_sign_in(8) <= VN573_sign_out(4);
    CN282_data_in(9) <= VN626_data_out(4);
    CN282_sign_in(9) <= VN626_sign_out(4);
    CN282_data_in(10) <= VN746_data_out(4);
    CN282_sign_in(10) <= VN746_sign_out(4);
    CN282_data_in(11) <= VN859_data_out(4);
    CN282_sign_in(11) <= VN859_sign_out(4);
    CN282_data_in(12) <= VN940_data_out(4);
    CN282_sign_in(12) <= VN940_sign_out(4);
    CN282_data_in(13) <= VN960_data_out(4);
    CN282_sign_in(13) <= VN960_sign_out(4);
    CN282_data_in(14) <= VN1043_data_out(4);
    CN282_sign_in(14) <= VN1043_sign_out(4);
    CN282_data_in(15) <= VN1203_data_out(4);
    CN282_sign_in(15) <= VN1203_sign_out(4);
    CN282_data_in(16) <= VN1265_data_out(4);
    CN282_sign_in(16) <= VN1265_sign_out(4);
    CN282_data_in(17) <= VN1298_data_out(4);
    CN282_sign_in(17) <= VN1298_sign_out(4);
    CN282_data_in(18) <= VN1331_data_out(4);
    CN282_sign_in(18) <= VN1331_sign_out(4);
    CN282_data_in(19) <= VN1361_data_out(4);
    CN282_sign_in(19) <= VN1361_sign_out(4);
    CN282_data_in(20) <= VN1388_data_out(4);
    CN282_sign_in(20) <= VN1388_sign_out(4);
    CN282_data_in(21) <= VN1541_data_out(4);
    CN282_sign_in(21) <= VN1541_sign_out(4);
    CN282_data_in(22) <= VN1605_data_out(4);
    CN282_sign_in(22) <= VN1605_sign_out(4);
    CN282_data_in(23) <= VN1627_data_out(4);
    CN282_sign_in(23) <= VN1627_sign_out(4);
    CN282_data_in(24) <= VN1766_data_out(4);
    CN282_sign_in(24) <= VN1766_sign_out(4);
    CN282_data_in(25) <= VN1785_data_out(4);
    CN282_sign_in(25) <= VN1785_sign_out(4);
    CN282_data_in(26) <= VN1974_data_out(4);
    CN282_sign_in(26) <= VN1974_sign_out(4);
    CN282_data_in(27) <= VN2003_data_out(4);
    CN282_sign_in(27) <= VN2003_sign_out(4);
    CN282_data_in(28) <= VN2009_data_out(4);
    CN282_sign_in(28) <= VN2009_sign_out(4);
    CN282_data_in(29) <= VN2040_data_out(4);
    CN282_sign_in(29) <= VN2040_sign_out(4);
    CN282_data_in(30) <= VN2041_data_out(4);
    CN282_sign_in(30) <= VN2041_sign_out(4);
    CN282_data_in(31) <= VN2047_data_out(4);
    CN282_sign_in(31) <= VN2047_sign_out(4);
    CN283_data_in(0) <= VN27_data_out(4);
    CN283_sign_in(0) <= VN27_sign_out(4);
    CN283_data_in(1) <= VN76_data_out(4);
    CN283_sign_in(1) <= VN76_sign_out(4);
    CN283_data_in(2) <= VN153_data_out(4);
    CN283_sign_in(2) <= VN153_sign_out(4);
    CN283_data_in(3) <= VN201_data_out(4);
    CN283_sign_in(3) <= VN201_sign_out(4);
    CN283_data_in(4) <= VN260_data_out(4);
    CN283_sign_in(4) <= VN260_sign_out(4);
    CN283_data_in(5) <= VN294_data_out(4);
    CN283_sign_in(5) <= VN294_sign_out(4);
    CN283_data_in(6) <= VN374_data_out(4);
    CN283_sign_in(6) <= VN374_sign_out(4);
    CN283_data_in(7) <= VN431_data_out(4);
    CN283_sign_in(7) <= VN431_sign_out(4);
    CN283_data_in(8) <= VN482_data_out(4);
    CN283_sign_in(8) <= VN482_sign_out(4);
    CN283_data_in(9) <= VN616_data_out(4);
    CN283_sign_in(9) <= VN616_sign_out(4);
    CN283_data_in(10) <= VN650_data_out(4);
    CN283_sign_in(10) <= VN650_sign_out(4);
    CN283_data_in(11) <= VN692_data_out(4);
    CN283_sign_in(11) <= VN692_sign_out(4);
    CN283_data_in(12) <= VN756_data_out(4);
    CN283_sign_in(12) <= VN756_sign_out(4);
    CN283_data_in(13) <= VN810_data_out(4);
    CN283_sign_in(13) <= VN810_sign_out(4);
    CN283_data_in(14) <= VN870_data_out(4);
    CN283_sign_in(14) <= VN870_sign_out(4);
    CN283_data_in(15) <= VN955_data_out(4);
    CN283_sign_in(15) <= VN955_sign_out(4);
    CN283_data_in(16) <= VN1012_data_out(4);
    CN283_sign_in(16) <= VN1012_sign_out(4);
    CN283_data_in(17) <= VN1075_data_out(4);
    CN283_sign_in(17) <= VN1075_sign_out(4);
    CN283_data_in(18) <= VN1147_data_out(4);
    CN283_sign_in(18) <= VN1147_sign_out(4);
    CN283_data_in(19) <= VN1276_data_out(4);
    CN283_sign_in(19) <= VN1276_sign_out(4);
    CN283_data_in(20) <= VN1351_data_out(4);
    CN283_sign_in(20) <= VN1351_sign_out(4);
    CN283_data_in(21) <= VN1396_data_out(4);
    CN283_sign_in(21) <= VN1396_sign_out(4);
    CN283_data_in(22) <= VN1435_data_out(4);
    CN283_sign_in(22) <= VN1435_sign_out(4);
    CN283_data_in(23) <= VN1491_data_out(4);
    CN283_sign_in(23) <= VN1491_sign_out(4);
    CN283_data_in(24) <= VN1524_data_out(4);
    CN283_sign_in(24) <= VN1524_sign_out(4);
    CN283_data_in(25) <= VN1585_data_out(4);
    CN283_sign_in(25) <= VN1585_sign_out(4);
    CN283_data_in(26) <= VN1697_data_out(4);
    CN283_sign_in(26) <= VN1697_sign_out(4);
    CN283_data_in(27) <= VN1829_data_out(4);
    CN283_sign_in(27) <= VN1829_sign_out(4);
    CN283_data_in(28) <= VN1835_data_out(4);
    CN283_sign_in(28) <= VN1835_sign_out(4);
    CN283_data_in(29) <= VN1900_data_out(4);
    CN283_sign_in(29) <= VN1900_sign_out(4);
    CN283_data_in(30) <= VN1947_data_out(4);
    CN283_sign_in(30) <= VN1947_sign_out(4);
    CN283_data_in(31) <= VN1955_data_out(4);
    CN283_sign_in(31) <= VN1955_sign_out(4);
    CN284_data_in(0) <= VN26_data_out(4);
    CN284_sign_in(0) <= VN26_sign_out(4);
    CN284_data_in(1) <= VN100_data_out(4);
    CN284_sign_in(1) <= VN100_sign_out(4);
    CN284_data_in(2) <= VN137_data_out(4);
    CN284_sign_in(2) <= VN137_sign_out(4);
    CN284_data_in(3) <= VN181_data_out(4);
    CN284_sign_in(3) <= VN181_sign_out(4);
    CN284_data_in(4) <= VN245_data_out(4);
    CN284_sign_in(4) <= VN245_sign_out(4);
    CN284_data_in(5) <= VN320_data_out(4);
    CN284_sign_in(5) <= VN320_sign_out(4);
    CN284_data_in(6) <= VN353_data_out(4);
    CN284_sign_in(6) <= VN353_sign_out(4);
    CN284_data_in(7) <= VN436_data_out(4);
    CN284_sign_in(7) <= VN436_sign_out(4);
    CN284_data_in(8) <= VN488_data_out(4);
    CN284_sign_in(8) <= VN488_sign_out(4);
    CN284_data_in(9) <= VN517_data_out(4);
    CN284_sign_in(9) <= VN517_sign_out(4);
    CN284_data_in(10) <= VN572_data_out(4);
    CN284_sign_in(10) <= VN572_sign_out(4);
    CN284_data_in(11) <= VN662_data_out(4);
    CN284_sign_in(11) <= VN662_sign_out(4);
    CN284_data_in(12) <= VN701_data_out(4);
    CN284_sign_in(12) <= VN701_sign_out(4);
    CN284_data_in(13) <= VN749_data_out(4);
    CN284_sign_in(13) <= VN749_sign_out(4);
    CN284_data_in(14) <= VN803_data_out(4);
    CN284_sign_in(14) <= VN803_sign_out(4);
    CN284_data_in(15) <= VN881_data_out(4);
    CN284_sign_in(15) <= VN881_sign_out(4);
    CN284_data_in(16) <= VN928_data_out(4);
    CN284_sign_in(16) <= VN928_sign_out(4);
    CN284_data_in(17) <= VN961_data_out(4);
    CN284_sign_in(17) <= VN961_sign_out(4);
    CN284_data_in(18) <= VN1018_data_out(4);
    CN284_sign_in(18) <= VN1018_sign_out(4);
    CN284_data_in(19) <= VN1088_data_out(4);
    CN284_sign_in(19) <= VN1088_sign_out(4);
    CN284_data_in(20) <= VN1128_data_out(4);
    CN284_sign_in(20) <= VN1128_sign_out(4);
    CN284_data_in(21) <= VN1164_data_out(4);
    CN284_sign_in(21) <= VN1164_sign_out(4);
    CN284_data_in(22) <= VN1211_data_out(4);
    CN284_sign_in(22) <= VN1211_sign_out(4);
    CN284_data_in(23) <= VN1252_data_out(4);
    CN284_sign_in(23) <= VN1252_sign_out(4);
    CN284_data_in(24) <= VN1291_data_out(4);
    CN284_sign_in(24) <= VN1291_sign_out(4);
    CN284_data_in(25) <= VN1374_data_out(4);
    CN284_sign_in(25) <= VN1374_sign_out(4);
    CN284_data_in(26) <= VN1418_data_out(4);
    CN284_sign_in(26) <= VN1418_sign_out(4);
    CN284_data_in(27) <= VN1432_data_out(4);
    CN284_sign_in(27) <= VN1432_sign_out(4);
    CN284_data_in(28) <= VN1583_data_out(4);
    CN284_sign_in(28) <= VN1583_sign_out(4);
    CN284_data_in(29) <= VN1640_data_out(4);
    CN284_sign_in(29) <= VN1640_sign_out(4);
    CN284_data_in(30) <= VN1684_data_out(4);
    CN284_sign_in(30) <= VN1684_sign_out(4);
    CN284_data_in(31) <= VN1792_data_out(4);
    CN284_sign_in(31) <= VN1792_sign_out(4);
    CN285_data_in(0) <= VN25_data_out(4);
    CN285_sign_in(0) <= VN25_sign_out(4);
    CN285_data_in(1) <= VN82_data_out(4);
    CN285_sign_in(1) <= VN82_sign_out(4);
    CN285_data_in(2) <= VN165_data_out(4);
    CN285_sign_in(2) <= VN165_sign_out(4);
    CN285_data_in(3) <= VN172_data_out(4);
    CN285_sign_in(3) <= VN172_sign_out(4);
    CN285_data_in(4) <= VN255_data_out(4);
    CN285_sign_in(4) <= VN255_sign_out(4);
    CN285_data_in(5) <= VN304_data_out(4);
    CN285_sign_in(5) <= VN304_sign_out(4);
    CN285_data_in(6) <= VN355_data_out(4);
    CN285_sign_in(6) <= VN355_sign_out(4);
    CN285_data_in(7) <= VN447_data_out(4);
    CN285_sign_in(7) <= VN447_sign_out(4);
    CN285_data_in(8) <= VN456_data_out(4);
    CN285_sign_in(8) <= VN456_sign_out(4);
    CN285_data_in(9) <= VN524_data_out(4);
    CN285_sign_in(9) <= VN524_sign_out(4);
    CN285_data_in(10) <= VN567_data_out(4);
    CN285_sign_in(10) <= VN567_sign_out(4);
    CN285_data_in(11) <= VN658_data_out(4);
    CN285_sign_in(11) <= VN658_sign_out(4);
    CN285_data_in(12) <= VN674_data_out(4);
    CN285_sign_in(12) <= VN674_sign_out(4);
    CN285_data_in(13) <= VN753_data_out(4);
    CN285_sign_in(13) <= VN753_sign_out(4);
    CN285_data_in(14) <= VN780_data_out(4);
    CN285_sign_in(14) <= VN780_sign_out(4);
    CN285_data_in(15) <= VN901_data_out(4);
    CN285_sign_in(15) <= VN901_sign_out(4);
    CN285_data_in(16) <= VN949_data_out(4);
    CN285_sign_in(16) <= VN949_sign_out(4);
    CN285_data_in(17) <= VN1081_data_out(4);
    CN285_sign_in(17) <= VN1081_sign_out(4);
    CN285_data_in(18) <= VN1139_data_out(4);
    CN285_sign_in(18) <= VN1139_sign_out(4);
    CN285_data_in(19) <= VN1178_data_out(4);
    CN285_sign_in(19) <= VN1178_sign_out(4);
    CN285_data_in(20) <= VN1232_data_out(4);
    CN285_sign_in(20) <= VN1232_sign_out(4);
    CN285_data_in(21) <= VN1281_data_out(4);
    CN285_sign_in(21) <= VN1281_sign_out(4);
    CN285_data_in(22) <= VN1288_data_out(4);
    CN285_sign_in(22) <= VN1288_sign_out(4);
    CN285_data_in(23) <= VN1380_data_out(4);
    CN285_sign_in(23) <= VN1380_sign_out(4);
    CN285_data_in(24) <= VN1419_data_out(4);
    CN285_sign_in(24) <= VN1419_sign_out(4);
    CN285_data_in(25) <= VN1474_data_out(4);
    CN285_sign_in(25) <= VN1474_sign_out(4);
    CN285_data_in(26) <= VN1504_data_out(4);
    CN285_sign_in(26) <= VN1504_sign_out(4);
    CN285_data_in(27) <= VN1593_data_out(4);
    CN285_sign_in(27) <= VN1593_sign_out(4);
    CN285_data_in(28) <= VN1701_data_out(4);
    CN285_sign_in(28) <= VN1701_sign_out(4);
    CN285_data_in(29) <= VN1731_data_out(4);
    CN285_sign_in(29) <= VN1731_sign_out(4);
    CN285_data_in(30) <= VN1755_data_out(4);
    CN285_sign_in(30) <= VN1755_sign_out(4);
    CN285_data_in(31) <= VN1865_data_out(4);
    CN285_sign_in(31) <= VN1865_sign_out(4);
    CN286_data_in(0) <= VN24_data_out(4);
    CN286_sign_in(0) <= VN24_sign_out(4);
    CN286_data_in(1) <= VN93_data_out(4);
    CN286_sign_in(1) <= VN93_sign_out(4);
    CN286_data_in(2) <= VN155_data_out(4);
    CN286_sign_in(2) <= VN155_sign_out(4);
    CN286_data_in(3) <= VN189_data_out(4);
    CN286_sign_in(3) <= VN189_sign_out(4);
    CN286_data_in(4) <= VN267_data_out(4);
    CN286_sign_in(4) <= VN267_sign_out(4);
    CN286_data_in(5) <= VN330_data_out(4);
    CN286_sign_in(5) <= VN330_sign_out(4);
    CN286_data_in(6) <= VN341_data_out(4);
    CN286_sign_in(6) <= VN341_sign_out(4);
    CN286_data_in(7) <= VN435_data_out(4);
    CN286_sign_in(7) <= VN435_sign_out(4);
    CN286_data_in(8) <= VN454_data_out(4);
    CN286_sign_in(8) <= VN454_sign_out(4);
    CN286_data_in(9) <= VN556_data_out(4);
    CN286_sign_in(9) <= VN556_sign_out(4);
    CN286_data_in(10) <= VN603_data_out(4);
    CN286_sign_in(10) <= VN603_sign_out(4);
    CN286_data_in(11) <= VN623_data_out(4);
    CN286_sign_in(11) <= VN623_sign_out(4);
    CN286_data_in(12) <= VN688_data_out(4);
    CN286_sign_in(12) <= VN688_sign_out(4);
    CN286_data_in(13) <= VN744_data_out(4);
    CN286_sign_in(13) <= VN744_sign_out(4);
    CN286_data_in(14) <= VN790_data_out(4);
    CN286_sign_in(14) <= VN790_sign_out(4);
    CN286_data_in(15) <= VN842_data_out(4);
    CN286_sign_in(15) <= VN842_sign_out(4);
    CN286_data_in(16) <= VN887_data_out(4);
    CN286_sign_in(16) <= VN887_sign_out(4);
    CN286_data_in(17) <= VN934_data_out(4);
    CN286_sign_in(17) <= VN934_sign_out(4);
    CN286_data_in(18) <= VN975_data_out(4);
    CN286_sign_in(18) <= VN975_sign_out(4);
    CN286_data_in(19) <= VN1005_data_out(4);
    CN286_sign_in(19) <= VN1005_sign_out(4);
    CN286_data_in(20) <= VN1148_data_out(4);
    CN286_sign_in(20) <= VN1148_sign_out(4);
    CN286_data_in(21) <= VN1192_data_out(4);
    CN286_sign_in(21) <= VN1192_sign_out(4);
    CN286_data_in(22) <= VN1254_data_out(4);
    CN286_sign_in(22) <= VN1254_sign_out(4);
    CN286_data_in(23) <= VN1333_data_out(4);
    CN286_sign_in(23) <= VN1333_sign_out(4);
    CN286_data_in(24) <= VN1364_data_out(4);
    CN286_sign_in(24) <= VN1364_sign_out(4);
    CN286_data_in(25) <= VN1507_data_out(4);
    CN286_sign_in(25) <= VN1507_sign_out(4);
    CN286_data_in(26) <= VN1589_data_out(4);
    CN286_sign_in(26) <= VN1589_sign_out(4);
    CN286_data_in(27) <= VN1643_data_out(4);
    CN286_sign_in(27) <= VN1643_sign_out(4);
    CN286_data_in(28) <= VN1659_data_out(4);
    CN286_sign_in(28) <= VN1659_sign_out(4);
    CN286_data_in(29) <= VN1752_data_out(4);
    CN286_sign_in(29) <= VN1752_sign_out(4);
    CN286_data_in(30) <= VN1764_data_out(4);
    CN286_sign_in(30) <= VN1764_sign_out(4);
    CN286_data_in(31) <= VN1866_data_out(4);
    CN286_sign_in(31) <= VN1866_sign_out(4);
    CN287_data_in(0) <= VN23_data_out(4);
    CN287_sign_in(0) <= VN23_sign_out(4);
    CN287_data_in(1) <= VN101_data_out(4);
    CN287_sign_in(1) <= VN101_sign_out(4);
    CN287_data_in(2) <= VN142_data_out(4);
    CN287_sign_in(2) <= VN142_sign_out(4);
    CN287_data_in(3) <= VN193_data_out(4);
    CN287_sign_in(3) <= VN193_sign_out(4);
    CN287_data_in(4) <= VN240_data_out(4);
    CN287_sign_in(4) <= VN240_sign_out(4);
    CN287_data_in(5) <= VN322_data_out(4);
    CN287_sign_in(5) <= VN322_sign_out(4);
    CN287_data_in(6) <= VN375_data_out(4);
    CN287_sign_in(6) <= VN375_sign_out(4);
    CN287_data_in(7) <= VN429_data_out(4);
    CN287_sign_in(7) <= VN429_sign_out(4);
    CN287_data_in(8) <= VN486_data_out(4);
    CN287_sign_in(8) <= VN486_sign_out(4);
    CN287_data_in(9) <= VN514_data_out(4);
    CN287_sign_in(9) <= VN514_sign_out(4);
    CN287_data_in(10) <= VN610_data_out(4);
    CN287_sign_in(10) <= VN610_sign_out(4);
    CN287_data_in(11) <= VN643_data_out(4);
    CN287_sign_in(11) <= VN643_sign_out(4);
    CN287_data_in(12) <= VN716_data_out(4);
    CN287_sign_in(12) <= VN716_sign_out(4);
    CN287_data_in(13) <= VN722_data_out(4);
    CN287_sign_in(13) <= VN722_sign_out(4);
    CN287_data_in(14) <= VN724_data_out(4);
    CN287_sign_in(14) <= VN724_sign_out(4);
    CN287_data_in(15) <= VN784_data_out(4);
    CN287_sign_in(15) <= VN784_sign_out(4);
    CN287_data_in(16) <= VN884_data_out(4);
    CN287_sign_in(16) <= VN884_sign_out(4);
    CN287_data_in(17) <= VN903_data_out(4);
    CN287_sign_in(17) <= VN903_sign_out(4);
    CN287_data_in(18) <= VN981_data_out(4);
    CN287_sign_in(18) <= VN981_sign_out(4);
    CN287_data_in(19) <= VN1028_data_out(4);
    CN287_sign_in(19) <= VN1028_sign_out(4);
    CN287_data_in(20) <= VN1068_data_out(4);
    CN287_sign_in(20) <= VN1068_sign_out(4);
    CN287_data_in(21) <= VN1121_data_out(4);
    CN287_sign_in(21) <= VN1121_sign_out(4);
    CN287_data_in(22) <= VN1188_data_out(4);
    CN287_sign_in(22) <= VN1188_sign_out(4);
    CN287_data_in(23) <= VN1267_data_out(4);
    CN287_sign_in(23) <= VN1267_sign_out(4);
    CN287_data_in(24) <= VN1296_data_out(4);
    CN287_sign_in(24) <= VN1296_sign_out(4);
    CN287_data_in(25) <= VN1334_data_out(4);
    CN287_sign_in(25) <= VN1334_sign_out(4);
    CN287_data_in(26) <= VN1366_data_out(4);
    CN287_sign_in(26) <= VN1366_sign_out(4);
    CN287_data_in(27) <= VN1476_data_out(4);
    CN287_sign_in(27) <= VN1476_sign_out(4);
    CN287_data_in(28) <= VN1551_data_out(4);
    CN287_sign_in(28) <= VN1551_sign_out(4);
    CN287_data_in(29) <= VN1611_data_out(4);
    CN287_sign_in(29) <= VN1611_sign_out(4);
    CN287_data_in(30) <= VN1687_data_out(4);
    CN287_sign_in(30) <= VN1687_sign_out(4);
    CN287_data_in(31) <= VN1793_data_out(4);
    CN287_sign_in(31) <= VN1793_sign_out(4);
    CN288_data_in(0) <= VN22_data_out(4);
    CN288_sign_in(0) <= VN22_sign_out(4);
    CN288_data_in(1) <= VN75_data_out(4);
    CN288_sign_in(1) <= VN75_sign_out(4);
    CN288_data_in(2) <= VN161_data_out(4);
    CN288_sign_in(2) <= VN161_sign_out(4);
    CN288_data_in(3) <= VN224_data_out(4);
    CN288_sign_in(3) <= VN224_sign_out(4);
    CN288_data_in(4) <= VN228_data_out(4);
    CN288_sign_in(4) <= VN228_sign_out(4);
    CN288_data_in(5) <= VN308_data_out(4);
    CN288_sign_in(5) <= VN308_sign_out(4);
    CN288_data_in(6) <= VN337_data_out(4);
    CN288_sign_in(6) <= VN337_sign_out(4);
    CN288_data_in(7) <= VN410_data_out(4);
    CN288_sign_in(7) <= VN410_sign_out(4);
    CN288_data_in(8) <= VN468_data_out(4);
    CN288_sign_in(8) <= VN468_sign_out(4);
    CN288_data_in(9) <= VN542_data_out(4);
    CN288_sign_in(9) <= VN542_sign_out(4);
    CN288_data_in(10) <= VN578_data_out(4);
    CN288_sign_in(10) <= VN578_sign_out(4);
    CN288_data_in(11) <= VN644_data_out(4);
    CN288_sign_in(11) <= VN644_sign_out(4);
    CN288_data_in(12) <= VN695_data_out(4);
    CN288_sign_in(12) <= VN695_sign_out(4);
    CN288_data_in(13) <= VN763_data_out(4);
    CN288_sign_in(13) <= VN763_sign_out(4);
    CN288_data_in(14) <= VN787_data_out(4);
    CN288_sign_in(14) <= VN787_sign_out(4);
    CN288_data_in(15) <= VN845_data_out(4);
    CN288_sign_in(15) <= VN845_sign_out(4);
    CN288_data_in(16) <= VN916_data_out(4);
    CN288_sign_in(16) <= VN916_sign_out(4);
    CN288_data_in(17) <= VN964_data_out(4);
    CN288_sign_in(17) <= VN964_sign_out(4);
    CN288_data_in(18) <= VN1010_data_out(4);
    CN288_sign_in(18) <= VN1010_sign_out(4);
    CN288_data_in(19) <= VN1061_data_out(4);
    CN288_sign_in(19) <= VN1061_sign_out(4);
    CN288_data_in(20) <= VN1135_data_out(4);
    CN288_sign_in(20) <= VN1135_sign_out(4);
    CN288_data_in(21) <= VN1168_data_out(4);
    CN288_sign_in(21) <= VN1168_sign_out(4);
    CN288_data_in(22) <= VN1206_data_out(4);
    CN288_sign_in(22) <= VN1206_sign_out(4);
    CN288_data_in(23) <= VN1263_data_out(4);
    CN288_sign_in(23) <= VN1263_sign_out(4);
    CN288_data_in(24) <= VN1324_data_out(4);
    CN288_sign_in(24) <= VN1324_sign_out(4);
    CN288_data_in(25) <= VN1405_data_out(4);
    CN288_sign_in(25) <= VN1405_sign_out(4);
    CN288_data_in(26) <= VN1473_data_out(4);
    CN288_sign_in(26) <= VN1473_sign_out(4);
    CN288_data_in(27) <= VN1487_data_out(4);
    CN288_sign_in(27) <= VN1487_sign_out(4);
    CN288_data_in(28) <= VN1619_data_out(4);
    CN288_sign_in(28) <= VN1619_sign_out(4);
    CN288_data_in(29) <= VN1658_data_out(4);
    CN288_sign_in(29) <= VN1658_sign_out(4);
    CN288_data_in(30) <= VN1713_data_out(4);
    CN288_sign_in(30) <= VN1713_sign_out(4);
    CN288_data_in(31) <= VN1794_data_out(4);
    CN288_sign_in(31) <= VN1794_sign_out(4);
    CN289_data_in(0) <= VN21_data_out(4);
    CN289_sign_in(0) <= VN21_sign_out(4);
    CN289_data_in(1) <= VN89_data_out(4);
    CN289_sign_in(1) <= VN89_sign_out(4);
    CN289_data_in(2) <= VN134_data_out(4);
    CN289_sign_in(2) <= VN134_sign_out(4);
    CN289_data_in(3) <= VN192_data_out(4);
    CN289_sign_in(3) <= VN192_sign_out(4);
    CN289_data_in(4) <= VN269_data_out(4);
    CN289_sign_in(4) <= VN269_sign_out(4);
    CN289_data_in(5) <= VN327_data_out(4);
    CN289_sign_in(5) <= VN327_sign_out(4);
    CN289_data_in(6) <= VN365_data_out(4);
    CN289_sign_in(6) <= VN365_sign_out(4);
    CN289_data_in(7) <= VN418_data_out(4);
    CN289_sign_in(7) <= VN418_sign_out(4);
    CN289_data_in(8) <= VN471_data_out(4);
    CN289_sign_in(8) <= VN471_sign_out(4);
    CN289_data_in(9) <= VN519_data_out(4);
    CN289_sign_in(9) <= VN519_sign_out(4);
    CN289_data_in(10) <= VN577_data_out(4);
    CN289_sign_in(10) <= VN577_sign_out(4);
    CN289_data_in(11) <= VN622_data_out(4);
    CN289_sign_in(11) <= VN622_sign_out(4);
    CN289_data_in(12) <= VN717_data_out(4);
    CN289_sign_in(12) <= VN717_sign_out(4);
    CN289_data_in(13) <= VN774_data_out(4);
    CN289_sign_in(13) <= VN774_sign_out(4);
    CN289_data_in(14) <= VN778_data_out(4);
    CN289_sign_in(14) <= VN778_sign_out(4);
    CN289_data_in(15) <= VN913_data_out(4);
    CN289_sign_in(15) <= VN913_sign_out(4);
    CN289_data_in(16) <= VN966_data_out(4);
    CN289_sign_in(16) <= VN966_sign_out(4);
    CN289_data_in(17) <= VN1021_data_out(4);
    CN289_sign_in(17) <= VN1021_sign_out(4);
    CN289_data_in(18) <= VN1065_data_out(4);
    CN289_sign_in(18) <= VN1065_sign_out(4);
    CN289_data_in(19) <= VN1110_data_out(4);
    CN289_sign_in(19) <= VN1110_sign_out(4);
    CN289_data_in(20) <= VN1173_data_out(4);
    CN289_sign_in(20) <= VN1173_sign_out(4);
    CN289_data_in(21) <= VN1227_data_out(4);
    CN289_sign_in(21) <= VN1227_sign_out(4);
    CN289_data_in(22) <= VN1283_data_out(4);
    CN289_sign_in(22) <= VN1283_sign_out(4);
    CN289_data_in(23) <= VN1372_data_out(4);
    CN289_sign_in(23) <= VN1372_sign_out(4);
    CN289_data_in(24) <= VN1410_data_out(4);
    CN289_sign_in(24) <= VN1410_sign_out(4);
    CN289_data_in(25) <= VN1441_data_out(4);
    CN289_sign_in(25) <= VN1441_sign_out(4);
    CN289_data_in(26) <= VN1479_data_out(4);
    CN289_sign_in(26) <= VN1479_sign_out(4);
    CN289_data_in(27) <= VN1510_data_out(4);
    CN289_sign_in(27) <= VN1510_sign_out(4);
    CN289_data_in(28) <= VN1614_data_out(4);
    CN289_sign_in(28) <= VN1614_sign_out(4);
    CN289_data_in(29) <= VN1654_data_out(4);
    CN289_sign_in(29) <= VN1654_sign_out(4);
    CN289_data_in(30) <= VN1994_data_out(4);
    CN289_sign_in(30) <= VN1994_sign_out(4);
    CN289_data_in(31) <= VN1998_data_out(4);
    CN289_sign_in(31) <= VN1998_sign_out(4);
    CN290_data_in(0) <= VN20_data_out(4);
    CN290_sign_in(0) <= VN20_sign_out(4);
    CN290_data_in(1) <= VN60_data_out(4);
    CN290_sign_in(1) <= VN60_sign_out(4);
    CN290_data_in(2) <= VN131_data_out(4);
    CN290_sign_in(2) <= VN131_sign_out(4);
    CN290_data_in(3) <= VN187_data_out(4);
    CN290_sign_in(3) <= VN187_sign_out(4);
    CN290_data_in(4) <= VN231_data_out(4);
    CN290_sign_in(4) <= VN231_sign_out(4);
    CN290_data_in(5) <= VN350_data_out(4);
    CN290_sign_in(5) <= VN350_sign_out(4);
    CN290_data_in(6) <= VN440_data_out(4);
    CN290_sign_in(6) <= VN440_sign_out(4);
    CN290_data_in(7) <= VN457_data_out(4);
    CN290_sign_in(7) <= VN457_sign_out(4);
    CN290_data_in(8) <= VN544_data_out(4);
    CN290_sign_in(8) <= VN544_sign_out(4);
    CN290_data_in(9) <= VN608_data_out(4);
    CN290_sign_in(9) <= VN608_sign_out(4);
    CN290_data_in(10) <= VN676_data_out(4);
    CN290_sign_in(10) <= VN676_sign_out(4);
    CN290_data_in(11) <= VN730_data_out(4);
    CN290_sign_in(11) <= VN730_sign_out(4);
    CN290_data_in(12) <= VN811_data_out(4);
    CN290_sign_in(12) <= VN811_sign_out(4);
    CN290_data_in(13) <= VN872_data_out(4);
    CN290_sign_in(13) <= VN872_sign_out(4);
    CN290_data_in(14) <= VN992_data_out(4);
    CN290_sign_in(14) <= VN992_sign_out(4);
    CN290_data_in(15) <= VN1107_data_out(4);
    CN290_sign_in(15) <= VN1107_sign_out(4);
    CN290_data_in(16) <= VN1142_data_out(4);
    CN290_sign_in(16) <= VN1142_sign_out(4);
    CN290_data_in(17) <= VN1174_data_out(4);
    CN290_sign_in(17) <= VN1174_sign_out(4);
    CN290_data_in(18) <= VN1247_data_out(4);
    CN290_sign_in(18) <= VN1247_sign_out(4);
    CN290_data_in(19) <= VN1328_data_out(4);
    CN290_sign_in(19) <= VN1328_sign_out(4);
    CN290_data_in(20) <= VN1483_data_out(4);
    CN290_sign_in(20) <= VN1483_sign_out(4);
    CN290_data_in(21) <= VN1552_data_out(4);
    CN290_sign_in(21) <= VN1552_sign_out(4);
    CN290_data_in(22) <= VN1558_data_out(4);
    CN290_sign_in(22) <= VN1558_sign_out(4);
    CN290_data_in(23) <= VN1563_data_out(4);
    CN290_sign_in(23) <= VN1563_sign_out(4);
    CN290_data_in(24) <= VN1620_data_out(4);
    CN290_sign_in(24) <= VN1620_sign_out(4);
    CN290_data_in(25) <= VN1712_data_out(4);
    CN290_sign_in(25) <= VN1712_sign_out(4);
    CN290_data_in(26) <= VN1783_data_out(4);
    CN290_sign_in(26) <= VN1783_sign_out(4);
    CN290_data_in(27) <= VN1820_data_out(4);
    CN290_sign_in(27) <= VN1820_sign_out(4);
    CN290_data_in(28) <= VN1850_data_out(4);
    CN290_sign_in(28) <= VN1850_sign_out(4);
    CN290_data_in(29) <= VN1886_data_out(4);
    CN290_sign_in(29) <= VN1886_sign_out(4);
    CN290_data_in(30) <= VN1972_data_out(4);
    CN290_sign_in(30) <= VN1972_sign_out(4);
    CN290_data_in(31) <= VN1977_data_out(4);
    CN290_sign_in(31) <= VN1977_sign_out(4);
    CN291_data_in(0) <= VN19_data_out(4);
    CN291_sign_in(0) <= VN19_sign_out(4);
    CN291_data_in(1) <= VN96_data_out(4);
    CN291_sign_in(1) <= VN96_sign_out(4);
    CN291_data_in(2) <= VN147_data_out(4);
    CN291_sign_in(2) <= VN147_sign_out(4);
    CN291_data_in(3) <= VN223_data_out(4);
    CN291_sign_in(3) <= VN223_sign_out(4);
    CN291_data_in(4) <= VN249_data_out(4);
    CN291_sign_in(4) <= VN249_sign_out(4);
    CN291_data_in(5) <= VN377_data_out(4);
    CN291_sign_in(5) <= VN377_sign_out(4);
    CN291_data_in(6) <= VN439_data_out(4);
    CN291_sign_in(6) <= VN439_sign_out(4);
    CN291_data_in(7) <= VN487_data_out(4);
    CN291_sign_in(7) <= VN487_sign_out(4);
    CN291_data_in(8) <= VN558_data_out(4);
    CN291_sign_in(8) <= VN558_sign_out(4);
    CN291_data_in(9) <= VN590_data_out(4);
    CN291_sign_in(9) <= VN590_sign_out(4);
    CN291_data_in(10) <= VN629_data_out(4);
    CN291_sign_in(10) <= VN629_sign_out(4);
    CN291_data_in(11) <= VN673_data_out(4);
    CN291_sign_in(11) <= VN673_sign_out(4);
    CN291_data_in(12) <= VN757_data_out(4);
    CN291_sign_in(12) <= VN757_sign_out(4);
    CN291_data_in(13) <= VN796_data_out(4);
    CN291_sign_in(13) <= VN796_sign_out(4);
    CN291_data_in(14) <= VN867_data_out(4);
    CN291_sign_in(14) <= VN867_sign_out(4);
    CN291_data_in(15) <= VN896_data_out(4);
    CN291_sign_in(15) <= VN896_sign_out(4);
    CN291_data_in(16) <= VN973_data_out(4);
    CN291_sign_in(16) <= VN973_sign_out(4);
    CN291_data_in(17) <= VN1004_data_out(4);
    CN291_sign_in(17) <= VN1004_sign_out(4);
    CN291_data_in(18) <= VN1089_data_out(4);
    CN291_sign_in(18) <= VN1089_sign_out(4);
    CN291_data_in(19) <= VN1205_data_out(4);
    CN291_sign_in(19) <= VN1205_sign_out(4);
    CN291_data_in(20) <= VN1248_data_out(4);
    CN291_sign_in(20) <= VN1248_sign_out(4);
    CN291_data_in(21) <= VN1336_data_out(4);
    CN291_sign_in(21) <= VN1336_sign_out(4);
    CN291_data_in(22) <= VN1409_data_out(4);
    CN291_sign_in(22) <= VN1409_sign_out(4);
    CN291_data_in(23) <= VN1450_data_out(4);
    CN291_sign_in(23) <= VN1450_sign_out(4);
    CN291_data_in(24) <= VN1465_data_out(4);
    CN291_sign_in(24) <= VN1465_sign_out(4);
    CN291_data_in(25) <= VN1494_data_out(4);
    CN291_sign_in(25) <= VN1494_sign_out(4);
    CN291_data_in(26) <= VN1512_data_out(4);
    CN291_sign_in(26) <= VN1512_sign_out(4);
    CN291_data_in(27) <= VN1529_data_out(4);
    CN291_sign_in(27) <= VN1529_sign_out(4);
    CN291_data_in(28) <= VN1568_data_out(4);
    CN291_sign_in(28) <= VN1568_sign_out(4);
    CN291_data_in(29) <= VN1610_data_out(4);
    CN291_sign_in(29) <= VN1610_sign_out(4);
    CN291_data_in(30) <= VN1767_data_out(4);
    CN291_sign_in(30) <= VN1767_sign_out(4);
    CN291_data_in(31) <= VN1867_data_out(4);
    CN291_sign_in(31) <= VN1867_sign_out(4);
    CN292_data_in(0) <= VN18_data_out(4);
    CN292_sign_in(0) <= VN18_sign_out(4);
    CN292_data_in(1) <= VN62_data_out(4);
    CN292_sign_in(1) <= VN62_sign_out(4);
    CN292_data_in(2) <= VN139_data_out(4);
    CN292_sign_in(2) <= VN139_sign_out(4);
    CN292_data_in(3) <= VN177_data_out(4);
    CN292_sign_in(3) <= VN177_sign_out(4);
    CN292_data_in(4) <= VN257_data_out(4);
    CN292_sign_in(4) <= VN257_sign_out(4);
    CN292_data_in(5) <= VN313_data_out(4);
    CN292_sign_in(5) <= VN313_sign_out(4);
    CN292_data_in(6) <= VN367_data_out(4);
    CN292_sign_in(6) <= VN367_sign_out(4);
    CN292_data_in(7) <= VN416_data_out(4);
    CN292_sign_in(7) <= VN416_sign_out(4);
    CN292_data_in(8) <= VN453_data_out(4);
    CN292_sign_in(8) <= VN453_sign_out(4);
    CN292_data_in(9) <= VN554_data_out(4);
    CN292_sign_in(9) <= VN554_sign_out(4);
    CN292_data_in(10) <= VN592_data_out(4);
    CN292_sign_in(10) <= VN592_sign_out(4);
    CN292_data_in(11) <= VN633_data_out(4);
    CN292_sign_in(11) <= VN633_sign_out(4);
    CN292_data_in(12) <= VN690_data_out(4);
    CN292_sign_in(12) <= VN690_sign_out(4);
    CN292_data_in(13) <= VN745_data_out(4);
    CN292_sign_in(13) <= VN745_sign_out(4);
    CN292_data_in(14) <= VN806_data_out(4);
    CN292_sign_in(14) <= VN806_sign_out(4);
    CN292_data_in(15) <= VN873_data_out(4);
    CN292_sign_in(15) <= VN873_sign_out(4);
    CN292_data_in(16) <= VN897_data_out(4);
    CN292_sign_in(16) <= VN897_sign_out(4);
    CN292_data_in(17) <= VN985_data_out(4);
    CN292_sign_in(17) <= VN985_sign_out(4);
    CN292_data_in(18) <= VN1017_data_out(4);
    CN292_sign_in(18) <= VN1017_sign_out(4);
    CN292_data_in(19) <= VN1074_data_out(4);
    CN292_sign_in(19) <= VN1074_sign_out(4);
    CN292_data_in(20) <= VN1122_data_out(4);
    CN292_sign_in(20) <= VN1122_sign_out(4);
    CN292_data_in(21) <= VN1197_data_out(4);
    CN292_sign_in(21) <= VN1197_sign_out(4);
    CN292_data_in(22) <= VN1226_data_out(4);
    CN292_sign_in(22) <= VN1226_sign_out(4);
    CN292_data_in(23) <= VN1321_data_out(4);
    CN292_sign_in(23) <= VN1321_sign_out(4);
    CN292_data_in(24) <= VN1365_data_out(4);
    CN292_sign_in(24) <= VN1365_sign_out(4);
    CN292_data_in(25) <= VN1403_data_out(4);
    CN292_sign_in(25) <= VN1403_sign_out(4);
    CN292_data_in(26) <= VN1575_data_out(4);
    CN292_sign_in(26) <= VN1575_sign_out(4);
    CN292_data_in(27) <= VN1594_data_out(4);
    CN292_sign_in(27) <= VN1594_sign_out(4);
    CN292_data_in(28) <= VN1630_data_out(4);
    CN292_sign_in(28) <= VN1630_sign_out(4);
    CN292_data_in(29) <= VN1663_data_out(4);
    CN292_sign_in(29) <= VN1663_sign_out(4);
    CN292_data_in(30) <= VN1705_data_out(4);
    CN292_sign_in(30) <= VN1705_sign_out(4);
    CN292_data_in(31) <= VN1795_data_out(4);
    CN292_sign_in(31) <= VN1795_sign_out(4);
    CN293_data_in(0) <= VN17_data_out(4);
    CN293_sign_in(0) <= VN17_sign_out(4);
    CN293_data_in(1) <= VN77_data_out(4);
    CN293_sign_in(1) <= VN77_sign_out(4);
    CN293_data_in(2) <= VN113_data_out(4);
    CN293_sign_in(2) <= VN113_sign_out(4);
    CN293_data_in(3) <= VN197_data_out(4);
    CN293_sign_in(3) <= VN197_sign_out(4);
    CN293_data_in(4) <= VN306_data_out(4);
    CN293_sign_in(4) <= VN306_sign_out(4);
    CN293_data_in(5) <= VN354_data_out(4);
    CN293_sign_in(5) <= VN354_sign_out(4);
    CN293_data_in(6) <= VN397_data_out(4);
    CN293_sign_in(6) <= VN397_sign_out(4);
    CN293_data_in(7) <= VN479_data_out(4);
    CN293_sign_in(7) <= VN479_sign_out(4);
    CN293_data_in(8) <= VN516_data_out(4);
    CN293_sign_in(8) <= VN516_sign_out(4);
    CN293_data_in(9) <= VN579_data_out(4);
    CN293_sign_in(9) <= VN579_sign_out(4);
    CN293_data_in(10) <= VN668_data_out(4);
    CN293_sign_in(10) <= VN668_sign_out(4);
    CN293_data_in(11) <= VN712_data_out(4);
    CN293_sign_in(11) <= VN712_sign_out(4);
    CN293_data_in(12) <= VN732_data_out(4);
    CN293_sign_in(12) <= VN732_sign_out(4);
    CN293_data_in(13) <= VN818_data_out(4);
    CN293_sign_in(13) <= VN818_sign_out(4);
    CN293_data_in(14) <= VN864_data_out(4);
    CN293_sign_in(14) <= VN864_sign_out(4);
    CN293_data_in(15) <= VN930_data_out(4);
    CN293_sign_in(15) <= VN930_sign_out(4);
    CN293_data_in(16) <= VN993_data_out(4);
    CN293_sign_in(16) <= VN993_sign_out(4);
    CN293_data_in(17) <= VN1045_data_out(4);
    CN293_sign_in(17) <= VN1045_sign_out(4);
    CN293_data_in(18) <= VN1085_data_out(4);
    CN293_sign_in(18) <= VN1085_sign_out(4);
    CN293_data_in(19) <= VN1119_data_out(4);
    CN293_sign_in(19) <= VN1119_sign_out(4);
    CN293_data_in(20) <= VN1214_data_out(4);
    CN293_sign_in(20) <= VN1214_sign_out(4);
    CN293_data_in(21) <= VN1274_data_out(4);
    CN293_sign_in(21) <= VN1274_sign_out(4);
    CN293_data_in(22) <= VN1302_data_out(4);
    CN293_sign_in(22) <= VN1302_sign_out(4);
    CN293_data_in(23) <= VN1379_data_out(4);
    CN293_sign_in(23) <= VN1379_sign_out(4);
    CN293_data_in(24) <= VN1448_data_out(4);
    CN293_sign_in(24) <= VN1448_sign_out(4);
    CN293_data_in(25) <= VN1548_data_out(4);
    CN293_sign_in(25) <= VN1548_sign_out(4);
    CN293_data_in(26) <= VN1567_data_out(4);
    CN293_sign_in(26) <= VN1567_sign_out(4);
    CN293_data_in(27) <= VN1582_data_out(4);
    CN293_sign_in(27) <= VN1582_sign_out(4);
    CN293_data_in(28) <= VN1636_data_out(4);
    CN293_sign_in(28) <= VN1636_sign_out(4);
    CN293_data_in(29) <= VN1662_data_out(4);
    CN293_sign_in(29) <= VN1662_sign_out(4);
    CN293_data_in(30) <= VN1696_data_out(4);
    CN293_sign_in(30) <= VN1696_sign_out(4);
    CN293_data_in(31) <= VN1796_data_out(4);
    CN293_sign_in(31) <= VN1796_sign_out(4);
    CN294_data_in(0) <= VN16_data_out(4);
    CN294_sign_in(0) <= VN16_sign_out(4);
    CN294_data_in(1) <= VN73_data_out(4);
    CN294_sign_in(1) <= VN73_sign_out(4);
    CN294_data_in(2) <= VN123_data_out(4);
    CN294_sign_in(2) <= VN123_sign_out(4);
    CN294_data_in(3) <= VN196_data_out(4);
    CN294_sign_in(3) <= VN196_sign_out(4);
    CN294_data_in(4) <= VN258_data_out(4);
    CN294_sign_in(4) <= VN258_sign_out(4);
    CN294_data_in(5) <= VN284_data_out(4);
    CN294_sign_in(5) <= VN284_sign_out(4);
    CN294_data_in(6) <= VN373_data_out(4);
    CN294_sign_in(6) <= VN373_sign_out(4);
    CN294_data_in(7) <= VN400_data_out(4);
    CN294_sign_in(7) <= VN400_sign_out(4);
    CN294_data_in(8) <= VN465_data_out(4);
    CN294_sign_in(8) <= VN465_sign_out(4);
    CN294_data_in(9) <= VN537_data_out(4);
    CN294_sign_in(9) <= VN537_sign_out(4);
    CN294_data_in(10) <= VN609_data_out(4);
    CN294_sign_in(10) <= VN609_sign_out(4);
    CN294_data_in(11) <= VN632_data_out(4);
    CN294_sign_in(11) <= VN632_sign_out(4);
    CN294_data_in(12) <= VN713_data_out(4);
    CN294_sign_in(12) <= VN713_sign_out(4);
    CN294_data_in(13) <= VN748_data_out(4);
    CN294_sign_in(13) <= VN748_sign_out(4);
    CN294_data_in(14) <= VN791_data_out(4);
    CN294_sign_in(14) <= VN791_sign_out(4);
    CN294_data_in(15) <= VN831_data_out(4);
    CN294_sign_in(15) <= VN831_sign_out(4);
    CN294_data_in(16) <= VN922_data_out(4);
    CN294_sign_in(16) <= VN922_sign_out(4);
    CN294_data_in(17) <= VN965_data_out(4);
    CN294_sign_in(17) <= VN965_sign_out(4);
    CN294_data_in(18) <= VN1024_data_out(4);
    CN294_sign_in(18) <= VN1024_sign_out(4);
    CN294_data_in(19) <= VN1094_data_out(4);
    CN294_sign_in(19) <= VN1094_sign_out(4);
    CN294_data_in(20) <= VN1138_data_out(4);
    CN294_sign_in(20) <= VN1138_sign_out(4);
    CN294_data_in(21) <= VN1217_data_out(4);
    CN294_sign_in(21) <= VN1217_sign_out(4);
    CN294_data_in(22) <= VN1235_data_out(4);
    CN294_sign_in(22) <= VN1235_sign_out(4);
    CN294_data_in(23) <= VN1287_data_out(4);
    CN294_sign_in(23) <= VN1287_sign_out(4);
    CN294_data_in(24) <= VN1353_data_out(4);
    CN294_sign_in(24) <= VN1353_sign_out(4);
    CN294_data_in(25) <= VN1393_data_out(4);
    CN294_sign_in(25) <= VN1393_sign_out(4);
    CN294_data_in(26) <= VN1555_data_out(4);
    CN294_sign_in(26) <= VN1555_sign_out(4);
    CN294_data_in(27) <= VN1562_data_out(4);
    CN294_sign_in(27) <= VN1562_sign_out(4);
    CN294_data_in(28) <= VN1624_data_out(4);
    CN294_sign_in(28) <= VN1624_sign_out(4);
    CN294_data_in(29) <= VN1686_data_out(4);
    CN294_sign_in(29) <= VN1686_sign_out(4);
    CN294_data_in(30) <= VN1689_data_out(4);
    CN294_sign_in(30) <= VN1689_sign_out(4);
    CN294_data_in(31) <= VN1797_data_out(4);
    CN294_sign_in(31) <= VN1797_sign_out(4);
    CN295_data_in(0) <= VN15_data_out(4);
    CN295_sign_in(0) <= VN15_sign_out(4);
    CN295_data_in(1) <= VN92_data_out(4);
    CN295_sign_in(1) <= VN92_sign_out(4);
    CN295_data_in(2) <= VN117_data_out(4);
    CN295_sign_in(2) <= VN117_sign_out(4);
    CN295_data_in(3) <= VN175_data_out(4);
    CN295_sign_in(3) <= VN175_sign_out(4);
    CN295_data_in(4) <= VN346_data_out(4);
    CN295_sign_in(4) <= VN346_sign_out(4);
    CN295_data_in(5) <= VN441_data_out(4);
    CN295_sign_in(5) <= VN441_sign_out(4);
    CN295_data_in(6) <= VN489_data_out(4);
    CN295_sign_in(6) <= VN489_sign_out(4);
    CN295_data_in(7) <= VN538_data_out(4);
    CN295_sign_in(7) <= VN538_sign_out(4);
    CN295_data_in(8) <= VN576_data_out(4);
    CN295_sign_in(8) <= VN576_sign_out(4);
    CN295_data_in(9) <= VN628_data_out(4);
    CN295_sign_in(9) <= VN628_sign_out(4);
    CN295_data_in(10) <= VN768_data_out(4);
    CN295_sign_in(10) <= VN768_sign_out(4);
    CN295_data_in(11) <= VN837_data_out(4);
    CN295_sign_in(11) <= VN837_sign_out(4);
    CN295_data_in(12) <= VN938_data_out(4);
    CN295_sign_in(12) <= VN938_sign_out(4);
    CN295_data_in(13) <= VN1047_data_out(4);
    CN295_sign_in(13) <= VN1047_sign_out(4);
    CN295_data_in(14) <= VN1160_data_out(4);
    CN295_sign_in(14) <= VN1160_sign_out(4);
    CN295_data_in(15) <= VN1169_data_out(4);
    CN295_sign_in(15) <= VN1169_sign_out(4);
    CN295_data_in(16) <= VN1299_data_out(4);
    CN295_sign_in(16) <= VN1299_sign_out(4);
    CN295_data_in(17) <= VN1415_data_out(4);
    CN295_sign_in(17) <= VN1415_sign_out(4);
    CN295_data_in(18) <= VN1439_data_out(4);
    CN295_sign_in(18) <= VN1439_sign_out(4);
    CN295_data_in(19) <= VN1519_data_out(4);
    CN295_sign_in(19) <= VN1519_sign_out(4);
    CN295_data_in(20) <= VN1535_data_out(4);
    CN295_sign_in(20) <= VN1535_sign_out(4);
    CN295_data_in(21) <= VN1670_data_out(4);
    CN295_sign_in(21) <= VN1670_sign_out(4);
    CN295_data_in(22) <= VN1699_data_out(4);
    CN295_sign_in(22) <= VN1699_sign_out(4);
    CN295_data_in(23) <= VN1737_data_out(4);
    CN295_sign_in(23) <= VN1737_sign_out(4);
    CN295_data_in(24) <= VN1756_data_out(4);
    CN295_sign_in(24) <= VN1756_sign_out(4);
    CN295_data_in(25) <= VN1826_data_out(4);
    CN295_sign_in(25) <= VN1826_sign_out(4);
    CN295_data_in(26) <= VN1843_data_out(4);
    CN295_sign_in(26) <= VN1843_sign_out(4);
    CN295_data_in(27) <= VN1931_data_out(4);
    CN295_sign_in(27) <= VN1931_sign_out(4);
    CN295_data_in(28) <= VN1975_data_out(4);
    CN295_sign_in(28) <= VN1975_sign_out(4);
    CN295_data_in(29) <= VN1982_data_out(4);
    CN295_sign_in(29) <= VN1982_sign_out(4);
    CN295_data_in(30) <= VN1987_data_out(4);
    CN295_sign_in(30) <= VN1987_sign_out(4);
    CN295_data_in(31) <= VN1989_data_out(4);
    CN295_sign_in(31) <= VN1989_sign_out(4);
    CN296_data_in(0) <= VN14_data_out(4);
    CN296_sign_in(0) <= VN14_sign_out(4);
    CN296_data_in(1) <= VN55_data_out(4);
    CN296_sign_in(1) <= VN55_sign_out(4);
    CN296_data_in(2) <= VN121_data_out(4);
    CN296_sign_in(2) <= VN121_sign_out(4);
    CN296_data_in(3) <= VN208_data_out(4);
    CN296_sign_in(3) <= VN208_sign_out(4);
    CN296_data_in(4) <= VN286_data_out(4);
    CN296_sign_in(4) <= VN286_sign_out(4);
    CN296_data_in(5) <= VN343_data_out(4);
    CN296_sign_in(5) <= VN343_sign_out(4);
    CN296_data_in(6) <= VN417_data_out(4);
    CN296_sign_in(6) <= VN417_sign_out(4);
    CN296_data_in(7) <= VN481_data_out(4);
    CN296_sign_in(7) <= VN481_sign_out(4);
    CN296_data_in(8) <= VN515_data_out(4);
    CN296_sign_in(8) <= VN515_sign_out(4);
    CN296_data_in(9) <= VN665_data_out(4);
    CN296_sign_in(9) <= VN665_sign_out(4);
    CN296_data_in(10) <= VN681_data_out(4);
    CN296_sign_in(10) <= VN681_sign_out(4);
    CN296_data_in(11) <= VN820_data_out(4);
    CN296_sign_in(11) <= VN820_sign_out(4);
    CN296_data_in(12) <= VN951_data_out(4);
    CN296_sign_in(12) <= VN951_sign_out(4);
    CN296_data_in(13) <= VN1109_data_out(4);
    CN296_sign_in(13) <= VN1109_sign_out(4);
    CN296_data_in(14) <= VN1161_data_out(4);
    CN296_sign_in(14) <= VN1161_sign_out(4);
    CN296_data_in(15) <= VN1216_data_out(4);
    CN296_sign_in(15) <= VN1216_sign_out(4);
    CN296_data_in(16) <= VN1307_data_out(4);
    CN296_sign_in(16) <= VN1307_sign_out(4);
    CN296_data_in(17) <= VN1413_data_out(4);
    CN296_sign_in(17) <= VN1413_sign_out(4);
    CN296_data_in(18) <= VN1469_data_out(4);
    CN296_sign_in(18) <= VN1469_sign_out(4);
    CN296_data_in(19) <= VN1525_data_out(4);
    CN296_sign_in(19) <= VN1525_sign_out(4);
    CN296_data_in(20) <= VN1577_data_out(4);
    CN296_sign_in(20) <= VN1577_sign_out(4);
    CN296_data_in(21) <= VN1646_data_out(4);
    CN296_sign_in(21) <= VN1646_sign_out(4);
    CN296_data_in(22) <= VN1671_data_out(4);
    CN296_sign_in(22) <= VN1671_sign_out(4);
    CN296_data_in(23) <= VN1832_data_out(4);
    CN296_sign_in(23) <= VN1832_sign_out(4);
    CN296_data_in(24) <= VN1838_data_out(4);
    CN296_sign_in(24) <= VN1838_sign_out(4);
    CN296_data_in(25) <= VN1880_data_out(4);
    CN296_sign_in(25) <= VN1880_sign_out(4);
    CN296_data_in(26) <= VN1882_data_out(4);
    CN296_sign_in(26) <= VN1882_sign_out(4);
    CN296_data_in(27) <= VN1897_data_out(4);
    CN296_sign_in(27) <= VN1897_sign_out(4);
    CN296_data_in(28) <= VN1902_data_out(4);
    CN296_sign_in(28) <= VN1902_sign_out(4);
    CN296_data_in(29) <= VN1933_data_out(4);
    CN296_sign_in(29) <= VN1933_sign_out(4);
    CN296_data_in(30) <= VN1950_data_out(4);
    CN296_sign_in(30) <= VN1950_sign_out(4);
    CN296_data_in(31) <= VN1956_data_out(4);
    CN296_sign_in(31) <= VN1956_sign_out(4);
    CN297_data_in(0) <= VN13_data_out(4);
    CN297_sign_in(0) <= VN13_sign_out(4);
    CN297_data_in(1) <= VN56_data_out(4);
    CN297_sign_in(1) <= VN56_sign_out(4);
    CN297_data_in(2) <= VN111_data_out(4);
    CN297_sign_in(2) <= VN111_sign_out(4);
    CN297_data_in(3) <= VN211_data_out(4);
    CN297_sign_in(3) <= VN211_sign_out(4);
    CN297_data_in(4) <= VN277_data_out(4);
    CN297_sign_in(4) <= VN277_sign_out(4);
    CN297_data_in(5) <= VN290_data_out(4);
    CN297_sign_in(5) <= VN290_sign_out(4);
    CN297_data_in(6) <= VN358_data_out(4);
    CN297_sign_in(6) <= VN358_sign_out(4);
    CN297_data_in(7) <= VN438_data_out(4);
    CN297_sign_in(7) <= VN438_sign_out(4);
    CN297_data_in(8) <= VN469_data_out(4);
    CN297_sign_in(8) <= VN469_sign_out(4);
    CN297_data_in(9) <= VN508_data_out(4);
    CN297_sign_in(9) <= VN508_sign_out(4);
    CN297_data_in(10) <= VN587_data_out(4);
    CN297_sign_in(10) <= VN587_sign_out(4);
    CN297_data_in(11) <= VN620_data_out(4);
    CN297_sign_in(11) <= VN620_sign_out(4);
    CN297_data_in(12) <= VN699_data_out(4);
    CN297_sign_in(12) <= VN699_sign_out(4);
    CN297_data_in(13) <= VN772_data_out(4);
    CN297_sign_in(13) <= VN772_sign_out(4);
    CN297_data_in(14) <= VN782_data_out(4);
    CN297_sign_in(14) <= VN782_sign_out(4);
    CN297_data_in(15) <= VN878_data_out(4);
    CN297_sign_in(15) <= VN878_sign_out(4);
    CN297_data_in(16) <= VN988_data_out(4);
    CN297_sign_in(16) <= VN988_sign_out(4);
    CN297_data_in(17) <= VN1058_data_out(4);
    CN297_sign_in(17) <= VN1058_sign_out(4);
    CN297_data_in(18) <= VN1096_data_out(4);
    CN297_sign_in(18) <= VN1096_sign_out(4);
    CN297_data_in(19) <= VN1137_data_out(4);
    CN297_sign_in(19) <= VN1137_sign_out(4);
    CN297_data_in(20) <= VN1165_data_out(4);
    CN297_sign_in(20) <= VN1165_sign_out(4);
    CN297_data_in(21) <= VN1239_data_out(4);
    CN297_sign_in(21) <= VN1239_sign_out(4);
    CN297_data_in(22) <= VN1284_data_out(4);
    CN297_sign_in(22) <= VN1284_sign_out(4);
    CN297_data_in(23) <= VN1367_data_out(4);
    CN297_sign_in(23) <= VN1367_sign_out(4);
    CN297_data_in(24) <= VN1502_data_out(4);
    CN297_sign_in(24) <= VN1502_sign_out(4);
    CN297_data_in(25) <= VN1629_data_out(4);
    CN297_sign_in(25) <= VN1629_sign_out(4);
    CN297_data_in(26) <= VN1734_data_out(4);
    CN297_sign_in(26) <= VN1734_sign_out(4);
    CN297_data_in(27) <= VN1744_data_out(4);
    CN297_sign_in(27) <= VN1744_sign_out(4);
    CN297_data_in(28) <= VN1763_data_out(4);
    CN297_sign_in(28) <= VN1763_sign_out(4);
    CN297_data_in(29) <= VN1781_data_out(4);
    CN297_sign_in(29) <= VN1781_sign_out(4);
    CN297_data_in(30) <= VN1784_data_out(4);
    CN297_sign_in(30) <= VN1784_sign_out(4);
    CN297_data_in(31) <= VN1868_data_out(4);
    CN297_sign_in(31) <= VN1868_sign_out(4);
    CN298_data_in(0) <= VN12_data_out(4);
    CN298_sign_in(0) <= VN12_sign_out(4);
    CN298_data_in(1) <= VN91_data_out(4);
    CN298_sign_in(1) <= VN91_sign_out(4);
    CN298_data_in(2) <= VN148_data_out(4);
    CN298_sign_in(2) <= VN148_sign_out(4);
    CN298_data_in(3) <= VN198_data_out(4);
    CN298_sign_in(3) <= VN198_sign_out(4);
    CN298_data_in(4) <= VN262_data_out(4);
    CN298_sign_in(4) <= VN262_sign_out(4);
    CN298_data_in(5) <= VN282_data_out(4);
    CN298_sign_in(5) <= VN282_sign_out(4);
    CN298_data_in(6) <= VN351_data_out(4);
    CN298_sign_in(6) <= VN351_sign_out(4);
    CN298_data_in(7) <= VN408_data_out(4);
    CN298_sign_in(7) <= VN408_sign_out(4);
    CN298_data_in(8) <= VN485_data_out(4);
    CN298_sign_in(8) <= VN485_sign_out(4);
    CN298_data_in(9) <= VN523_data_out(4);
    CN298_sign_in(9) <= VN523_sign_out(4);
    CN298_data_in(10) <= VN611_data_out(4);
    CN298_sign_in(10) <= VN611_sign_out(4);
    CN298_data_in(11) <= VN639_data_out(4);
    CN298_sign_in(11) <= VN639_sign_out(4);
    CN298_data_in(12) <= VN704_data_out(4);
    CN298_sign_in(12) <= VN704_sign_out(4);
    CN298_data_in(13) <= VN776_data_out(4);
    CN298_sign_in(13) <= VN776_sign_out(4);
    CN298_data_in(14) <= VN800_data_out(4);
    CN298_sign_in(14) <= VN800_sign_out(4);
    CN298_data_in(15) <= VN849_data_out(4);
    CN298_sign_in(15) <= VN849_sign_out(4);
    CN298_data_in(16) <= VN942_data_out(4);
    CN298_sign_in(16) <= VN942_sign_out(4);
    CN298_data_in(17) <= VN953_data_out(4);
    CN298_sign_in(17) <= VN953_sign_out(4);
    CN298_data_in(18) <= VN1020_data_out(4);
    CN298_sign_in(18) <= VN1020_sign_out(4);
    CN298_data_in(19) <= VN1129_data_out(4);
    CN298_sign_in(19) <= VN1129_sign_out(4);
    CN298_data_in(20) <= VN1194_data_out(4);
    CN298_sign_in(20) <= VN1194_sign_out(4);
    CN298_data_in(21) <= VN1224_data_out(4);
    CN298_sign_in(21) <= VN1224_sign_out(4);
    CN298_data_in(22) <= VN1234_data_out(4);
    CN298_sign_in(22) <= VN1234_sign_out(4);
    CN298_data_in(23) <= VN1323_data_out(4);
    CN298_sign_in(23) <= VN1323_sign_out(4);
    CN298_data_in(24) <= VN1495_data_out(4);
    CN298_sign_in(24) <= VN1495_sign_out(4);
    CN298_data_in(25) <= VN1508_data_out(4);
    CN298_sign_in(25) <= VN1508_sign_out(4);
    CN298_data_in(26) <= VN1572_data_out(4);
    CN298_sign_in(26) <= VN1572_sign_out(4);
    CN298_data_in(27) <= VN1602_data_out(4);
    CN298_sign_in(27) <= VN1602_sign_out(4);
    CN298_data_in(28) <= VN1639_data_out(4);
    CN298_sign_in(28) <= VN1639_sign_out(4);
    CN298_data_in(29) <= VN1772_data_out(4);
    CN298_sign_in(29) <= VN1772_sign_out(4);
    CN298_data_in(30) <= VN1776_data_out(4);
    CN298_sign_in(30) <= VN1776_sign_out(4);
    CN298_data_in(31) <= VN1869_data_out(4);
    CN298_sign_in(31) <= VN1869_sign_out(4);
    CN299_data_in(0) <= VN83_data_out(4);
    CN299_sign_in(0) <= VN83_sign_out(4);
    CN299_data_in(1) <= VN130_data_out(4);
    CN299_sign_in(1) <= VN130_sign_out(4);
    CN299_data_in(2) <= VN176_data_out(4);
    CN299_sign_in(2) <= VN176_sign_out(4);
    CN299_data_in(3) <= VN264_data_out(4);
    CN299_sign_in(3) <= VN264_sign_out(4);
    CN299_data_in(4) <= VN314_data_out(4);
    CN299_sign_in(4) <= VN314_sign_out(4);
    CN299_data_in(5) <= VN385_data_out(4);
    CN299_sign_in(5) <= VN385_sign_out(4);
    CN299_data_in(6) <= VN393_data_out(4);
    CN299_sign_in(6) <= VN393_sign_out(4);
    CN299_data_in(7) <= VN462_data_out(4);
    CN299_sign_in(7) <= VN462_sign_out(4);
    CN299_data_in(8) <= VN527_data_out(4);
    CN299_sign_in(8) <= VN527_sign_out(4);
    CN299_data_in(9) <= VN637_data_out(4);
    CN299_sign_in(9) <= VN637_sign_out(4);
    CN299_data_in(10) <= VN767_data_out(4);
    CN299_sign_in(10) <= VN767_sign_out(4);
    CN299_data_in(11) <= VN808_data_out(4);
    CN299_sign_in(11) <= VN808_sign_out(4);
    CN299_data_in(12) <= VN885_data_out(4);
    CN299_sign_in(12) <= VN885_sign_out(4);
    CN299_data_in(13) <= VN936_data_out(4);
    CN299_sign_in(13) <= VN936_sign_out(4);
    CN299_data_in(14) <= VN967_data_out(4);
    CN299_sign_in(14) <= VN967_sign_out(4);
    CN299_data_in(15) <= VN1040_data_out(4);
    CN299_sign_in(15) <= VN1040_sign_out(4);
    CN299_data_in(16) <= VN1079_data_out(4);
    CN299_sign_in(16) <= VN1079_sign_out(4);
    CN299_data_in(17) <= VN1146_data_out(4);
    CN299_sign_in(17) <= VN1146_sign_out(4);
    CN299_data_in(18) <= VN1201_data_out(4);
    CN299_sign_in(18) <= VN1201_sign_out(4);
    CN299_data_in(19) <= VN1271_data_out(4);
    CN299_sign_in(19) <= VN1271_sign_out(4);
    CN299_data_in(20) <= VN1382_data_out(4);
    CN299_sign_in(20) <= VN1382_sign_out(4);
    CN299_data_in(21) <= VN1451_data_out(4);
    CN299_sign_in(21) <= VN1451_sign_out(4);
    CN299_data_in(22) <= VN1467_data_out(4);
    CN299_sign_in(22) <= VN1467_sign_out(4);
    CN299_data_in(23) <= VN1477_data_out(4);
    CN299_sign_in(23) <= VN1477_sign_out(4);
    CN299_data_in(24) <= VN1498_data_out(4);
    CN299_sign_in(24) <= VN1498_sign_out(4);
    CN299_data_in(25) <= VN1538_data_out(4);
    CN299_sign_in(25) <= VN1538_sign_out(4);
    CN299_data_in(26) <= VN1647_data_out(4);
    CN299_sign_in(26) <= VN1647_sign_out(4);
    CN299_data_in(27) <= VN1733_data_out(4);
    CN299_sign_in(27) <= VN1733_sign_out(4);
    CN299_data_in(28) <= VN1746_data_out(4);
    CN299_sign_in(28) <= VN1746_sign_out(4);
    CN299_data_in(29) <= VN1883_data_out(4);
    CN299_sign_in(29) <= VN1883_sign_out(4);
    CN299_data_in(30) <= VN1889_data_out(4);
    CN299_sign_in(30) <= VN1889_sign_out(4);
    CN299_data_in(31) <= VN1912_data_out(4);
    CN299_sign_in(31) <= VN1912_sign_out(4);
    CN300_data_in(0) <= VN11_data_out(4);
    CN300_sign_in(0) <= VN11_sign_out(4);
    CN300_data_in(1) <= VN99_data_out(4);
    CN300_sign_in(1) <= VN99_sign_out(4);
    CN300_data_in(2) <= VN143_data_out(4);
    CN300_sign_in(2) <= VN143_sign_out(4);
    CN300_data_in(3) <= VN195_data_out(4);
    CN300_sign_in(3) <= VN195_sign_out(4);
    CN300_data_in(4) <= VN299_data_out(4);
    CN300_sign_in(4) <= VN299_sign_out(4);
    CN300_data_in(5) <= VN335_data_out(4);
    CN300_sign_in(5) <= VN335_sign_out(4);
    CN300_data_in(6) <= VN419_data_out(4);
    CN300_sign_in(6) <= VN419_sign_out(4);
    CN300_data_in(7) <= VN459_data_out(4);
    CN300_sign_in(7) <= VN459_sign_out(4);
    CN300_data_in(8) <= VN591_data_out(4);
    CN300_sign_in(8) <= VN591_sign_out(4);
    CN300_data_in(9) <= VN618_data_out(4);
    CN300_sign_in(9) <= VN618_sign_out(4);
    CN300_data_in(10) <= VN703_data_out(4);
    CN300_sign_in(10) <= VN703_sign_out(4);
    CN300_data_in(11) <= VN735_data_out(4);
    CN300_sign_in(11) <= VN735_sign_out(4);
    CN300_data_in(12) <= VN804_data_out(4);
    CN300_sign_in(12) <= VN804_sign_out(4);
    CN300_data_in(13) <= VN841_data_out(4);
    CN300_sign_in(13) <= VN841_sign_out(4);
    CN300_data_in(14) <= VN920_data_out(4);
    CN300_sign_in(14) <= VN920_sign_out(4);
    CN300_data_in(15) <= VN1041_data_out(4);
    CN300_sign_in(15) <= VN1041_sign_out(4);
    CN300_data_in(16) <= VN1087_data_out(4);
    CN300_sign_in(16) <= VN1087_sign_out(4);
    CN300_data_in(17) <= VN1151_data_out(4);
    CN300_sign_in(17) <= VN1151_sign_out(4);
    CN300_data_in(18) <= VN1326_data_out(4);
    CN300_sign_in(18) <= VN1326_sign_out(4);
    CN300_data_in(19) <= VN1348_data_out(4);
    CN300_sign_in(19) <= VN1348_sign_out(4);
    CN300_data_in(20) <= VN1426_data_out(4);
    CN300_sign_in(20) <= VN1426_sign_out(4);
    CN300_data_in(21) <= VN1497_data_out(4);
    CN300_sign_in(21) <= VN1497_sign_out(4);
    CN300_data_in(22) <= VN1518_data_out(4);
    CN300_sign_in(22) <= VN1518_sign_out(4);
    CN300_data_in(23) <= VN1522_data_out(4);
    CN300_sign_in(23) <= VN1522_sign_out(4);
    CN300_data_in(24) <= VN1557_data_out(4);
    CN300_sign_in(24) <= VN1557_sign_out(4);
    CN300_data_in(25) <= VN1587_data_out(4);
    CN300_sign_in(25) <= VN1587_sign_out(4);
    CN300_data_in(26) <= VN1625_data_out(4);
    CN300_sign_in(26) <= VN1625_sign_out(4);
    CN300_data_in(27) <= VN1680_data_out(4);
    CN300_sign_in(27) <= VN1680_sign_out(4);
    CN300_data_in(28) <= VN1774_data_out(4);
    CN300_sign_in(28) <= VN1774_sign_out(4);
    CN300_data_in(29) <= VN1831_data_out(4);
    CN300_sign_in(29) <= VN1831_sign_out(4);
    CN300_data_in(30) <= VN1859_data_out(4);
    CN300_sign_in(30) <= VN1859_sign_out(4);
    CN300_data_in(31) <= VN1894_data_out(4);
    CN300_sign_in(31) <= VN1894_sign_out(4);
    CN301_data_in(0) <= VN10_data_out(4);
    CN301_sign_in(0) <= VN10_sign_out(4);
    CN301_data_in(1) <= VN103_data_out(4);
    CN301_sign_in(1) <= VN103_sign_out(4);
    CN301_data_in(2) <= VN154_data_out(4);
    CN301_sign_in(2) <= VN154_sign_out(4);
    CN301_data_in(3) <= VN220_data_out(4);
    CN301_sign_in(3) <= VN220_sign_out(4);
    CN301_data_in(4) <= VN270_data_out(4);
    CN301_sign_in(4) <= VN270_sign_out(4);
    CN301_data_in(5) <= VN309_data_out(4);
    CN301_sign_in(5) <= VN309_sign_out(4);
    CN301_data_in(6) <= VN389_data_out(4);
    CN301_sign_in(6) <= VN389_sign_out(4);
    CN301_data_in(7) <= VN409_data_out(4);
    CN301_sign_in(7) <= VN409_sign_out(4);
    CN301_data_in(8) <= VN474_data_out(4);
    CN301_sign_in(8) <= VN474_sign_out(4);
    CN301_data_in(9) <= VN526_data_out(4);
    CN301_sign_in(9) <= VN526_sign_out(4);
    CN301_data_in(10) <= VN697_data_out(4);
    CN301_sign_in(10) <= VN697_sign_out(4);
    CN301_data_in(11) <= VN741_data_out(4);
    CN301_sign_in(11) <= VN741_sign_out(4);
    CN301_data_in(12) <= VN809_data_out(4);
    CN301_sign_in(12) <= VN809_sign_out(4);
    CN301_data_in(13) <= VN850_data_out(4);
    CN301_sign_in(13) <= VN850_sign_out(4);
    CN301_data_in(14) <= VN983_data_out(4);
    CN301_sign_in(14) <= VN983_sign_out(4);
    CN301_data_in(15) <= VN1019_data_out(4);
    CN301_sign_in(15) <= VN1019_sign_out(4);
    CN301_data_in(16) <= VN1082_data_out(4);
    CN301_sign_in(16) <= VN1082_sign_out(4);
    CN301_data_in(17) <= VN1243_data_out(4);
    CN301_sign_in(17) <= VN1243_sign_out(4);
    CN301_data_in(18) <= VN1349_data_out(4);
    CN301_sign_in(18) <= VN1349_sign_out(4);
    CN301_data_in(19) <= VN1428_data_out(4);
    CN301_sign_in(19) <= VN1428_sign_out(4);
    CN301_data_in(20) <= VN1514_data_out(4);
    CN301_sign_in(20) <= VN1514_sign_out(4);
    CN301_data_in(21) <= VN1553_data_out(4);
    CN301_sign_in(21) <= VN1553_sign_out(4);
    CN301_data_in(22) <= VN1691_data_out(4);
    CN301_sign_in(22) <= VN1691_sign_out(4);
    CN301_data_in(23) <= VN1773_data_out(4);
    CN301_sign_in(23) <= VN1773_sign_out(4);
    CN301_data_in(24) <= VN1812_data_out(4);
    CN301_sign_in(24) <= VN1812_sign_out(4);
    CN301_data_in(25) <= VN1847_data_out(4);
    CN301_sign_in(25) <= VN1847_sign_out(4);
    CN301_data_in(26) <= VN1855_data_out(4);
    CN301_sign_in(26) <= VN1855_sign_out(4);
    CN301_data_in(27) <= VN1856_data_out(4);
    CN301_sign_in(27) <= VN1856_sign_out(4);
    CN301_data_in(28) <= VN1903_data_out(4);
    CN301_sign_in(28) <= VN1903_sign_out(4);
    CN301_data_in(29) <= VN1904_data_out(4);
    CN301_sign_in(29) <= VN1904_sign_out(4);
    CN301_data_in(30) <= VN1916_data_out(4);
    CN301_sign_in(30) <= VN1916_sign_out(4);
    CN301_data_in(31) <= VN1920_data_out(4);
    CN301_sign_in(31) <= VN1920_sign_out(4);
    CN302_data_in(0) <= VN9_data_out(4);
    CN302_sign_in(0) <= VN9_sign_out(4);
    CN302_data_in(1) <= VN110_data_out(4);
    CN302_sign_in(1) <= VN110_sign_out(4);
    CN302_data_in(2) <= VN124_data_out(4);
    CN302_sign_in(2) <= VN124_sign_out(4);
    CN302_data_in(3) <= VN206_data_out(4);
    CN302_sign_in(3) <= VN206_sign_out(4);
    CN302_data_in(4) <= VN227_data_out(4);
    CN302_sign_in(4) <= VN227_sign_out(4);
    CN302_data_in(5) <= VN321_data_out(4);
    CN302_sign_in(5) <= VN321_sign_out(4);
    CN302_data_in(6) <= VN398_data_out(4);
    CN302_sign_in(6) <= VN398_sign_out(4);
    CN302_data_in(7) <= VN521_data_out(4);
    CN302_sign_in(7) <= VN521_sign_out(4);
    CN302_data_in(8) <= VN583_data_out(4);
    CN302_sign_in(8) <= VN583_sign_out(4);
    CN302_data_in(9) <= VN679_data_out(4);
    CN302_sign_in(9) <= VN679_sign_out(4);
    CN302_data_in(10) <= VN725_data_out(4);
    CN302_sign_in(10) <= VN725_sign_out(4);
    CN302_data_in(11) <= VN877_data_out(4);
    CN302_sign_in(11) <= VN877_sign_out(4);
    CN302_data_in(12) <= VN892_data_out(4);
    CN302_sign_in(12) <= VN892_sign_out(4);
    CN302_data_in(13) <= VN946_data_out(4);
    CN302_sign_in(13) <= VN946_sign_out(4);
    CN302_data_in(14) <= VN1011_data_out(4);
    CN302_sign_in(14) <= VN1011_sign_out(4);
    CN302_data_in(15) <= VN1150_data_out(4);
    CN302_sign_in(15) <= VN1150_sign_out(4);
    CN302_data_in(16) <= VN1199_data_out(4);
    CN302_sign_in(16) <= VN1199_sign_out(4);
    CN302_data_in(17) <= VN1381_data_out(4);
    CN302_sign_in(17) <= VN1381_sign_out(4);
    CN302_data_in(18) <= VN1412_data_out(4);
    CN302_sign_in(18) <= VN1412_sign_out(4);
    CN302_data_in(19) <= VN1443_data_out(4);
    CN302_sign_in(19) <= VN1443_sign_out(4);
    CN302_data_in(20) <= VN1573_data_out(4);
    CN302_sign_in(20) <= VN1573_sign_out(4);
    CN302_data_in(21) <= VN1590_data_out(4);
    CN302_sign_in(21) <= VN1590_sign_out(4);
    CN302_data_in(22) <= VN1649_data_out(4);
    CN302_sign_in(22) <= VN1649_sign_out(4);
    CN302_data_in(23) <= VN1759_data_out(4);
    CN302_sign_in(23) <= VN1759_sign_out(4);
    CN302_data_in(24) <= VN1769_data_out(4);
    CN302_sign_in(24) <= VN1769_sign_out(4);
    CN302_data_in(25) <= VN1816_data_out(4);
    CN302_sign_in(25) <= VN1816_sign_out(4);
    CN302_data_in(26) <= VN1818_data_out(4);
    CN302_sign_in(26) <= VN1818_sign_out(4);
    CN302_data_in(27) <= VN1821_data_out(4);
    CN302_sign_in(27) <= VN1821_sign_out(4);
    CN302_data_in(28) <= VN1823_data_out(4);
    CN302_sign_in(28) <= VN1823_sign_out(4);
    CN302_data_in(29) <= VN1885_data_out(4);
    CN302_sign_in(29) <= VN1885_sign_out(4);
    CN302_data_in(30) <= VN1914_data_out(4);
    CN302_sign_in(30) <= VN1914_sign_out(4);
    CN302_data_in(31) <= VN1917_data_out(4);
    CN302_sign_in(31) <= VN1917_sign_out(4);
    CN303_data_in(0) <= VN8_data_out(4);
    CN303_sign_in(0) <= VN8_sign_out(4);
    CN303_data_in(1) <= VN102_data_out(4);
    CN303_sign_in(1) <= VN102_sign_out(4);
    CN303_data_in(2) <= VN112_data_out(4);
    CN303_sign_in(2) <= VN112_sign_out(4);
    CN303_data_in(3) <= VN178_data_out(4);
    CN303_sign_in(3) <= VN178_sign_out(4);
    CN303_data_in(4) <= VN235_data_out(4);
    CN303_sign_in(4) <= VN235_sign_out(4);
    CN303_data_in(5) <= VN293_data_out(4);
    CN303_sign_in(5) <= VN293_sign_out(4);
    CN303_data_in(6) <= VN382_data_out(4);
    CN303_sign_in(6) <= VN382_sign_out(4);
    CN303_data_in(7) <= VN415_data_out(4);
    CN303_sign_in(7) <= VN415_sign_out(4);
    CN303_data_in(8) <= VN497_data_out(4);
    CN303_sign_in(8) <= VN497_sign_out(4);
    CN303_data_in(9) <= VN506_data_out(4);
    CN303_sign_in(9) <= VN506_sign_out(4);
    CN303_data_in(10) <= VN581_data_out(4);
    CN303_sign_in(10) <= VN581_sign_out(4);
    CN303_data_in(11) <= VN640_data_out(4);
    CN303_sign_in(11) <= VN640_sign_out(4);
    CN303_data_in(12) <= VN686_data_out(4);
    CN303_sign_in(12) <= VN686_sign_out(4);
    CN303_data_in(13) <= VN727_data_out(4);
    CN303_sign_in(13) <= VN727_sign_out(4);
    CN303_data_in(14) <= VN823_data_out(4);
    CN303_sign_in(14) <= VN823_sign_out(4);
    CN303_data_in(15) <= VN836_data_out(4);
    CN303_sign_in(15) <= VN836_sign_out(4);
    CN303_data_in(16) <= VN890_data_out(4);
    CN303_sign_in(16) <= VN890_sign_out(4);
    CN303_data_in(17) <= VN947_data_out(4);
    CN303_sign_in(17) <= VN947_sign_out(4);
    CN303_data_in(18) <= VN1003_data_out(4);
    CN303_sign_in(18) <= VN1003_sign_out(4);
    CN303_data_in(19) <= VN1027_data_out(4);
    CN303_sign_in(19) <= VN1027_sign_out(4);
    CN303_data_in(20) <= VN1078_data_out(4);
    CN303_sign_in(20) <= VN1078_sign_out(4);
    CN303_data_in(21) <= VN1144_data_out(4);
    CN303_sign_in(21) <= VN1144_sign_out(4);
    CN303_data_in(22) <= VN1181_data_out(4);
    CN303_sign_in(22) <= VN1181_sign_out(4);
    CN303_data_in(23) <= VN1373_data_out(4);
    CN303_sign_in(23) <= VN1373_sign_out(4);
    CN303_data_in(24) <= VN1468_data_out(4);
    CN303_sign_in(24) <= VN1468_sign_out(4);
    CN303_data_in(25) <= VN1520_data_out(4);
    CN303_sign_in(25) <= VN1520_sign_out(4);
    CN303_data_in(26) <= VN1546_data_out(4);
    CN303_sign_in(26) <= VN1546_sign_out(4);
    CN303_data_in(27) <= VN1592_data_out(4);
    CN303_sign_in(27) <= VN1592_sign_out(4);
    CN303_data_in(28) <= VN1642_data_out(4);
    CN303_sign_in(28) <= VN1642_sign_out(4);
    CN303_data_in(29) <= VN1681_data_out(4);
    CN303_sign_in(29) <= VN1681_sign_out(4);
    CN303_data_in(30) <= VN1762_data_out(4);
    CN303_sign_in(30) <= VN1762_sign_out(4);
    CN303_data_in(31) <= VN1870_data_out(4);
    CN303_sign_in(31) <= VN1870_sign_out(4);
    CN304_data_in(0) <= VN7_data_out(4);
    CN304_sign_in(0) <= VN7_sign_out(4);
    CN304_data_in(1) <= VN97_data_out(4);
    CN304_sign_in(1) <= VN97_sign_out(4);
    CN304_data_in(2) <= VN157_data_out(4);
    CN304_sign_in(2) <= VN157_sign_out(4);
    CN304_data_in(3) <= VN222_data_out(4);
    CN304_sign_in(3) <= VN222_sign_out(4);
    CN304_data_in(4) <= VN263_data_out(4);
    CN304_sign_in(4) <= VN263_sign_out(4);
    CN304_data_in(5) <= VN283_data_out(4);
    CN304_sign_in(5) <= VN283_sign_out(4);
    CN304_data_in(6) <= VN359_data_out(4);
    CN304_sign_in(6) <= VN359_sign_out(4);
    CN304_data_in(7) <= VN446_data_out(4);
    CN304_sign_in(7) <= VN446_sign_out(4);
    CN304_data_in(8) <= VN451_data_out(4);
    CN304_sign_in(8) <= VN451_sign_out(4);
    CN304_data_in(9) <= VN512_data_out(4);
    CN304_sign_in(9) <= VN512_sign_out(4);
    CN304_data_in(10) <= VN595_data_out(4);
    CN304_sign_in(10) <= VN595_sign_out(4);
    CN304_data_in(11) <= VN619_data_out(4);
    CN304_sign_in(11) <= VN619_sign_out(4);
    CN304_data_in(12) <= VN709_data_out(4);
    CN304_sign_in(12) <= VN709_sign_out(4);
    CN304_data_in(13) <= VN751_data_out(4);
    CN304_sign_in(13) <= VN751_sign_out(4);
    CN304_data_in(14) <= VN828_data_out(4);
    CN304_sign_in(14) <= VN828_sign_out(4);
    CN304_data_in(15) <= VN865_data_out(4);
    CN304_sign_in(15) <= VN865_sign_out(4);
    CN304_data_in(16) <= VN925_data_out(4);
    CN304_sign_in(16) <= VN925_sign_out(4);
    CN304_data_in(17) <= VN982_data_out(4);
    CN304_sign_in(17) <= VN982_sign_out(4);
    CN304_data_in(18) <= VN1031_data_out(4);
    CN304_sign_in(18) <= VN1031_sign_out(4);
    CN304_data_in(19) <= VN1098_data_out(4);
    CN304_sign_in(19) <= VN1098_sign_out(4);
    CN304_data_in(20) <= VN1126_data_out(4);
    CN304_sign_in(20) <= VN1126_sign_out(4);
    CN304_data_in(21) <= VN1167_data_out(4);
    CN304_sign_in(21) <= VN1167_sign_out(4);
    CN304_data_in(22) <= VN1184_data_out(4);
    CN304_sign_in(22) <= VN1184_sign_out(4);
    CN304_data_in(23) <= VN1256_data_out(4);
    CN304_sign_in(23) <= VN1256_sign_out(4);
    CN304_data_in(24) <= VN1301_data_out(4);
    CN304_sign_in(24) <= VN1301_sign_out(4);
    CN304_data_in(25) <= VN1423_data_out(4);
    CN304_sign_in(25) <= VN1423_sign_out(4);
    CN304_data_in(26) <= VN1571_data_out(4);
    CN304_sign_in(26) <= VN1571_sign_out(4);
    CN304_data_in(27) <= VN1586_data_out(4);
    CN304_sign_in(27) <= VN1586_sign_out(4);
    CN304_data_in(28) <= VN1613_data_out(4);
    CN304_sign_in(28) <= VN1613_sign_out(4);
    CN304_data_in(29) <= VN1716_data_out(4);
    CN304_sign_in(29) <= VN1716_sign_out(4);
    CN304_data_in(30) <= VN1809_data_out(4);
    CN304_sign_in(30) <= VN1809_sign_out(4);
    CN304_data_in(31) <= VN1871_data_out(4);
    CN304_sign_in(31) <= VN1871_sign_out(4);
    CN305_data_in(0) <= VN6_data_out(4);
    CN305_sign_in(0) <= VN6_sign_out(4);
    CN305_data_in(1) <= VN80_data_out(4);
    CN305_sign_in(1) <= VN80_sign_out(4);
    CN305_data_in(2) <= VN115_data_out(4);
    CN305_sign_in(2) <= VN115_sign_out(4);
    CN305_data_in(3) <= VN209_data_out(4);
    CN305_sign_in(3) <= VN209_sign_out(4);
    CN305_data_in(4) <= VN276_data_out(4);
    CN305_sign_in(4) <= VN276_sign_out(4);
    CN305_data_in(5) <= VN323_data_out(4);
    CN305_sign_in(5) <= VN323_sign_out(4);
    CN305_data_in(6) <= VN342_data_out(4);
    CN305_sign_in(6) <= VN342_sign_out(4);
    CN305_data_in(7) <= VN443_data_out(4);
    CN305_sign_in(7) <= VN443_sign_out(4);
    CN305_data_in(8) <= VN501_data_out(4);
    CN305_sign_in(8) <= VN501_sign_out(4);
    CN305_data_in(9) <= VN533_data_out(4);
    CN305_sign_in(9) <= VN533_sign_out(4);
    CN305_data_in(10) <= VN588_data_out(4);
    CN305_sign_in(10) <= VN588_sign_out(4);
    CN305_data_in(11) <= VN636_data_out(4);
    CN305_sign_in(11) <= VN636_sign_out(4);
    CN305_data_in(12) <= VN707_data_out(4);
    CN305_sign_in(12) <= VN707_sign_out(4);
    CN305_data_in(13) <= VN733_data_out(4);
    CN305_sign_in(13) <= VN733_sign_out(4);
    CN305_data_in(14) <= VN813_data_out(4);
    CN305_sign_in(14) <= VN813_sign_out(4);
    CN305_data_in(15) <= VN844_data_out(4);
    CN305_sign_in(15) <= VN844_sign_out(4);
    CN305_data_in(16) <= VN906_data_out(4);
    CN305_sign_in(16) <= VN906_sign_out(4);
    CN305_data_in(17) <= VN974_data_out(4);
    CN305_sign_in(17) <= VN974_sign_out(4);
    CN305_data_in(18) <= VN1104_data_out(4);
    CN305_sign_in(18) <= VN1104_sign_out(4);
    CN305_data_in(19) <= VN1112_data_out(4);
    CN305_sign_in(19) <= VN1112_sign_out(4);
    CN305_data_in(20) <= VN1133_data_out(4);
    CN305_sign_in(20) <= VN1133_sign_out(4);
    CN305_data_in(21) <= VN1170_data_out(4);
    CN305_sign_in(21) <= VN1170_sign_out(4);
    CN305_data_in(22) <= VN1258_data_out(4);
    CN305_sign_in(22) <= VN1258_sign_out(4);
    CN305_data_in(23) <= VN1292_data_out(4);
    CN305_sign_in(23) <= VN1292_sign_out(4);
    CN305_data_in(24) <= VN1338_data_out(4);
    CN305_sign_in(24) <= VN1338_sign_out(4);
    CN305_data_in(25) <= VN1436_data_out(4);
    CN305_sign_in(25) <= VN1436_sign_out(4);
    CN305_data_in(26) <= VN1505_data_out(4);
    CN305_sign_in(26) <= VN1505_sign_out(4);
    CN305_data_in(27) <= VN1604_data_out(4);
    CN305_sign_in(27) <= VN1604_sign_out(4);
    CN305_data_in(28) <= VN1626_data_out(4);
    CN305_sign_in(28) <= VN1626_sign_out(4);
    CN305_data_in(29) <= VN1685_data_out(4);
    CN305_sign_in(29) <= VN1685_sign_out(4);
    CN305_data_in(30) <= VN1702_data_out(4);
    CN305_sign_in(30) <= VN1702_sign_out(4);
    CN305_data_in(31) <= VN1798_data_out(4);
    CN305_sign_in(31) <= VN1798_sign_out(4);
    CN306_data_in(0) <= VN5_data_out(4);
    CN306_sign_in(0) <= VN5_sign_out(4);
    CN306_data_in(1) <= VN87_data_out(4);
    CN306_sign_in(1) <= VN87_sign_out(4);
    CN306_data_in(2) <= VN136_data_out(4);
    CN306_sign_in(2) <= VN136_sign_out(4);
    CN306_data_in(3) <= VN174_data_out(4);
    CN306_sign_in(3) <= VN174_sign_out(4);
    CN306_data_in(4) <= VN402_data_out(4);
    CN306_sign_in(4) <= VN402_sign_out(4);
    CN306_data_in(5) <= VN448_data_out(4);
    CN306_sign_in(5) <= VN448_sign_out(4);
    CN306_data_in(6) <= VN531_data_out(4);
    CN306_sign_in(6) <= VN531_sign_out(4);
    CN306_data_in(7) <= VN564_data_out(4);
    CN306_sign_in(7) <= VN564_sign_out(4);
    CN306_data_in(8) <= VN663_data_out(4);
    CN306_sign_in(8) <= VN663_sign_out(4);
    CN306_data_in(9) <= VN684_data_out(4);
    CN306_sign_in(9) <= VN684_sign_out(4);
    CN306_data_in(10) <= VN815_data_out(4);
    CN306_sign_in(10) <= VN815_sign_out(4);
    CN306_data_in(11) <= VN909_data_out(4);
    CN306_sign_in(11) <= VN909_sign_out(4);
    CN306_data_in(12) <= VN1030_data_out(4);
    CN306_sign_in(12) <= VN1030_sign_out(4);
    CN306_data_in(13) <= VN1156_data_out(4);
    CN306_sign_in(13) <= VN1156_sign_out(4);
    CN306_data_in(14) <= VN1200_data_out(4);
    CN306_sign_in(14) <= VN1200_sign_out(4);
    CN306_data_in(15) <= VN1244_data_out(4);
    CN306_sign_in(15) <= VN1244_sign_out(4);
    CN306_data_in(16) <= VN1312_data_out(4);
    CN306_sign_in(16) <= VN1312_sign_out(4);
    CN306_data_in(17) <= VN1387_data_out(4);
    CN306_sign_in(17) <= VN1387_sign_out(4);
    CN306_data_in(18) <= VN1462_data_out(4);
    CN306_sign_in(18) <= VN1462_sign_out(4);
    CN306_data_in(19) <= VN1536_data_out(4);
    CN306_sign_in(19) <= VN1536_sign_out(4);
    CN306_data_in(20) <= VN1623_data_out(4);
    CN306_sign_in(20) <= VN1623_sign_out(4);
    CN306_data_in(21) <= VN1667_data_out(4);
    CN306_sign_in(21) <= VN1667_sign_out(4);
    CN306_data_in(22) <= VN1732_data_out(4);
    CN306_sign_in(22) <= VN1732_sign_out(4);
    CN306_data_in(23) <= VN1861_data_out(4);
    CN306_sign_in(23) <= VN1861_sign_out(4);
    CN306_data_in(24) <= VN1876_data_out(4);
    CN306_sign_in(24) <= VN1876_sign_out(4);
    CN306_data_in(25) <= VN1878_data_out(4);
    CN306_sign_in(25) <= VN1878_sign_out(4);
    CN306_data_in(26) <= VN1887_data_out(4);
    CN306_sign_in(26) <= VN1887_sign_out(4);
    CN306_data_in(27) <= VN1890_data_out(4);
    CN306_sign_in(27) <= VN1890_sign_out(4);
    CN306_data_in(28) <= VN1942_data_out(4);
    CN306_sign_in(28) <= VN1942_sign_out(4);
    CN306_data_in(29) <= VN1944_data_out(4);
    CN306_sign_in(29) <= VN1944_sign_out(4);
    CN306_data_in(30) <= VN2016_data_out(4);
    CN306_sign_in(30) <= VN2016_sign_out(4);
    CN306_data_in(31) <= VN2026_data_out(4);
    CN306_sign_in(31) <= VN2026_sign_out(4);
    CN307_data_in(0) <= VN4_data_out(4);
    CN307_sign_in(0) <= VN4_sign_out(4);
    CN307_data_in(1) <= VN107_data_out(4);
    CN307_sign_in(1) <= VN107_sign_out(4);
    CN307_data_in(2) <= VN145_data_out(4);
    CN307_sign_in(2) <= VN145_sign_out(4);
    CN307_data_in(3) <= VN202_data_out(4);
    CN307_sign_in(3) <= VN202_sign_out(4);
    CN307_data_in(4) <= VN230_data_out(4);
    CN307_sign_in(4) <= VN230_sign_out(4);
    CN307_data_in(5) <= VN302_data_out(4);
    CN307_sign_in(5) <= VN302_sign_out(4);
    CN307_data_in(6) <= VN366_data_out(4);
    CN307_sign_in(6) <= VN366_sign_out(4);
    CN307_data_in(7) <= VN395_data_out(4);
    CN307_sign_in(7) <= VN395_sign_out(4);
    CN307_data_in(8) <= VN494_data_out(4);
    CN307_sign_in(8) <= VN494_sign_out(4);
    CN307_data_in(9) <= VN510_data_out(4);
    CN307_sign_in(9) <= VN510_sign_out(4);
    CN307_data_in(10) <= VN574_data_out(4);
    CN307_sign_in(10) <= VN574_sign_out(4);
    CN307_data_in(11) <= VN649_data_out(4);
    CN307_sign_in(11) <= VN649_sign_out(4);
    CN307_data_in(12) <= VN719_data_out(4);
    CN307_sign_in(12) <= VN719_sign_out(4);
    CN307_data_in(13) <= VN752_data_out(4);
    CN307_sign_in(13) <= VN752_sign_out(4);
    CN307_data_in(14) <= VN785_data_out(4);
    CN307_sign_in(14) <= VN785_sign_out(4);
    CN307_data_in(15) <= VN879_data_out(4);
    CN307_sign_in(15) <= VN879_sign_out(4);
    CN307_data_in(16) <= VN893_data_out(4);
    CN307_sign_in(16) <= VN893_sign_out(4);
    CN307_data_in(17) <= VN996_data_out(4);
    CN307_sign_in(17) <= VN996_sign_out(4);
    CN307_data_in(18) <= VN1025_data_out(4);
    CN307_sign_in(18) <= VN1025_sign_out(4);
    CN307_data_in(19) <= VN1091_data_out(4);
    CN307_sign_in(19) <= VN1091_sign_out(4);
    CN307_data_in(20) <= VN1154_data_out(4);
    CN307_sign_in(20) <= VN1154_sign_out(4);
    CN307_data_in(21) <= VN1318_data_out(4);
    CN307_sign_in(21) <= VN1318_sign_out(4);
    CN307_data_in(22) <= VN1470_data_out(4);
    CN307_sign_in(22) <= VN1470_sign_out(4);
    CN307_data_in(23) <= VN1521_data_out(4);
    CN307_sign_in(23) <= VN1521_sign_out(4);
    CN307_data_in(24) <= VN1537_data_out(4);
    CN307_sign_in(24) <= VN1537_sign_out(4);
    CN307_data_in(25) <= VN1637_data_out(4);
    CN307_sign_in(25) <= VN1637_sign_out(4);
    CN307_data_in(26) <= VN1665_data_out(4);
    CN307_sign_in(26) <= VN1665_sign_out(4);
    CN307_data_in(27) <= VN1745_data_out(4);
    CN307_sign_in(27) <= VN1745_sign_out(4);
    CN307_data_in(28) <= VN1748_data_out(4);
    CN307_sign_in(28) <= VN1748_sign_out(4);
    CN307_data_in(29) <= VN1923_data_out(4);
    CN307_sign_in(29) <= VN1923_sign_out(4);
    CN307_data_in(30) <= VN1932_data_out(4);
    CN307_sign_in(30) <= VN1932_sign_out(4);
    CN307_data_in(31) <= VN1940_data_out(4);
    CN307_sign_in(31) <= VN1940_sign_out(4);
    CN308_data_in(0) <= VN140_data_out(4);
    CN308_sign_in(0) <= VN140_sign_out(4);
    CN308_data_in(1) <= VN199_data_out(4);
    CN308_sign_in(1) <= VN199_sign_out(4);
    CN308_data_in(2) <= VN251_data_out(4);
    CN308_sign_in(2) <= VN251_sign_out(4);
    CN308_data_in(3) <= VN311_data_out(4);
    CN308_sign_in(3) <= VN311_sign_out(4);
    CN308_data_in(4) <= VN336_data_out(4);
    CN308_sign_in(4) <= VN336_sign_out(4);
    CN308_data_in(5) <= VN426_data_out(4);
    CN308_sign_in(5) <= VN426_sign_out(4);
    CN308_data_in(6) <= VN475_data_out(4);
    CN308_sign_in(6) <= VN475_sign_out(4);
    CN308_data_in(7) <= VN547_data_out(4);
    CN308_sign_in(7) <= VN547_sign_out(4);
    CN308_data_in(8) <= VN568_data_out(4);
    CN308_sign_in(8) <= VN568_sign_out(4);
    CN308_data_in(9) <= VN669_data_out(4);
    CN308_sign_in(9) <= VN669_sign_out(4);
    CN308_data_in(10) <= VN726_data_out(4);
    CN308_sign_in(10) <= VN726_sign_out(4);
    CN308_data_in(11) <= VN821_data_out(4);
    CN308_sign_in(11) <= VN821_sign_out(4);
    CN308_data_in(12) <= VN876_data_out(4);
    CN308_sign_in(12) <= VN876_sign_out(4);
    CN308_data_in(13) <= VN926_data_out(4);
    CN308_sign_in(13) <= VN926_sign_out(4);
    CN308_data_in(14) <= VN1008_data_out(4);
    CN308_sign_in(14) <= VN1008_sign_out(4);
    CN308_data_in(15) <= VN1063_data_out(4);
    CN308_sign_in(15) <= VN1063_sign_out(4);
    CN308_data_in(16) <= VN1131_data_out(4);
    CN308_sign_in(16) <= VN1131_sign_out(4);
    CN308_data_in(17) <= VN1241_data_out(4);
    CN308_sign_in(17) <= VN1241_sign_out(4);
    CN308_data_in(18) <= VN1280_data_out(4);
    CN308_sign_in(18) <= VN1280_sign_out(4);
    CN308_data_in(19) <= VN1392_data_out(4);
    CN308_sign_in(19) <= VN1392_sign_out(4);
    CN308_data_in(20) <= VN1438_data_out(4);
    CN308_sign_in(20) <= VN1438_sign_out(4);
    CN308_data_in(21) <= VN1503_data_out(4);
    CN308_sign_in(21) <= VN1503_sign_out(4);
    CN308_data_in(22) <= VN1597_data_out(4);
    CN308_sign_in(22) <= VN1597_sign_out(4);
    CN308_data_in(23) <= VN1674_data_out(4);
    CN308_sign_in(23) <= VN1674_sign_out(4);
    CN308_data_in(24) <= VN1703_data_out(4);
    CN308_sign_in(24) <= VN1703_sign_out(4);
    CN308_data_in(25) <= VN1741_data_out(4);
    CN308_sign_in(25) <= VN1741_sign_out(4);
    CN308_data_in(26) <= VN1930_data_out(4);
    CN308_sign_in(26) <= VN1930_sign_out(4);
    CN308_data_in(27) <= VN1946_data_out(4);
    CN308_sign_in(27) <= VN1946_sign_out(4);
    CN308_data_in(28) <= VN1966_data_out(4);
    CN308_sign_in(28) <= VN1966_sign_out(4);
    CN308_data_in(29) <= VN1979_data_out(4);
    CN308_sign_in(29) <= VN1979_sign_out(4);
    CN308_data_in(30) <= VN2018_data_out(4);
    CN308_sign_in(30) <= VN2018_sign_out(4);
    CN308_data_in(31) <= VN2024_data_out(4);
    CN308_sign_in(31) <= VN2024_sign_out(4);
    CN309_data_in(0) <= VN3_data_out(4);
    CN309_sign_in(0) <= VN3_sign_out(4);
    CN309_data_in(1) <= VN86_data_out(4);
    CN309_sign_in(1) <= VN86_sign_out(4);
    CN309_data_in(2) <= VN146_data_out(4);
    CN309_sign_in(2) <= VN146_sign_out(4);
    CN309_data_in(3) <= VN214_data_out(4);
    CN309_sign_in(3) <= VN214_sign_out(4);
    CN309_data_in(4) <= VN265_data_out(4);
    CN309_sign_in(4) <= VN265_sign_out(4);
    CN309_data_in(5) <= VN307_data_out(4);
    CN309_sign_in(5) <= VN307_sign_out(4);
    CN309_data_in(6) <= VN384_data_out(4);
    CN309_sign_in(6) <= VN384_sign_out(4);
    CN309_data_in(7) <= VN437_data_out(4);
    CN309_sign_in(7) <= VN437_sign_out(4);
    CN309_data_in(8) <= VN458_data_out(4);
    CN309_sign_in(8) <= VN458_sign_out(4);
    CN309_data_in(9) <= VN550_data_out(4);
    CN309_sign_in(9) <= VN550_sign_out(4);
    CN309_data_in(10) <= VN571_data_out(4);
    CN309_sign_in(10) <= VN571_sign_out(4);
    CN309_data_in(11) <= VN664_data_out(4);
    CN309_sign_in(11) <= VN664_sign_out(4);
    CN309_data_in(12) <= VN710_data_out(4);
    CN309_sign_in(12) <= VN710_sign_out(4);
    CN309_data_in(13) <= VN740_data_out(4);
    CN309_sign_in(13) <= VN740_sign_out(4);
    CN309_data_in(14) <= VN779_data_out(4);
    CN309_sign_in(14) <= VN779_sign_out(4);
    CN309_data_in(15) <= VN839_data_out(4);
    CN309_sign_in(15) <= VN839_sign_out(4);
    CN309_data_in(16) <= VN889_data_out(4);
    CN309_sign_in(16) <= VN889_sign_out(4);
    CN309_data_in(17) <= VN995_data_out(4);
    CN309_sign_in(17) <= VN995_sign_out(4);
    CN309_data_in(18) <= VN1015_data_out(4);
    CN309_sign_in(18) <= VN1015_sign_out(4);
    CN309_data_in(19) <= VN1097_data_out(4);
    CN309_sign_in(19) <= VN1097_sign_out(4);
    CN309_data_in(20) <= VN1177_data_out(4);
    CN309_sign_in(20) <= VN1177_sign_out(4);
    CN309_data_in(21) <= VN1268_data_out(4);
    CN309_sign_in(21) <= VN1268_sign_out(4);
    CN309_data_in(22) <= VN1304_data_out(4);
    CN309_sign_in(22) <= VN1304_sign_out(4);
    CN309_data_in(23) <= VN1370_data_out(4);
    CN309_sign_in(23) <= VN1370_sign_out(4);
    CN309_data_in(24) <= VN1420_data_out(4);
    CN309_sign_in(24) <= VN1420_sign_out(4);
    CN309_data_in(25) <= VN1427_data_out(4);
    CN309_sign_in(25) <= VN1427_sign_out(4);
    CN309_data_in(26) <= VN1481_data_out(4);
    CN309_sign_in(26) <= VN1481_sign_out(4);
    CN309_data_in(27) <= VN1513_data_out(4);
    CN309_sign_in(27) <= VN1513_sign_out(4);
    CN309_data_in(28) <= VN1715_data_out(4);
    CN309_sign_in(28) <= VN1715_sign_out(4);
    CN309_data_in(29) <= VN1730_data_out(4);
    CN309_sign_in(29) <= VN1730_sign_out(4);
    CN309_data_in(30) <= VN1742_data_out(4);
    CN309_sign_in(30) <= VN1742_sign_out(4);
    CN309_data_in(31) <= VN1872_data_out(4);
    CN309_sign_in(31) <= VN1872_sign_out(4);
    CN310_data_in(0) <= VN2_data_out(4);
    CN310_sign_in(0) <= VN2_sign_out(4);
    CN310_data_in(1) <= VN65_data_out(4);
    CN310_sign_in(1) <= VN65_sign_out(4);
    CN310_data_in(2) <= VN135_data_out(4);
    CN310_sign_in(2) <= VN135_sign_out(4);
    CN310_data_in(3) <= VN261_data_out(4);
    CN310_sign_in(3) <= VN261_sign_out(4);
    CN310_data_in(4) <= VN312_data_out(4);
    CN310_sign_in(4) <= VN312_sign_out(4);
    CN310_data_in(5) <= VN369_data_out(4);
    CN310_sign_in(5) <= VN369_sign_out(4);
    CN310_data_in(6) <= VN430_data_out(4);
    CN310_sign_in(6) <= VN430_sign_out(4);
    CN310_data_in(7) <= VN470_data_out(4);
    CN310_sign_in(7) <= VN470_sign_out(4);
    CN310_data_in(8) <= VN534_data_out(4);
    CN310_sign_in(8) <= VN534_sign_out(4);
    CN310_data_in(9) <= VN561_data_out(4);
    CN310_sign_in(9) <= VN561_sign_out(4);
    CN310_data_in(10) <= VN653_data_out(4);
    CN310_sign_in(10) <= VN653_sign_out(4);
    CN310_data_in(11) <= VN685_data_out(4);
    CN310_sign_in(11) <= VN685_sign_out(4);
    CN310_data_in(12) <= VN786_data_out(4);
    CN310_sign_in(12) <= VN786_sign_out(4);
    CN310_data_in(13) <= VN861_data_out(4);
    CN310_sign_in(13) <= VN861_sign_out(4);
    CN310_data_in(14) <= VN917_data_out(4);
    CN310_sign_in(14) <= VN917_sign_out(4);
    CN310_data_in(15) <= VN990_data_out(4);
    CN310_sign_in(15) <= VN990_sign_out(4);
    CN310_data_in(16) <= VN1036_data_out(4);
    CN310_sign_in(16) <= VN1036_sign_out(4);
    CN310_data_in(17) <= VN1202_data_out(4);
    CN310_sign_in(17) <= VN1202_sign_out(4);
    CN310_data_in(18) <= VN1219_data_out(4);
    CN310_sign_in(18) <= VN1219_sign_out(4);
    CN310_data_in(19) <= VN1253_data_out(4);
    CN310_sign_in(19) <= VN1253_sign_out(4);
    CN310_data_in(20) <= VN1417_data_out(4);
    CN310_sign_in(20) <= VN1417_sign_out(4);
    CN310_data_in(21) <= VN1506_data_out(4);
    CN310_sign_in(21) <= VN1506_sign_out(4);
    CN310_data_in(22) <= VN1527_data_out(4);
    CN310_sign_in(22) <= VN1527_sign_out(4);
    CN310_data_in(23) <= VN1694_data_out(4);
    CN310_sign_in(23) <= VN1694_sign_out(4);
    CN310_data_in(24) <= VN1819_data_out(4);
    CN310_sign_in(24) <= VN1819_sign_out(4);
    CN310_data_in(25) <= VN1828_data_out(4);
    CN310_sign_in(25) <= VN1828_sign_out(4);
    CN310_data_in(26) <= VN1860_data_out(4);
    CN310_sign_in(26) <= VN1860_sign_out(4);
    CN310_data_in(27) <= VN1879_data_out(4);
    CN310_sign_in(27) <= VN1879_sign_out(4);
    CN310_data_in(28) <= VN1909_data_out(4);
    CN310_sign_in(28) <= VN1909_sign_out(4);
    CN310_data_in(29) <= VN1937_data_out(4);
    CN310_sign_in(29) <= VN1937_sign_out(4);
    CN310_data_in(30) <= VN1957_data_out(4);
    CN310_sign_in(30) <= VN1957_sign_out(4);
    CN310_data_in(31) <= VN1967_data_out(4);
    CN310_sign_in(31) <= VN1967_sign_out(4);
    CN311_data_in(0) <= VN1_data_out(4);
    CN311_sign_in(0) <= VN1_sign_out(4);
    CN311_data_in(1) <= VN68_data_out(4);
    CN311_sign_in(1) <= VN68_sign_out(4);
    CN311_data_in(2) <= VN160_data_out(4);
    CN311_sign_in(2) <= VN160_sign_out(4);
    CN311_data_in(3) <= VN225_data_out(4);
    CN311_sign_in(3) <= VN225_sign_out(4);
    CN311_data_in(4) <= VN301_data_out(4);
    CN311_sign_in(4) <= VN301_sign_out(4);
    CN311_data_in(5) <= VN387_data_out(4);
    CN311_sign_in(5) <= VN387_sign_out(4);
    CN311_data_in(6) <= VN434_data_out(4);
    CN311_sign_in(6) <= VN434_sign_out(4);
    CN311_data_in(7) <= VN480_data_out(4);
    CN311_sign_in(7) <= VN480_sign_out(4);
    CN311_data_in(8) <= VN511_data_out(4);
    CN311_sign_in(8) <= VN511_sign_out(4);
    CN311_data_in(9) <= VN596_data_out(4);
    CN311_sign_in(9) <= VN596_sign_out(4);
    CN311_data_in(10) <= VN617_data_out(4);
    CN311_sign_in(10) <= VN617_sign_out(4);
    CN311_data_in(11) <= VN706_data_out(4);
    CN311_sign_in(11) <= VN706_sign_out(4);
    CN311_data_in(12) <= VN747_data_out(4);
    CN311_sign_in(12) <= VN747_sign_out(4);
    CN311_data_in(13) <= VN814_data_out(4);
    CN311_sign_in(13) <= VN814_sign_out(4);
    CN311_data_in(14) <= VN862_data_out(4);
    CN311_sign_in(14) <= VN862_sign_out(4);
    CN311_data_in(15) <= VN902_data_out(4);
    CN311_sign_in(15) <= VN902_sign_out(4);
    CN311_data_in(16) <= VN971_data_out(4);
    CN311_sign_in(16) <= VN971_sign_out(4);
    CN311_data_in(17) <= VN1034_data_out(4);
    CN311_sign_in(17) <= VN1034_sign_out(4);
    CN311_data_in(18) <= VN1064_data_out(4);
    CN311_sign_in(18) <= VN1064_sign_out(4);
    CN311_data_in(19) <= VN1157_data_out(4);
    CN311_sign_in(19) <= VN1157_sign_out(4);
    CN311_data_in(20) <= VN1193_data_out(4);
    CN311_sign_in(20) <= VN1193_sign_out(4);
    CN311_data_in(21) <= VN1221_data_out(4);
    CN311_sign_in(21) <= VN1221_sign_out(4);
    CN311_data_in(22) <= VN1310_data_out(4);
    CN311_sign_in(22) <= VN1310_sign_out(4);
    CN311_data_in(23) <= VN1344_data_out(4);
    CN311_sign_in(23) <= VN1344_sign_out(4);
    CN311_data_in(24) <= VN1466_data_out(4);
    CN311_sign_in(24) <= VN1466_sign_out(4);
    CN311_data_in(25) <= VN1523_data_out(4);
    CN311_sign_in(25) <= VN1523_sign_out(4);
    CN311_data_in(26) <= VN1660_data_out(4);
    CN311_sign_in(26) <= VN1660_sign_out(4);
    CN311_data_in(27) <= VN1750_data_out(4);
    CN311_sign_in(27) <= VN1750_sign_out(4);
    CN311_data_in(28) <= VN1760_data_out(4);
    CN311_sign_in(28) <= VN1760_sign_out(4);
    CN311_data_in(29) <= VN1804_data_out(4);
    CN311_sign_in(29) <= VN1804_sign_out(4);
    CN311_data_in(30) <= VN1899_data_out(4);
    CN311_sign_in(30) <= VN1899_sign_out(4);
    CN311_data_in(31) <= VN1913_data_out(4);
    CN311_sign_in(31) <= VN1913_sign_out(4);
    CN312_data_in(0) <= VN0_data_out(4);
    CN312_sign_in(0) <= VN0_sign_out(4);
    CN312_data_in(1) <= VN108_data_out(4);
    CN312_sign_in(1) <= VN108_sign_out(4);
    CN312_data_in(2) <= VN167_data_out(4);
    CN312_sign_in(2) <= VN167_sign_out(4);
    CN312_data_in(3) <= VN246_data_out(4);
    CN312_sign_in(3) <= VN246_sign_out(4);
    CN312_data_in(4) <= VN326_data_out(4);
    CN312_sign_in(4) <= VN326_sign_out(4);
    CN312_data_in(5) <= VN348_data_out(4);
    CN312_sign_in(5) <= VN348_sign_out(4);
    CN312_data_in(6) <= VN452_data_out(4);
    CN312_sign_in(6) <= VN452_sign_out(4);
    CN312_data_in(7) <= VN530_data_out(4);
    CN312_sign_in(7) <= VN530_sign_out(4);
    CN312_data_in(8) <= VN580_data_out(4);
    CN312_sign_in(8) <= VN580_sign_out(4);
    CN312_data_in(9) <= VN645_data_out(4);
    CN312_sign_in(9) <= VN645_sign_out(4);
    CN312_data_in(10) <= VN770_data_out(4);
    CN312_sign_in(10) <= VN770_sign_out(4);
    CN312_data_in(11) <= VN827_data_out(4);
    CN312_sign_in(11) <= VN827_sign_out(4);
    CN312_data_in(12) <= VN838_data_out(4);
    CN312_sign_in(12) <= VN838_sign_out(4);
    CN312_data_in(13) <= VN927_data_out(4);
    CN312_sign_in(13) <= VN927_sign_out(4);
    CN312_data_in(14) <= VN979_data_out(4);
    CN312_sign_in(14) <= VN979_sign_out(4);
    CN312_data_in(15) <= VN1090_data_out(4);
    CN312_sign_in(15) <= VN1090_sign_out(4);
    CN312_data_in(16) <= VN1132_data_out(4);
    CN312_sign_in(16) <= VN1132_sign_out(4);
    CN312_data_in(17) <= VN1182_data_out(4);
    CN312_sign_in(17) <= VN1182_sign_out(4);
    CN312_data_in(18) <= VN1270_data_out(4);
    CN312_sign_in(18) <= VN1270_sign_out(4);
    CN312_data_in(19) <= VN1322_data_out(4);
    CN312_sign_in(19) <= VN1322_sign_out(4);
    CN312_data_in(20) <= VN1342_data_out(4);
    CN312_sign_in(20) <= VN1342_sign_out(4);
    CN312_data_in(21) <= VN1425_data_out(4);
    CN312_sign_in(21) <= VN1425_sign_out(4);
    CN312_data_in(22) <= VN1446_data_out(4);
    CN312_sign_in(22) <= VN1446_sign_out(4);
    CN312_data_in(23) <= VN1482_data_out(4);
    CN312_sign_in(23) <= VN1482_sign_out(4);
    CN312_data_in(24) <= VN1645_data_out(4);
    CN312_sign_in(24) <= VN1645_sign_out(4);
    CN312_data_in(25) <= VN1655_data_out(4);
    CN312_sign_in(25) <= VN1655_sign_out(4);
    CN312_data_in(26) <= VN1698_data_out(4);
    CN312_sign_in(26) <= VN1698_sign_out(4);
    CN312_data_in(27) <= VN1729_data_out(4);
    CN312_sign_in(27) <= VN1729_sign_out(4);
    CN312_data_in(28) <= VN1925_data_out(4);
    CN312_sign_in(28) <= VN1925_sign_out(4);
    CN312_data_in(29) <= VN1969_data_out(4);
    CN312_sign_in(29) <= VN1969_sign_out(4);
    CN312_data_in(30) <= VN2021_data_out(4);
    CN312_sign_in(30) <= VN2021_sign_out(4);
    CN312_data_in(31) <= VN2027_data_out(4);
    CN312_sign_in(31) <= VN2027_sign_out(4);
    CN313_data_in(0) <= VN150_data_out(4);
    CN313_sign_in(0) <= VN150_sign_out(4);
    CN313_data_in(1) <= VN188_data_out(4);
    CN313_sign_in(1) <= VN188_sign_out(4);
    CN313_data_in(2) <= VN247_data_out(4);
    CN313_sign_in(2) <= VN247_sign_out(4);
    CN313_data_in(3) <= VN356_data_out(4);
    CN313_sign_in(3) <= VN356_sign_out(4);
    CN313_data_in(4) <= VN403_data_out(4);
    CN313_sign_in(4) <= VN403_sign_out(4);
    CN313_data_in(5) <= VN496_data_out(4);
    CN313_sign_in(5) <= VN496_sign_out(4);
    CN313_data_in(6) <= VN642_data_out(4);
    CN313_sign_in(6) <= VN642_sign_out(4);
    CN313_data_in(7) <= VN728_data_out(4);
    CN313_sign_in(7) <= VN728_sign_out(4);
    CN313_data_in(8) <= VN886_data_out(4);
    CN313_sign_in(8) <= VN886_sign_out(4);
    CN313_data_in(9) <= VN919_data_out(4);
    CN313_sign_in(9) <= VN919_sign_out(4);
    CN313_data_in(10) <= VN1001_data_out(4);
    CN313_sign_in(10) <= VN1001_sign_out(4);
    CN313_data_in(11) <= VN1050_data_out(4);
    CN313_sign_in(11) <= VN1050_sign_out(4);
    CN313_data_in(12) <= VN1103_data_out(4);
    CN313_sign_in(12) <= VN1103_sign_out(4);
    CN313_data_in(13) <= VN1278_data_out(4);
    CN313_sign_in(13) <= VN1278_sign_out(4);
    CN313_data_in(14) <= VN1376_data_out(4);
    CN313_sign_in(14) <= VN1376_sign_out(4);
    CN313_data_in(15) <= VN1400_data_out(4);
    CN313_sign_in(15) <= VN1400_sign_out(4);
    CN313_data_in(16) <= VN1489_data_out(4);
    CN313_sign_in(16) <= VN1489_sign_out(4);
    CN313_data_in(17) <= VN1528_data_out(4);
    CN313_sign_in(17) <= VN1528_sign_out(4);
    CN313_data_in(18) <= VN1596_data_out(4);
    CN313_sign_in(18) <= VN1596_sign_out(4);
    CN313_data_in(19) <= VN1710_data_out(4);
    CN313_sign_in(19) <= VN1710_sign_out(4);
    CN313_data_in(20) <= VN1723_data_out(4);
    CN313_sign_in(20) <= VN1723_sign_out(4);
    CN313_data_in(21) <= VN1814_data_out(4);
    CN313_sign_in(21) <= VN1814_sign_out(4);
    CN313_data_in(22) <= VN1830_data_out(4);
    CN313_sign_in(22) <= VN1830_sign_out(4);
    CN313_data_in(23) <= VN1881_data_out(4);
    CN313_sign_in(23) <= VN1881_sign_out(4);
    CN313_data_in(24) <= VN1919_data_out(4);
    CN313_sign_in(24) <= VN1919_sign_out(4);
    CN313_data_in(25) <= VN1953_data_out(4);
    CN313_sign_in(25) <= VN1953_sign_out(4);
    CN313_data_in(26) <= VN1973_data_out(4);
    CN313_sign_in(26) <= VN1973_sign_out(4);
    CN313_data_in(27) <= VN1983_data_out(4);
    CN313_sign_in(27) <= VN1983_sign_out(4);
    CN313_data_in(28) <= VN2022_data_out(4);
    CN313_sign_in(28) <= VN2022_sign_out(4);
    CN313_data_in(29) <= VN2034_data_out(4);
    CN313_sign_in(29) <= VN2034_sign_out(4);
    CN313_data_in(30) <= VN2038_data_out(4);
    CN313_sign_in(30) <= VN2038_sign_out(4);
    CN313_data_in(31) <= VN2044_data_out(4);
    CN313_sign_in(31) <= VN2044_sign_out(4);
    CN314_data_in(0) <= VN191_data_out(4);
    CN314_sign_in(0) <= VN191_sign_out(4);
    CN314_data_in(1) <= VN278_data_out(4);
    CN314_sign_in(1) <= VN278_sign_out(4);
    CN314_data_in(2) <= VN316_data_out(4);
    CN314_sign_in(2) <= VN316_sign_out(4);
    CN314_data_in(3) <= VN352_data_out(4);
    CN314_sign_in(3) <= VN352_sign_out(4);
    CN314_data_in(4) <= VN442_data_out(4);
    CN314_sign_in(4) <= VN442_sign_out(4);
    CN314_data_in(5) <= VN483_data_out(4);
    CN314_sign_in(5) <= VN483_sign_out(4);
    CN314_data_in(6) <= VN543_data_out(4);
    CN314_sign_in(6) <= VN543_sign_out(4);
    CN314_data_in(7) <= VN602_data_out(4);
    CN314_sign_in(7) <= VN602_sign_out(4);
    CN314_data_in(8) <= VN656_data_out(4);
    CN314_sign_in(8) <= VN656_sign_out(4);
    CN314_data_in(9) <= VN687_data_out(4);
    CN314_sign_in(9) <= VN687_sign_out(4);
    CN314_data_in(10) <= VN781_data_out(4);
    CN314_sign_in(10) <= VN781_sign_out(4);
    CN314_data_in(11) <= VN848_data_out(4);
    CN314_sign_in(11) <= VN848_sign_out(4);
    CN314_data_in(12) <= VN907_data_out(4);
    CN314_sign_in(12) <= VN907_sign_out(4);
    CN314_data_in(13) <= VN1053_data_out(4);
    CN314_sign_in(13) <= VN1053_sign_out(4);
    CN314_data_in(14) <= VN1123_data_out(4);
    CN314_sign_in(14) <= VN1123_sign_out(4);
    CN314_data_in(15) <= VN1357_data_out(4);
    CN314_sign_in(15) <= VN1357_sign_out(4);
    CN314_data_in(16) <= VN1389_data_out(4);
    CN314_sign_in(16) <= VN1389_sign_out(4);
    CN314_data_in(17) <= VN1411_data_out(4);
    CN314_sign_in(17) <= VN1411_sign_out(4);
    CN314_data_in(18) <= VN1461_data_out(4);
    CN314_sign_in(18) <= VN1461_sign_out(4);
    CN314_data_in(19) <= VN1556_data_out(4);
    CN314_sign_in(19) <= VN1556_sign_out(4);
    CN314_data_in(20) <= VN1648_data_out(4);
    CN314_sign_in(20) <= VN1648_sign_out(4);
    CN314_data_in(21) <= VN1651_data_out(4);
    CN314_sign_in(21) <= VN1651_sign_out(4);
    CN314_data_in(22) <= VN1717_data_out(4);
    CN314_sign_in(22) <= VN1717_sign_out(4);
    CN314_data_in(23) <= VN1749_data_out(4);
    CN314_sign_in(23) <= VN1749_sign_out(4);
    CN314_data_in(24) <= VN1836_data_out(4);
    CN314_sign_in(24) <= VN1836_sign_out(4);
    CN314_data_in(25) <= VN1853_data_out(4);
    CN314_sign_in(25) <= VN1853_sign_out(4);
    CN314_data_in(26) <= VN1907_data_out(4);
    CN314_sign_in(26) <= VN1907_sign_out(4);
    CN314_data_in(27) <= VN1926_data_out(4);
    CN314_sign_in(27) <= VN1926_sign_out(4);
    CN314_data_in(28) <= VN1928_data_out(4);
    CN314_sign_in(28) <= VN1928_sign_out(4);
    CN314_data_in(29) <= VN1938_data_out(4);
    CN314_sign_in(29) <= VN1938_sign_out(4);
    CN314_data_in(30) <= VN1958_data_out(4);
    CN314_sign_in(30) <= VN1958_sign_out(4);
    CN314_data_in(31) <= VN1968_data_out(4);
    CN314_sign_in(31) <= VN1968_sign_out(4);
    CN315_data_in(0) <= VN78_data_out(4);
    CN315_sign_in(0) <= VN78_sign_out(4);
    CN315_data_in(1) <= VN119_data_out(4);
    CN315_sign_in(1) <= VN119_sign_out(4);
    CN315_data_in(2) <= VN183_data_out(4);
    CN315_sign_in(2) <= VN183_sign_out(4);
    CN315_data_in(3) <= VN271_data_out(4);
    CN315_sign_in(3) <= VN271_sign_out(4);
    CN315_data_in(4) <= VN318_data_out(4);
    CN315_sign_in(4) <= VN318_sign_out(4);
    CN315_data_in(5) <= VN357_data_out(4);
    CN315_sign_in(5) <= VN357_sign_out(4);
    CN315_data_in(6) <= VN399_data_out(4);
    CN315_sign_in(6) <= VN399_sign_out(4);
    CN315_data_in(7) <= VN499_data_out(4);
    CN315_sign_in(7) <= VN499_sign_out(4);
    CN315_data_in(8) <= VN513_data_out(4);
    CN315_sign_in(8) <= VN513_sign_out(4);
    CN315_data_in(9) <= VN575_data_out(4);
    CN315_sign_in(9) <= VN575_sign_out(4);
    CN315_data_in(10) <= VN651_data_out(4);
    CN315_sign_in(10) <= VN651_sign_out(4);
    CN315_data_in(11) <= VN678_data_out(4);
    CN315_sign_in(11) <= VN678_sign_out(4);
    CN315_data_in(12) <= VN743_data_out(4);
    CN315_sign_in(12) <= VN743_sign_out(4);
    CN315_data_in(13) <= VN802_data_out(4);
    CN315_sign_in(13) <= VN802_sign_out(4);
    CN315_data_in(14) <= VN853_data_out(4);
    CN315_sign_in(14) <= VN853_sign_out(4);
    CN315_data_in(15) <= VN924_data_out(4);
    CN315_sign_in(15) <= VN924_sign_out(4);
    CN315_data_in(16) <= VN977_data_out(4);
    CN315_sign_in(16) <= VN977_sign_out(4);
    CN315_data_in(17) <= VN1037_data_out(4);
    CN315_sign_in(17) <= VN1037_sign_out(4);
    CN315_data_in(18) <= VN1111_data_out(4);
    CN315_sign_in(18) <= VN1111_sign_out(4);
    CN315_data_in(19) <= VN1172_data_out(4);
    CN315_sign_in(19) <= VN1172_sign_out(4);
    CN315_data_in(20) <= VN1249_data_out(4);
    CN315_sign_in(20) <= VN1249_sign_out(4);
    CN315_data_in(21) <= VN1317_data_out(4);
    CN315_sign_in(21) <= VN1317_sign_out(4);
    CN315_data_in(22) <= VN1359_data_out(4);
    CN315_sign_in(22) <= VN1359_sign_out(4);
    CN315_data_in(23) <= VN1404_data_out(4);
    CN315_sign_in(23) <= VN1404_sign_out(4);
    CN315_data_in(24) <= VN1447_data_out(4);
    CN315_sign_in(24) <= VN1447_sign_out(4);
    CN315_data_in(25) <= VN1457_data_out(4);
    CN315_sign_in(25) <= VN1457_sign_out(4);
    CN315_data_in(26) <= VN1488_data_out(4);
    CN315_sign_in(26) <= VN1488_sign_out(4);
    CN315_data_in(27) <= VN1511_data_out(4);
    CN315_sign_in(27) <= VN1511_sign_out(4);
    CN315_data_in(28) <= VN1675_data_out(4);
    CN315_sign_in(28) <= VN1675_sign_out(4);
    CN315_data_in(29) <= VN1714_data_out(4);
    CN315_sign_in(29) <= VN1714_sign_out(4);
    CN315_data_in(30) <= VN1722_data_out(4);
    CN315_sign_in(30) <= VN1722_sign_out(4);
    CN315_data_in(31) <= VN1799_data_out(4);
    CN315_sign_in(31) <= VN1799_sign_out(4);
    CN316_data_in(0) <= VN61_data_out(4);
    CN316_sign_in(0) <= VN61_sign_out(4);
    CN316_data_in(1) <= VN158_data_out(4);
    CN316_sign_in(1) <= VN158_sign_out(4);
    CN316_data_in(2) <= VN234_data_out(4);
    CN316_sign_in(2) <= VN234_sign_out(4);
    CN316_data_in(3) <= VN288_data_out(4);
    CN316_sign_in(3) <= VN288_sign_out(4);
    CN316_data_in(4) <= VN347_data_out(4);
    CN316_sign_in(4) <= VN347_sign_out(4);
    CN316_data_in(5) <= VN560_data_out(4);
    CN316_sign_in(5) <= VN560_sign_out(4);
    CN316_data_in(6) <= VN563_data_out(4);
    CN316_sign_in(6) <= VN563_sign_out(4);
    CN316_data_in(7) <= VN625_data_out(4);
    CN316_sign_in(7) <= VN625_sign_out(4);
    CN316_data_in(8) <= VN720_data_out(4);
    CN316_sign_in(8) <= VN720_sign_out(4);
    CN316_data_in(9) <= VN764_data_out(4);
    CN316_sign_in(9) <= VN764_sign_out(4);
    CN316_data_in(10) <= VN816_data_out(4);
    CN316_sign_in(10) <= VN816_sign_out(4);
    CN316_data_in(11) <= VN898_data_out(4);
    CN316_sign_in(11) <= VN898_sign_out(4);
    CN316_data_in(12) <= VN956_data_out(4);
    CN316_sign_in(12) <= VN956_sign_out(4);
    CN316_data_in(13) <= VN1014_data_out(4);
    CN316_sign_in(13) <= VN1014_sign_out(4);
    CN316_data_in(14) <= VN1080_data_out(4);
    CN316_sign_in(14) <= VN1080_sign_out(4);
    CN316_data_in(15) <= VN1134_data_out(4);
    CN316_sign_in(15) <= VN1134_sign_out(4);
    CN316_data_in(16) <= VN1186_data_out(4);
    CN316_sign_in(16) <= VN1186_sign_out(4);
    CN316_data_in(17) <= VN1220_data_out(4);
    CN316_sign_in(17) <= VN1220_sign_out(4);
    CN316_data_in(18) <= VN1246_data_out(4);
    CN316_sign_in(18) <= VN1246_sign_out(4);
    CN316_data_in(19) <= VN1293_data_out(4);
    CN316_sign_in(19) <= VN1293_sign_out(4);
    CN316_data_in(20) <= VN1345_data_out(4);
    CN316_sign_in(20) <= VN1345_sign_out(4);
    CN316_data_in(21) <= VN1408_data_out(4);
    CN316_sign_in(21) <= VN1408_sign_out(4);
    CN316_data_in(22) <= VN1501_data_out(4);
    CN316_sign_in(22) <= VN1501_sign_out(4);
    CN316_data_in(23) <= VN1569_data_out(4);
    CN316_sign_in(23) <= VN1569_sign_out(4);
    CN316_data_in(24) <= VN1664_data_out(4);
    CN316_sign_in(24) <= VN1664_sign_out(4);
    CN316_data_in(25) <= VN1721_data_out(4);
    CN316_sign_in(25) <= VN1721_sign_out(4);
    CN316_data_in(26) <= VN1727_data_out(4);
    CN316_sign_in(26) <= VN1727_sign_out(4);
    CN316_data_in(27) <= VN1754_data_out(4);
    CN316_sign_in(27) <= VN1754_sign_out(4);
    CN316_data_in(28) <= VN1961_data_out(4);
    CN316_sign_in(28) <= VN1961_sign_out(4);
    CN316_data_in(29) <= VN2014_data_out(4);
    CN316_sign_in(29) <= VN2014_sign_out(4);
    CN316_data_in(30) <= VN2035_data_out(4);
    CN316_sign_in(30) <= VN2035_sign_out(4);
    CN316_data_in(31) <= VN2039_data_out(4);
    CN316_sign_in(31) <= VN2039_sign_out(4);
    CN317_data_in(0) <= VN88_data_out(4);
    CN317_sign_in(0) <= VN88_sign_out(4);
    CN317_data_in(1) <= VN238_data_out(4);
    CN317_sign_in(1) <= VN238_sign_out(4);
    CN317_data_in(2) <= VN324_data_out(4);
    CN317_sign_in(2) <= VN324_sign_out(4);
    CN317_data_in(3) <= VN372_data_out(4);
    CN317_sign_in(3) <= VN372_sign_out(4);
    CN317_data_in(4) <= VN472_data_out(4);
    CN317_sign_in(4) <= VN472_sign_out(4);
    CN317_data_in(5) <= VN548_data_out(4);
    CN317_sign_in(5) <= VN548_sign_out(4);
    CN317_data_in(6) <= VN604_data_out(4);
    CN317_sign_in(6) <= VN604_sign_out(4);
    CN317_data_in(7) <= VN634_data_out(4);
    CN317_sign_in(7) <= VN634_sign_out(4);
    CN317_data_in(8) <= VN683_data_out(4);
    CN317_sign_in(8) <= VN683_sign_out(4);
    CN317_data_in(9) <= VN765_data_out(4);
    CN317_sign_in(9) <= VN765_sign_out(4);
    CN317_data_in(10) <= VN812_data_out(4);
    CN317_sign_in(10) <= VN812_sign_out(4);
    CN317_data_in(11) <= VN852_data_out(4);
    CN317_sign_in(11) <= VN852_sign_out(4);
    CN317_data_in(12) <= VN895_data_out(4);
    CN317_sign_in(12) <= VN895_sign_out(4);
    CN317_data_in(13) <= VN959_data_out(4);
    CN317_sign_in(13) <= VN959_sign_out(4);
    CN317_data_in(14) <= VN1092_data_out(4);
    CN317_sign_in(14) <= VN1092_sign_out(4);
    CN317_data_in(15) <= VN1125_data_out(4);
    CN317_sign_in(15) <= VN1125_sign_out(4);
    CN317_data_in(16) <= VN1179_data_out(4);
    CN317_sign_in(16) <= VN1179_sign_out(4);
    CN317_data_in(17) <= VN1261_data_out(4);
    CN317_sign_in(17) <= VN1261_sign_out(4);
    CN317_data_in(18) <= VN1325_data_out(4);
    CN317_sign_in(18) <= VN1325_sign_out(4);
    CN317_data_in(19) <= VN1332_data_out(4);
    CN317_sign_in(19) <= VN1332_sign_out(4);
    CN317_data_in(20) <= VN1377_data_out(4);
    CN317_sign_in(20) <= VN1377_sign_out(4);
    CN317_data_in(21) <= VN1397_data_out(4);
    CN317_sign_in(21) <= VN1397_sign_out(4);
    CN317_data_in(22) <= VN1719_data_out(4);
    CN317_sign_in(22) <= VN1719_sign_out(4);
    CN317_data_in(23) <= VN1775_data_out(4);
    CN317_sign_in(23) <= VN1775_sign_out(4);
    CN317_data_in(24) <= VN1811_data_out(4);
    CN317_sign_in(24) <= VN1811_sign_out(4);
    CN317_data_in(25) <= VN1839_data_out(4);
    CN317_sign_in(25) <= VN1839_sign_out(4);
    CN317_data_in(26) <= VN1939_data_out(4);
    CN317_sign_in(26) <= VN1939_sign_out(4);
    CN317_data_in(27) <= VN1952_data_out(4);
    CN317_sign_in(27) <= VN1952_sign_out(4);
    CN317_data_in(28) <= VN1960_data_out(4);
    CN317_sign_in(28) <= VN1960_sign_out(4);
    CN317_data_in(29) <= VN1999_data_out(4);
    CN317_sign_in(29) <= VN1999_sign_out(4);
    CN317_data_in(30) <= VN2001_data_out(4);
    CN317_sign_in(30) <= VN2001_sign_out(4);
    CN317_data_in(31) <= VN2012_data_out(4);
    CN317_sign_in(31) <= VN2012_sign_out(4);
    CN318_data_in(0) <= VN120_data_out(4);
    CN318_sign_in(0) <= VN120_sign_out(4);
    CN318_data_in(1) <= VN210_data_out(4);
    CN318_sign_in(1) <= VN210_sign_out(4);
    CN318_data_in(2) <= VN279_data_out(4);
    CN318_sign_in(2) <= VN279_sign_out(4);
    CN318_data_in(3) <= VN379_data_out(4);
    CN318_sign_in(3) <= VN379_sign_out(4);
    CN318_data_in(4) <= VN425_data_out(4);
    CN318_sign_in(4) <= VN425_sign_out(4);
    CN318_data_in(5) <= VN467_data_out(4);
    CN318_sign_in(5) <= VN467_sign_out(4);
    CN318_data_in(6) <= VN566_data_out(4);
    CN318_sign_in(6) <= VN566_sign_out(4);
    CN318_data_in(7) <= VN742_data_out(4);
    CN318_sign_in(7) <= VN742_sign_out(4);
    CN318_data_in(8) <= VN846_data_out(4);
    CN318_sign_in(8) <= VN846_sign_out(4);
    CN318_data_in(9) <= VN911_data_out(4);
    CN318_sign_in(9) <= VN911_sign_out(4);
    CN318_data_in(10) <= VN1002_data_out(4);
    CN318_sign_in(10) <= VN1002_sign_out(4);
    CN318_data_in(11) <= VN1006_data_out(4);
    CN318_sign_in(11) <= VN1006_sign_out(4);
    CN318_data_in(12) <= VN1059_data_out(4);
    CN318_sign_in(12) <= VN1059_sign_out(4);
    CN318_data_in(13) <= VN1210_data_out(4);
    CN318_sign_in(13) <= VN1210_sign_out(4);
    CN318_data_in(14) <= VN1295_data_out(4);
    CN318_sign_in(14) <= VN1295_sign_out(4);
    CN318_data_in(15) <= VN1341_data_out(4);
    CN318_sign_in(15) <= VN1341_sign_out(4);
    CN318_data_in(16) <= VN1540_data_out(4);
    CN318_sign_in(16) <= VN1540_sign_out(4);
    CN318_data_in(17) <= VN1566_data_out(4);
    CN318_sign_in(17) <= VN1566_sign_out(4);
    CN318_data_in(18) <= VN1598_data_out(4);
    CN318_sign_in(18) <= VN1598_sign_out(4);
    CN318_data_in(19) <= VN1634_data_out(4);
    CN318_sign_in(19) <= VN1634_sign_out(4);
    CN318_data_in(20) <= VN1720_data_out(4);
    CN318_sign_in(20) <= VN1720_sign_out(4);
    CN318_data_in(21) <= VN1805_data_out(4);
    CN318_sign_in(21) <= VN1805_sign_out(4);
    CN318_data_in(22) <= VN1837_data_out(4);
    CN318_sign_in(22) <= VN1837_sign_out(4);
    CN318_data_in(23) <= VN1877_data_out(4);
    CN318_sign_in(23) <= VN1877_sign_out(4);
    CN318_data_in(24) <= VN1935_data_out(4);
    CN318_sign_in(24) <= VN1935_sign_out(4);
    CN318_data_in(25) <= VN1976_data_out(4);
    CN318_sign_in(25) <= VN1976_sign_out(4);
    CN318_data_in(26) <= VN1980_data_out(4);
    CN318_sign_in(26) <= VN1980_sign_out(4);
    CN318_data_in(27) <= VN2005_data_out(4);
    CN318_sign_in(27) <= VN2005_sign_out(4);
    CN318_data_in(28) <= VN2008_data_out(4);
    CN318_sign_in(28) <= VN2008_sign_out(4);
    CN318_data_in(29) <= VN2036_data_out(4);
    CN318_sign_in(29) <= VN2036_sign_out(4);
    CN318_data_in(30) <= VN2037_data_out(4);
    CN318_sign_in(30) <= VN2037_sign_out(4);
    CN318_data_in(31) <= VN2045_data_out(4);
    CN318_sign_in(31) <= VN2045_sign_out(4);
    CN319_data_in(0) <= VN52_data_out(4);
    CN319_sign_in(0) <= VN52_sign_out(4);
    CN319_data_in(1) <= VN66_data_out(4);
    CN319_sign_in(1) <= VN66_sign_out(4);
    CN319_data_in(2) <= VN151_data_out(4);
    CN319_sign_in(2) <= VN151_sign_out(4);
    CN319_data_in(3) <= VN221_data_out(4);
    CN319_sign_in(3) <= VN221_sign_out(4);
    CN319_data_in(4) <= VN237_data_out(4);
    CN319_sign_in(4) <= VN237_sign_out(4);
    CN319_data_in(5) <= VN289_data_out(4);
    CN319_sign_in(5) <= VN289_sign_out(4);
    CN319_data_in(6) <= VN361_data_out(4);
    CN319_sign_in(6) <= VN361_sign_out(4);
    CN319_data_in(7) <= VN411_data_out(4);
    CN319_sign_in(7) <= VN411_sign_out(4);
    CN319_data_in(8) <= VN473_data_out(4);
    CN319_sign_in(8) <= VN473_sign_out(4);
    CN319_data_in(9) <= VN539_data_out(4);
    CN319_sign_in(9) <= VN539_sign_out(4);
    CN319_data_in(10) <= VN585_data_out(4);
    CN319_sign_in(10) <= VN585_sign_out(4);
    CN319_data_in(11) <= VN631_data_out(4);
    CN319_sign_in(11) <= VN631_sign_out(4);
    CN319_data_in(12) <= VN711_data_out(4);
    CN319_sign_in(12) <= VN711_sign_out(4);
    CN319_data_in(13) <= VN734_data_out(4);
    CN319_sign_in(13) <= VN734_sign_out(4);
    CN319_data_in(14) <= VN797_data_out(4);
    CN319_sign_in(14) <= VN797_sign_out(4);
    CN319_data_in(15) <= VN883_data_out(4);
    CN319_sign_in(15) <= VN883_sign_out(4);
    CN319_data_in(16) <= VN904_data_out(4);
    CN319_sign_in(16) <= VN904_sign_out(4);
    CN319_data_in(17) <= VN978_data_out(4);
    CN319_sign_in(17) <= VN978_sign_out(4);
    CN319_data_in(18) <= VN1046_data_out(4);
    CN319_sign_in(18) <= VN1046_sign_out(4);
    CN319_data_in(19) <= VN1106_data_out(4);
    CN319_sign_in(19) <= VN1106_sign_out(4);
    CN319_data_in(20) <= VN1130_data_out(4);
    CN319_sign_in(20) <= VN1130_sign_out(4);
    CN319_data_in(21) <= VN1231_data_out(4);
    CN319_sign_in(21) <= VN1231_sign_out(4);
    CN319_data_in(22) <= VN1305_data_out(4);
    CN319_sign_in(22) <= VN1305_sign_out(4);
    CN319_data_in(23) <= VN1368_data_out(4);
    CN319_sign_in(23) <= VN1368_sign_out(4);
    CN319_data_in(24) <= VN1416_data_out(4);
    CN319_sign_in(24) <= VN1416_sign_out(4);
    CN319_data_in(25) <= VN1475_data_out(4);
    CN319_sign_in(25) <= VN1475_sign_out(4);
    CN319_data_in(26) <= VN1485_data_out(4);
    CN319_sign_in(26) <= VN1485_sign_out(4);
    CN319_data_in(27) <= VN1515_data_out(4);
    CN319_sign_in(27) <= VN1515_sign_out(4);
    CN319_data_in(28) <= VN1595_data_out(4);
    CN319_sign_in(28) <= VN1595_sign_out(4);
    CN319_data_in(29) <= VN1661_data_out(4);
    CN319_sign_in(29) <= VN1661_sign_out(4);
    CN319_data_in(30) <= VN1695_data_out(4);
    CN319_sign_in(30) <= VN1695_sign_out(4);
    CN319_data_in(31) <= VN1800_data_out(4);
    CN319_sign_in(31) <= VN1800_sign_out(4);
    CN320_data_in(0) <= VN53_data_out(5);
    CN320_sign_in(0) <= VN53_sign_out(5);
    CN320_data_in(1) <= VN126_data_out(5);
    CN320_sign_in(1) <= VN126_sign_out(5);
    CN320_data_in(2) <= VN196_data_out(5);
    CN320_sign_in(2) <= VN196_sign_out(5);
    CN320_data_in(3) <= VN295_data_out(5);
    CN320_sign_in(3) <= VN295_sign_out(5);
    CN320_data_in(4) <= VN338_data_out(5);
    CN320_sign_in(4) <= VN338_sign_out(5);
    CN320_data_in(5) <= VN439_data_out(5);
    CN320_sign_in(5) <= VN439_sign_out(5);
    CN320_data_in(6) <= VN454_data_out(5);
    CN320_sign_in(6) <= VN454_sign_out(5);
    CN320_data_in(7) <= VN531_data_out(5);
    CN320_sign_in(7) <= VN531_sign_out(5);
    CN320_data_in(8) <= VN577_data_out(5);
    CN320_sign_in(8) <= VN577_sign_out(5);
    CN320_data_in(9) <= VN637_data_out(5);
    CN320_sign_in(9) <= VN637_sign_out(5);
    CN320_data_in(10) <= VN707_data_out(5);
    CN320_sign_in(10) <= VN707_sign_out(5);
    CN320_data_in(11) <= VN759_data_out(5);
    CN320_sign_in(11) <= VN759_sign_out(5);
    CN320_data_in(12) <= VN792_data_out(5);
    CN320_sign_in(12) <= VN792_sign_out(5);
    CN320_data_in(13) <= VN856_data_out(5);
    CN320_sign_in(13) <= VN856_sign_out(5);
    CN320_data_in(14) <= VN890_data_out(5);
    CN320_sign_in(14) <= VN890_sign_out(5);
    CN320_data_in(15) <= VN1034_data_out(5);
    CN320_sign_in(15) <= VN1034_sign_out(5);
    CN320_data_in(16) <= VN1070_data_out(5);
    CN320_sign_in(16) <= VN1070_sign_out(5);
    CN320_data_in(17) <= VN1154_data_out(5);
    CN320_sign_in(17) <= VN1154_sign_out(5);
    CN320_data_in(18) <= VN1342_data_out(5);
    CN320_sign_in(18) <= VN1342_sign_out(5);
    CN320_data_in(19) <= VN1413_data_out(5);
    CN320_sign_in(19) <= VN1413_sign_out(5);
    CN320_data_in(20) <= VN1453_data_out(5);
    CN320_sign_in(20) <= VN1453_sign_out(5);
    CN320_data_in(21) <= VN1484_data_out(5);
    CN320_sign_in(21) <= VN1484_sign_out(5);
    CN320_data_in(22) <= VN1572_data_out(5);
    CN320_sign_in(22) <= VN1572_sign_out(5);
    CN320_data_in(23) <= VN1579_data_out(5);
    CN320_sign_in(23) <= VN1579_sign_out(5);
    CN320_data_in(24) <= VN1662_data_out(5);
    CN320_sign_in(24) <= VN1662_sign_out(5);
    CN320_data_in(25) <= VN1725_data_out(5);
    CN320_sign_in(25) <= VN1725_sign_out(5);
    CN320_data_in(26) <= VN1741_data_out(5);
    CN320_sign_in(26) <= VN1741_sign_out(5);
    CN320_data_in(27) <= VN1761_data_out(5);
    CN320_sign_in(27) <= VN1761_sign_out(5);
    CN320_data_in(28) <= VN1816_data_out(5);
    CN320_sign_in(28) <= VN1816_sign_out(5);
    CN320_data_in(29) <= VN1836_data_out(5);
    CN320_sign_in(29) <= VN1836_sign_out(5);
    CN320_data_in(30) <= VN1856_data_out(5);
    CN320_sign_in(30) <= VN1856_sign_out(5);
    CN320_data_in(31) <= VN1895_data_out(5);
    CN320_sign_in(31) <= VN1895_sign_out(5);
    CN321_data_in(0) <= VN51_data_out(5);
    CN321_sign_in(0) <= VN51_sign_out(5);
    CN321_data_in(1) <= VN65_data_out(5);
    CN321_sign_in(1) <= VN65_sign_out(5);
    CN321_data_in(2) <= VN150_data_out(5);
    CN321_sign_in(2) <= VN150_sign_out(5);
    CN321_data_in(3) <= VN220_data_out(5);
    CN321_sign_in(3) <= VN220_sign_out(5);
    CN321_data_in(4) <= VN236_data_out(5);
    CN321_sign_in(4) <= VN236_sign_out(5);
    CN321_data_in(5) <= VN288_data_out(5);
    CN321_sign_in(5) <= VN288_sign_out(5);
    CN321_data_in(6) <= VN360_data_out(5);
    CN321_sign_in(6) <= VN360_sign_out(5);
    CN321_data_in(7) <= VN410_data_out(5);
    CN321_sign_in(7) <= VN410_sign_out(5);
    CN321_data_in(8) <= VN472_data_out(5);
    CN321_sign_in(8) <= VN472_sign_out(5);
    CN321_data_in(9) <= VN538_data_out(5);
    CN321_sign_in(9) <= VN538_sign_out(5);
    CN321_data_in(10) <= VN584_data_out(5);
    CN321_sign_in(10) <= VN584_sign_out(5);
    CN321_data_in(11) <= VN630_data_out(5);
    CN321_sign_in(11) <= VN630_sign_out(5);
    CN321_data_in(12) <= VN733_data_out(5);
    CN321_sign_in(12) <= VN733_sign_out(5);
    CN321_data_in(13) <= VN882_data_out(5);
    CN321_sign_in(13) <= VN882_sign_out(5);
    CN321_data_in(14) <= VN903_data_out(5);
    CN321_sign_in(14) <= VN903_sign_out(5);
    CN321_data_in(15) <= VN977_data_out(5);
    CN321_sign_in(15) <= VN977_sign_out(5);
    CN321_data_in(16) <= VN1045_data_out(5);
    CN321_sign_in(16) <= VN1045_sign_out(5);
    CN321_data_in(17) <= VN1105_data_out(5);
    CN321_sign_in(17) <= VN1105_sign_out(5);
    CN321_data_in(18) <= VN1217_data_out(5);
    CN321_sign_in(18) <= VN1217_sign_out(5);
    CN321_data_in(19) <= VN1230_data_out(5);
    CN321_sign_in(19) <= VN1230_sign_out(5);
    CN321_data_in(20) <= VN1304_data_out(5);
    CN321_sign_in(20) <= VN1304_sign_out(5);
    CN321_data_in(21) <= VN1367_data_out(5);
    CN321_sign_in(21) <= VN1367_sign_out(5);
    CN321_data_in(22) <= VN1474_data_out(5);
    CN321_sign_in(22) <= VN1474_sign_out(5);
    CN321_data_in(23) <= VN1558_data_out(5);
    CN321_sign_in(23) <= VN1558_sign_out(5);
    CN321_data_in(24) <= VN1594_data_out(5);
    CN321_sign_in(24) <= VN1594_sign_out(5);
    CN321_data_in(25) <= VN1660_data_out(5);
    CN321_sign_in(25) <= VN1660_sign_out(5);
    CN321_data_in(26) <= VN1759_data_out(5);
    CN321_sign_in(26) <= VN1759_sign_out(5);
    CN321_data_in(27) <= VN1831_data_out(5);
    CN321_sign_in(27) <= VN1831_sign_out(5);
    CN321_data_in(28) <= VN1929_data_out(5);
    CN321_sign_in(28) <= VN1929_sign_out(5);
    CN321_data_in(29) <= VN1992_data_out(5);
    CN321_sign_in(29) <= VN1992_sign_out(5);
    CN321_data_in(30) <= VN2003_data_out(5);
    CN321_sign_in(30) <= VN2003_sign_out(5);
    CN321_data_in(31) <= VN2013_data_out(5);
    CN321_sign_in(31) <= VN2013_sign_out(5);
    CN322_data_in(0) <= VN50_data_out(5);
    CN322_sign_in(0) <= VN50_sign_out(5);
    CN322_data_in(1) <= VN84_data_out(5);
    CN322_sign_in(1) <= VN84_sign_out(5);
    CN322_data_in(2) <= VN165_data_out(5);
    CN322_sign_in(2) <= VN165_sign_out(5);
    CN322_data_in(3) <= VN231_data_out(5);
    CN322_sign_in(3) <= VN231_sign_out(5);
    CN322_data_in(4) <= VN316_data_out(5);
    CN322_sign_in(4) <= VN316_sign_out(5);
    CN322_data_in(5) <= VN362_data_out(5);
    CN322_sign_in(5) <= VN362_sign_out(5);
    CN322_data_in(6) <= VN427_data_out(5);
    CN322_sign_in(6) <= VN427_sign_out(5);
    CN322_data_in(7) <= VN462_data_out(5);
    CN322_sign_in(7) <= VN462_sign_out(5);
    CN322_data_in(8) <= VN535_data_out(5);
    CN322_sign_in(8) <= VN535_sign_out(5);
    CN322_data_in(9) <= VN592_data_out(5);
    CN322_sign_in(9) <= VN592_sign_out(5);
    CN322_data_in(10) <= VN623_data_out(5);
    CN322_sign_in(10) <= VN623_sign_out(5);
    CN322_data_in(11) <= VN749_data_out(5);
    CN322_sign_in(11) <= VN749_sign_out(5);
    CN322_data_in(12) <= VN797_data_out(5);
    CN322_sign_in(12) <= VN797_sign_out(5);
    CN322_data_in(13) <= VN834_data_out(5);
    CN322_sign_in(13) <= VN834_sign_out(5);
    CN322_data_in(14) <= VN932_data_out(5);
    CN322_sign_in(14) <= VN932_sign_out(5);
    CN322_data_in(15) <= VN998_data_out(5);
    CN322_sign_in(15) <= VN998_sign_out(5);
    CN322_data_in(16) <= VN1015_data_out(5);
    CN322_sign_in(16) <= VN1015_sign_out(5);
    CN322_data_in(17) <= VN1060_data_out(5);
    CN322_sign_in(17) <= VN1060_sign_out(5);
    CN322_data_in(18) <= VN1075_data_out(5);
    CN322_sign_in(18) <= VN1075_sign_out(5);
    CN322_data_in(19) <= VN1161_data_out(5);
    CN322_sign_in(19) <= VN1161_sign_out(5);
    CN322_data_in(20) <= VN1302_data_out(5);
    CN322_sign_in(20) <= VN1302_sign_out(5);
    CN322_data_in(21) <= VN1353_data_out(5);
    CN322_sign_in(21) <= VN1353_sign_out(5);
    CN322_data_in(22) <= VN1463_data_out(5);
    CN322_sign_in(22) <= VN1463_sign_out(5);
    CN322_data_in(23) <= VN1492_data_out(5);
    CN322_sign_in(23) <= VN1492_sign_out(5);
    CN322_data_in(24) <= VN1537_data_out(5);
    CN322_sign_in(24) <= VN1537_sign_out(5);
    CN322_data_in(25) <= VN1756_data_out(5);
    CN322_sign_in(25) <= VN1756_sign_out(5);
    CN322_data_in(26) <= VN1813_data_out(5);
    CN322_sign_in(26) <= VN1813_sign_out(5);
    CN322_data_in(27) <= VN1868_data_out(5);
    CN322_sign_in(27) <= VN1868_sign_out(5);
    CN322_data_in(28) <= VN1878_data_out(5);
    CN322_sign_in(28) <= VN1878_sign_out(5);
    CN322_data_in(29) <= VN1911_data_out(5);
    CN322_sign_in(29) <= VN1911_sign_out(5);
    CN322_data_in(30) <= VN1953_data_out(5);
    CN322_sign_in(30) <= VN1953_sign_out(5);
    CN322_data_in(31) <= VN1969_data_out(5);
    CN322_sign_in(31) <= VN1969_sign_out(5);
    CN323_data_in(0) <= VN56_data_out(5);
    CN323_sign_in(0) <= VN56_sign_out(5);
    CN323_data_in(1) <= VN136_data_out(5);
    CN323_sign_in(1) <= VN136_sign_out(5);
    CN323_data_in(2) <= VN184_data_out(5);
    CN323_sign_in(2) <= VN184_sign_out(5);
    CN323_data_in(3) <= VN268_data_out(5);
    CN323_sign_in(3) <= VN268_sign_out(5);
    CN323_data_in(4) <= VN330_data_out(5);
    CN323_sign_in(4) <= VN330_sign_out(5);
    CN323_data_in(5) <= VN390_data_out(5);
    CN323_sign_in(5) <= VN390_sign_out(5);
    CN323_data_in(6) <= VN392_data_out(5);
    CN323_sign_in(6) <= VN392_sign_out(5);
    CN323_data_in(7) <= VN484_data_out(5);
    CN323_sign_in(7) <= VN484_sign_out(5);
    CN323_data_in(8) <= VN552_data_out(5);
    CN323_sign_in(8) <= VN552_sign_out(5);
    CN323_data_in(9) <= VN588_data_out(5);
    CN323_sign_in(9) <= VN588_sign_out(5);
    CN323_data_in(10) <= VN656_data_out(5);
    CN323_sign_in(10) <= VN656_sign_out(5);
    CN323_data_in(11) <= VN717_data_out(5);
    CN323_sign_in(11) <= VN717_sign_out(5);
    CN323_data_in(12) <= VN754_data_out(5);
    CN323_sign_in(12) <= VN754_sign_out(5);
    CN323_data_in(13) <= VN828_data_out(5);
    CN323_sign_in(13) <= VN828_sign_out(5);
    CN323_data_in(14) <= VN967_data_out(5);
    CN323_sign_in(14) <= VN967_sign_out(5);
    CN323_data_in(15) <= VN1007_data_out(5);
    CN323_sign_in(15) <= VN1007_sign_out(5);
    CN323_data_in(16) <= VN1076_data_out(5);
    CN323_sign_in(16) <= VN1076_sign_out(5);
    CN323_data_in(17) <= VN1158_data_out(5);
    CN323_sign_in(17) <= VN1158_sign_out(5);
    CN323_data_in(18) <= VN1221_data_out(5);
    CN323_sign_in(18) <= VN1221_sign_out(5);
    CN323_data_in(19) <= VN1234_data_out(5);
    CN323_sign_in(19) <= VN1234_sign_out(5);
    CN323_data_in(20) <= VN1319_data_out(5);
    CN323_sign_in(20) <= VN1319_sign_out(5);
    CN323_data_in(21) <= VN1546_data_out(5);
    CN323_sign_in(21) <= VN1546_sign_out(5);
    CN323_data_in(22) <= VN1573_data_out(5);
    CN323_sign_in(22) <= VN1573_sign_out(5);
    CN323_data_in(23) <= VN1583_data_out(5);
    CN323_sign_in(23) <= VN1583_sign_out(5);
    CN323_data_in(24) <= VN1631_data_out(5);
    CN323_sign_in(24) <= VN1631_sign_out(5);
    CN323_data_in(25) <= VN1701_data_out(5);
    CN323_sign_in(25) <= VN1701_sign_out(5);
    CN323_data_in(26) <= VN1783_data_out(5);
    CN323_sign_in(26) <= VN1783_sign_out(5);
    CN323_data_in(27) <= VN1832_data_out(5);
    CN323_sign_in(27) <= VN1832_sign_out(5);
    CN323_data_in(28) <= VN1833_data_out(5);
    CN323_sign_in(28) <= VN1833_sign_out(5);
    CN323_data_in(29) <= VN1846_data_out(5);
    CN323_sign_in(29) <= VN1846_sign_out(5);
    CN323_data_in(30) <= VN1860_data_out(5);
    CN323_sign_in(30) <= VN1860_sign_out(5);
    CN323_data_in(31) <= VN1896_data_out(5);
    CN323_sign_in(31) <= VN1896_sign_out(5);
    CN324_data_in(0) <= VN49_data_out(5);
    CN324_sign_in(0) <= VN49_sign_out(5);
    CN324_data_in(1) <= VN109_data_out(5);
    CN324_sign_in(1) <= VN109_sign_out(5);
    CN324_data_in(2) <= VN113_data_out(5);
    CN324_sign_in(2) <= VN113_sign_out(5);
    CN324_data_in(3) <= VN223_data_out(5);
    CN324_sign_in(3) <= VN223_sign_out(5);
    CN324_data_in(4) <= VN273_data_out(5);
    CN324_sign_in(4) <= VN273_sign_out(5);
    CN324_data_in(5) <= VN302_data_out(5);
    CN324_sign_in(5) <= VN302_sign_out(5);
    CN324_data_in(6) <= VN369_data_out(5);
    CN324_sign_in(6) <= VN369_sign_out(5);
    CN324_data_in(7) <= VN400_data_out(5);
    CN324_sign_in(7) <= VN400_sign_out(5);
    CN324_data_in(8) <= VN490_data_out(5);
    CN324_sign_in(8) <= VN490_sign_out(5);
    CN324_data_in(9) <= VN544_data_out(5);
    CN324_sign_in(9) <= VN544_sign_out(5);
    CN324_data_in(10) <= VN593_data_out(5);
    CN324_sign_in(10) <= VN593_sign_out(5);
    CN324_data_in(11) <= VN640_data_out(5);
    CN324_sign_in(11) <= VN640_sign_out(5);
    CN324_data_in(12) <= VN693_data_out(5);
    CN324_sign_in(12) <= VN693_sign_out(5);
    CN324_data_in(13) <= VN821_data_out(5);
    CN324_sign_in(13) <= VN821_sign_out(5);
    CN324_data_in(14) <= VN855_data_out(5);
    CN324_sign_in(14) <= VN855_sign_out(5);
    CN324_data_in(15) <= VN936_data_out(5);
    CN324_sign_in(15) <= VN936_sign_out(5);
    CN324_data_in(16) <= VN951_data_out(5);
    CN324_sign_in(16) <= VN951_sign_out(5);
    CN324_data_in(17) <= VN1050_data_out(5);
    CN324_sign_in(17) <= VN1050_sign_out(5);
    CN324_data_in(18) <= VN1104_data_out(5);
    CN324_sign_in(18) <= VN1104_sign_out(5);
    CN324_data_in(19) <= VN1116_data_out(5);
    CN324_sign_in(19) <= VN1116_sign_out(5);
    CN324_data_in(20) <= VN1169_data_out(5);
    CN324_sign_in(20) <= VN1169_sign_out(5);
    CN324_data_in(21) <= VN1206_data_out(5);
    CN324_sign_in(21) <= VN1206_sign_out(5);
    CN324_data_in(22) <= VN1237_data_out(5);
    CN324_sign_in(22) <= VN1237_sign_out(5);
    CN324_data_in(23) <= VN1288_data_out(5);
    CN324_sign_in(23) <= VN1288_sign_out(5);
    CN324_data_in(24) <= VN1369_data_out(5);
    CN324_sign_in(24) <= VN1369_sign_out(5);
    CN324_data_in(25) <= VN1411_data_out(5);
    CN324_sign_in(25) <= VN1411_sign_out(5);
    CN324_data_in(26) <= VN1427_data_out(5);
    CN324_sign_in(26) <= VN1427_sign_out(5);
    CN324_data_in(27) <= VN1499_data_out(5);
    CN324_sign_in(27) <= VN1499_sign_out(5);
    CN324_data_in(28) <= VN1614_data_out(5);
    CN324_sign_in(28) <= VN1614_sign_out(5);
    CN324_data_in(29) <= VN1653_data_out(5);
    CN324_sign_in(29) <= VN1653_sign_out(5);
    CN324_data_in(30) <= VN1704_data_out(5);
    CN324_sign_in(30) <= VN1704_sign_out(5);
    CN324_data_in(31) <= VN1801_data_out(5);
    CN324_sign_in(31) <= VN1801_sign_out(5);
    CN325_data_in(0) <= VN48_data_out(5);
    CN325_sign_in(0) <= VN48_sign_out(5);
    CN325_data_in(1) <= VN70_data_out(5);
    CN325_sign_in(1) <= VN70_sign_out(5);
    CN325_data_in(2) <= VN137_data_out(5);
    CN325_sign_in(2) <= VN137_sign_out(5);
    CN325_data_in(3) <= VN185_data_out(5);
    CN325_sign_in(3) <= VN185_sign_out(5);
    CN325_data_in(4) <= VN242_data_out(5);
    CN325_sign_in(4) <= VN242_sign_out(5);
    CN325_data_in(5) <= VN284_data_out(5);
    CN325_sign_in(5) <= VN284_sign_out(5);
    CN325_data_in(6) <= VN382_data_out(5);
    CN325_sign_in(6) <= VN382_sign_out(5);
    CN325_data_in(7) <= VN395_data_out(5);
    CN325_sign_in(7) <= VN395_sign_out(5);
    CN325_data_in(8) <= VN476_data_out(5);
    CN325_sign_in(8) <= VN476_sign_out(5);
    CN325_data_in(9) <= VN518_data_out(5);
    CN325_sign_in(9) <= VN518_sign_out(5);
    CN325_data_in(10) <= VN583_data_out(5);
    CN325_sign_in(10) <= VN583_sign_out(5);
    CN325_data_in(11) <= VN653_data_out(5);
    CN325_sign_in(11) <= VN653_sign_out(5);
    CN325_data_in(12) <= VN704_data_out(5);
    CN325_sign_in(12) <= VN704_sign_out(5);
    CN325_data_in(13) <= VN753_data_out(5);
    CN325_sign_in(13) <= VN753_sign_out(5);
    CN325_data_in(14) <= VN784_data_out(5);
    CN325_sign_in(14) <= VN784_sign_out(5);
    CN325_data_in(15) <= VN832_data_out(5);
    CN325_sign_in(15) <= VN832_sign_out(5);
    CN325_data_in(16) <= VN940_data_out(5);
    CN325_sign_in(16) <= VN940_sign_out(5);
    CN325_data_in(17) <= VN979_data_out(5);
    CN325_sign_in(17) <= VN979_sign_out(5);
    CN325_data_in(18) <= VN1012_data_out(5);
    CN325_sign_in(18) <= VN1012_sign_out(5);
    CN325_data_in(19) <= VN1097_data_out(5);
    CN325_sign_in(19) <= VN1097_sign_out(5);
    CN325_data_in(20) <= VN1186_data_out(5);
    CN325_sign_in(20) <= VN1186_sign_out(5);
    CN325_data_in(21) <= VN1227_data_out(5);
    CN325_sign_in(21) <= VN1227_sign_out(5);
    CN325_data_in(22) <= VN1289_data_out(5);
    CN325_sign_in(22) <= VN1289_sign_out(5);
    CN325_data_in(23) <= VN1357_data_out(5);
    CN325_sign_in(23) <= VN1357_sign_out(5);
    CN325_data_in(24) <= VN1398_data_out(5);
    CN325_sign_in(24) <= VN1398_sign_out(5);
    CN325_data_in(25) <= VN1436_data_out(5);
    CN325_sign_in(25) <= VN1436_sign_out(5);
    CN325_data_in(26) <= VN1462_data_out(5);
    CN325_sign_in(26) <= VN1462_sign_out(5);
    CN325_data_in(27) <= VN1512_data_out(5);
    CN325_sign_in(27) <= VN1512_sign_out(5);
    CN325_data_in(28) <= VN1554_data_out(5);
    CN325_sign_in(28) <= VN1554_sign_out(5);
    CN325_data_in(29) <= VN1617_data_out(5);
    CN325_sign_in(29) <= VN1617_sign_out(5);
    CN325_data_in(30) <= VN1718_data_out(5);
    CN325_sign_in(30) <= VN1718_sign_out(5);
    CN325_data_in(31) <= VN1802_data_out(5);
    CN325_sign_in(31) <= VN1802_sign_out(5);
    CN326_data_in(0) <= VN47_data_out(5);
    CN326_sign_in(0) <= VN47_sign_out(5);
    CN326_data_in(1) <= VN62_data_out(5);
    CN326_sign_in(1) <= VN62_sign_out(5);
    CN326_data_in(2) <= VN203_data_out(5);
    CN326_sign_in(2) <= VN203_sign_out(5);
    CN326_data_in(3) <= VN241_data_out(5);
    CN326_sign_in(3) <= VN241_sign_out(5);
    CN326_data_in(4) <= VN304_data_out(5);
    CN326_sign_in(4) <= VN304_sign_out(5);
    CN326_data_in(5) <= VN527_data_out(5);
    CN326_sign_in(5) <= VN527_sign_out(5);
    CN326_data_in(6) <= VN606_data_out(5);
    CN326_sign_in(6) <= VN606_sign_out(5);
    CN326_data_in(7) <= VN663_data_out(5);
    CN326_sign_in(7) <= VN663_sign_out(5);
    CN326_data_in(8) <= VN697_data_out(5);
    CN326_sign_in(8) <= VN697_sign_out(5);
    CN326_data_in(9) <= VN722_data_out(5);
    CN326_sign_in(9) <= VN722_sign_out(5);
    CN326_data_in(10) <= VN748_data_out(5);
    CN326_sign_in(10) <= VN748_sign_out(5);
    CN326_data_in(11) <= VN788_data_out(5);
    CN326_sign_in(11) <= VN788_sign_out(5);
    CN326_data_in(12) <= VN867_data_out(5);
    CN326_sign_in(12) <= VN867_sign_out(5);
    CN326_data_in(13) <= VN969_data_out(5);
    CN326_sign_in(13) <= VN969_sign_out(5);
    CN326_data_in(14) <= VN1041_data_out(5);
    CN326_sign_in(14) <= VN1041_sign_out(5);
    CN326_data_in(15) <= VN1061_data_out(5);
    CN326_sign_in(15) <= VN1061_sign_out(5);
    CN326_data_in(16) <= VN1140_data_out(5);
    CN326_sign_in(16) <= VN1140_sign_out(5);
    CN326_data_in(17) <= VN1170_data_out(5);
    CN326_sign_in(17) <= VN1170_sign_out(5);
    CN326_data_in(18) <= VN1261_data_out(5);
    CN326_sign_in(18) <= VN1261_sign_out(5);
    CN326_data_in(19) <= VN1318_data_out(5);
    CN326_sign_in(19) <= VN1318_sign_out(5);
    CN326_data_in(20) <= VN1374_data_out(5);
    CN326_sign_in(20) <= VN1374_sign_out(5);
    CN326_data_in(21) <= VN1485_data_out(5);
    CN326_sign_in(21) <= VN1485_sign_out(5);
    CN326_data_in(22) <= VN1548_data_out(5);
    CN326_sign_in(22) <= VN1548_sign_out(5);
    CN326_data_in(23) <= VN1569_data_out(5);
    CN326_sign_in(23) <= VN1569_sign_out(5);
    CN326_data_in(24) <= VN1671_data_out(5);
    CN326_sign_in(24) <= VN1671_sign_out(5);
    CN326_data_in(25) <= VN1764_data_out(5);
    CN326_sign_in(25) <= VN1764_sign_out(5);
    CN326_data_in(26) <= VN1827_data_out(5);
    CN326_sign_in(26) <= VN1827_sign_out(5);
    CN326_data_in(27) <= VN1909_data_out(5);
    CN326_sign_in(27) <= VN1909_sign_out(5);
    CN326_data_in(28) <= VN1922_data_out(5);
    CN326_sign_in(28) <= VN1922_sign_out(5);
    CN326_data_in(29) <= VN1926_data_out(5);
    CN326_sign_in(29) <= VN1926_sign_out(5);
    CN326_data_in(30) <= VN1972_data_out(5);
    CN326_sign_in(30) <= VN1972_sign_out(5);
    CN326_data_in(31) <= VN1981_data_out(5);
    CN326_sign_in(31) <= VN1981_sign_out(5);
    CN327_data_in(0) <= VN46_data_out(5);
    CN327_sign_in(0) <= VN46_sign_out(5);
    CN327_data_in(1) <= VN94_data_out(5);
    CN327_sign_in(1) <= VN94_sign_out(5);
    CN327_data_in(2) <= VN148_data_out(5);
    CN327_sign_in(2) <= VN148_sign_out(5);
    CN327_data_in(3) <= VN211_data_out(5);
    CN327_sign_in(3) <= VN211_sign_out(5);
    CN327_data_in(4) <= VN272_data_out(5);
    CN327_sign_in(4) <= VN272_sign_out(5);
    CN327_data_in(5) <= VN318_data_out(5);
    CN327_sign_in(5) <= VN318_sign_out(5);
    CN327_data_in(6) <= VN361_data_out(5);
    CN327_sign_in(6) <= VN361_sign_out(5);
    CN327_data_in(7) <= VN446_data_out(5);
    CN327_sign_in(7) <= VN446_sign_out(5);
    CN327_data_in(8) <= VN502_data_out(5);
    CN327_sign_in(8) <= VN502_sign_out(5);
    CN327_data_in(9) <= VN521_data_out(5);
    CN327_sign_in(9) <= VN521_sign_out(5);
    CN327_data_in(10) <= VN612_data_out(5);
    CN327_sign_in(10) <= VN612_sign_out(5);
    CN327_data_in(11) <= VN634_data_out(5);
    CN327_sign_in(11) <= VN634_sign_out(5);
    CN327_data_in(12) <= VN701_data_out(5);
    CN327_sign_in(12) <= VN701_sign_out(5);
    CN327_data_in(13) <= VN777_data_out(5);
    CN327_sign_in(13) <= VN777_sign_out(5);
    CN327_data_in(14) <= VN870_data_out(5);
    CN327_sign_in(14) <= VN870_sign_out(5);
    CN327_data_in(15) <= VN911_data_out(5);
    CN327_sign_in(15) <= VN911_sign_out(5);
    CN327_data_in(16) <= VN956_data_out(5);
    CN327_sign_in(16) <= VN956_sign_out(5);
    CN327_data_in(17) <= VN1038_data_out(5);
    CN327_sign_in(17) <= VN1038_sign_out(5);
    CN327_data_in(18) <= VN1066_data_out(5);
    CN327_sign_in(18) <= VN1066_sign_out(5);
    CN327_data_in(19) <= VN1151_data_out(5);
    CN327_sign_in(19) <= VN1151_sign_out(5);
    CN327_data_in(20) <= VN1182_data_out(5);
    CN327_sign_in(20) <= VN1182_sign_out(5);
    CN327_data_in(21) <= VN1244_data_out(5);
    CN327_sign_in(21) <= VN1244_sign_out(5);
    CN327_data_in(22) <= VN1310_data_out(5);
    CN327_sign_in(22) <= VN1310_sign_out(5);
    CN327_data_in(23) <= VN1349_data_out(5);
    CN327_sign_in(23) <= VN1349_sign_out(5);
    CN327_data_in(24) <= VN1401_data_out(5);
    CN327_sign_in(24) <= VN1401_sign_out(5);
    CN327_data_in(25) <= VN1456_data_out(5);
    CN327_sign_in(25) <= VN1456_sign_out(5);
    CN327_data_in(26) <= VN1479_data_out(5);
    CN327_sign_in(26) <= VN1479_sign_out(5);
    CN327_data_in(27) <= VN1500_data_out(5);
    CN327_sign_in(27) <= VN1500_sign_out(5);
    CN327_data_in(28) <= VN1632_data_out(5);
    CN327_sign_in(28) <= VN1632_sign_out(5);
    CN327_data_in(29) <= VN1699_data_out(5);
    CN327_sign_in(29) <= VN1699_sign_out(5);
    CN327_data_in(30) <= VN1730_data_out(5);
    CN327_sign_in(30) <= VN1730_sign_out(5);
    CN327_data_in(31) <= VN1873_data_out(5);
    CN327_sign_in(31) <= VN1873_sign_out(5);
    CN328_data_in(0) <= VN45_data_out(5);
    CN328_sign_in(0) <= VN45_sign_out(5);
    CN328_data_in(1) <= VN103_data_out(5);
    CN328_sign_in(1) <= VN103_sign_out(5);
    CN328_data_in(2) <= VN168_data_out(5);
    CN328_sign_in(2) <= VN168_sign_out(5);
    CN328_data_in(3) <= VN314_data_out(5);
    CN328_sign_in(3) <= VN314_sign_out(5);
    CN328_data_in(4) <= VN377_data_out(5);
    CN328_sign_in(4) <= VN377_sign_out(5);
    CN328_data_in(5) <= VN413_data_out(5);
    CN328_sign_in(5) <= VN413_sign_out(5);
    CN328_data_in(6) <= VN483_data_out(5);
    CN328_sign_in(6) <= VN483_sign_out(5);
    CN328_data_in(7) <= VN524_data_out(5);
    CN328_sign_in(7) <= VN524_sign_out(5);
    CN328_data_in(8) <= VN597_data_out(5);
    CN328_sign_in(8) <= VN597_sign_out(5);
    CN328_data_in(9) <= VN690_data_out(5);
    CN328_sign_in(9) <= VN690_sign_out(5);
    CN328_data_in(10) <= VN737_data_out(5);
    CN328_sign_in(10) <= VN737_sign_out(5);
    CN328_data_in(11) <= VN787_data_out(5);
    CN328_sign_in(11) <= VN787_sign_out(5);
    CN328_data_in(12) <= VN857_data_out(5);
    CN328_sign_in(12) <= VN857_sign_out(5);
    CN328_data_in(13) <= VN893_data_out(5);
    CN328_sign_in(13) <= VN893_sign_out(5);
    CN328_data_in(14) <= VN975_data_out(5);
    CN328_sign_in(14) <= VN975_sign_out(5);
    CN328_data_in(15) <= VN1055_data_out(5);
    CN328_sign_in(15) <= VN1055_sign_out(5);
    CN328_data_in(16) <= VN1144_data_out(5);
    CN328_sign_in(16) <= VN1144_sign_out(5);
    CN328_data_in(17) <= VN1328_data_out(5);
    CN328_sign_in(17) <= VN1328_sign_out(5);
    CN328_data_in(18) <= VN1346_data_out(5);
    CN328_sign_in(18) <= VN1346_sign_out(5);
    CN328_data_in(19) <= VN1421_data_out(5);
    CN328_sign_in(19) <= VN1421_sign_out(5);
    CN328_data_in(20) <= VN1439_data_out(5);
    CN328_sign_in(20) <= VN1439_sign_out(5);
    CN328_data_in(21) <= VN1486_data_out(5);
    CN328_sign_in(21) <= VN1486_sign_out(5);
    CN328_data_in(22) <= VN1491_data_out(5);
    CN328_sign_in(22) <= VN1491_sign_out(5);
    CN328_data_in(23) <= VN1509_data_out(5);
    CN328_sign_in(23) <= VN1509_sign_out(5);
    CN328_data_in(24) <= VN1672_data_out(5);
    CN328_sign_in(24) <= VN1672_sign_out(5);
    CN328_data_in(25) <= VN1688_data_out(5);
    CN328_sign_in(25) <= VN1688_sign_out(5);
    CN328_data_in(26) <= VN1742_data_out(5);
    CN328_sign_in(26) <= VN1742_sign_out(5);
    CN328_data_in(27) <= VN1796_data_out(5);
    CN328_sign_in(27) <= VN1796_sign_out(5);
    CN328_data_in(28) <= VN1814_data_out(5);
    CN328_sign_in(28) <= VN1814_sign_out(5);
    CN328_data_in(29) <= VN1936_data_out(5);
    CN328_sign_in(29) <= VN1936_sign_out(5);
    CN328_data_in(30) <= VN1946_data_out(5);
    CN328_sign_in(30) <= VN1946_sign_out(5);
    CN328_data_in(31) <= VN1957_data_out(5);
    CN328_sign_in(31) <= VN1957_sign_out(5);
    CN329_data_in(0) <= VN44_data_out(5);
    CN329_sign_in(0) <= VN44_sign_out(5);
    CN329_data_in(1) <= VN97_data_out(5);
    CN329_sign_in(1) <= VN97_sign_out(5);
    CN329_data_in(2) <= VN131_data_out(5);
    CN329_sign_in(2) <= VN131_sign_out(5);
    CN329_data_in(3) <= VN212_data_out(5);
    CN329_sign_in(3) <= VN212_sign_out(5);
    CN329_data_in(4) <= VN255_data_out(5);
    CN329_sign_in(4) <= VN255_sign_out(5);
    CN329_data_in(5) <= VN280_data_out(5);
    CN329_sign_in(5) <= VN280_sign_out(5);
    CN329_data_in(6) <= VN348_data_out(5);
    CN329_sign_in(6) <= VN348_sign_out(5);
    CN329_data_in(7) <= VN420_data_out(5);
    CN329_sign_in(7) <= VN420_sign_out(5);
    CN329_data_in(8) <= VN494_data_out(5);
    CN329_sign_in(8) <= VN494_sign_out(5);
    CN329_data_in(9) <= VN516_data_out(5);
    CN329_sign_in(9) <= VN516_sign_out(5);
    CN329_data_in(10) <= VN599_data_out(5);
    CN329_sign_in(10) <= VN599_sign_out(5);
    CN329_data_in(11) <= VN665_data_out(5);
    CN329_sign_in(11) <= VN665_sign_out(5);
    CN329_data_in(12) <= VN671_data_out(5);
    CN329_sign_in(12) <= VN671_sign_out(5);
    CN329_data_in(13) <= VN760_data_out(5);
    CN329_sign_in(13) <= VN760_sign_out(5);
    CN329_data_in(14) <= VN782_data_out(5);
    CN329_sign_in(14) <= VN782_sign_out(5);
    CN329_data_in(15) <= VN833_data_out(5);
    CN329_sign_in(15) <= VN833_sign_out(5);
    CN329_data_in(16) <= VN907_data_out(5);
    CN329_sign_in(16) <= VN907_sign_out(5);
    CN329_data_in(17) <= VN947_data_out(5);
    CN329_sign_in(17) <= VN947_sign_out(5);
    CN329_data_in(18) <= VN1047_data_out(5);
    CN329_sign_in(18) <= VN1047_sign_out(5);
    CN329_data_in(19) <= VN1065_data_out(5);
    CN329_sign_in(19) <= VN1065_sign_out(5);
    CN329_data_in(20) <= VN1148_data_out(5);
    CN329_sign_in(20) <= VN1148_sign_out(5);
    CN329_data_in(21) <= VN1268_data_out(5);
    CN329_sign_in(21) <= VN1268_sign_out(5);
    CN329_data_in(22) <= VN1278_data_out(5);
    CN329_sign_in(22) <= VN1278_sign_out(5);
    CN329_data_in(23) <= VN1361_data_out(5);
    CN329_sign_in(23) <= VN1361_sign_out(5);
    CN329_data_in(24) <= VN1515_data_out(5);
    CN329_sign_in(24) <= VN1515_sign_out(5);
    CN329_data_in(25) <= VN1530_data_out(5);
    CN329_sign_in(25) <= VN1530_sign_out(5);
    CN329_data_in(26) <= VN1538_data_out(5);
    CN329_sign_in(26) <= VN1538_sign_out(5);
    CN329_data_in(27) <= VN1560_data_out(5);
    CN329_sign_in(27) <= VN1560_sign_out(5);
    CN329_data_in(28) <= VN1607_data_out(5);
    CN329_sign_in(28) <= VN1607_sign_out(5);
    CN329_data_in(29) <= VN1626_data_out(5);
    CN329_sign_in(29) <= VN1626_sign_out(5);
    CN329_data_in(30) <= VN1667_data_out(5);
    CN329_sign_in(30) <= VN1667_sign_out(5);
    CN329_data_in(31) <= VN1803_data_out(5);
    CN329_sign_in(31) <= VN1803_sign_out(5);
    CN330_data_in(0) <= VN43_data_out(5);
    CN330_sign_in(0) <= VN43_sign_out(5);
    CN330_data_in(1) <= VN101_data_out(5);
    CN330_sign_in(1) <= VN101_sign_out(5);
    CN330_data_in(2) <= VN132_data_out(5);
    CN330_sign_in(2) <= VN132_sign_out(5);
    CN330_data_in(3) <= VN202_data_out(5);
    CN330_sign_in(3) <= VN202_sign_out(5);
    CN330_data_in(4) <= VN243_data_out(5);
    CN330_sign_in(4) <= VN243_sign_out(5);
    CN330_data_in(5) <= VN385_data_out(5);
    CN330_sign_in(5) <= VN385_sign_out(5);
    CN330_data_in(6) <= VN404_data_out(5);
    CN330_sign_in(6) <= VN404_sign_out(5);
    CN330_data_in(7) <= VN503_data_out(5);
    CN330_sign_in(7) <= VN503_sign_out(5);
    CN330_data_in(8) <= VN553_data_out(5);
    CN330_sign_in(8) <= VN553_sign_out(5);
    CN330_data_in(9) <= VN569_data_out(5);
    CN330_sign_in(9) <= VN569_sign_out(5);
    CN330_data_in(10) <= VN626_data_out(5);
    CN330_sign_in(10) <= VN626_sign_out(5);
    CN330_data_in(11) <= VN710_data_out(5);
    CN330_sign_in(11) <= VN710_sign_out(5);
    CN330_data_in(12) <= VN758_data_out(5);
    CN330_sign_in(12) <= VN758_sign_out(5);
    CN330_data_in(13) <= VN819_data_out(5);
    CN330_sign_in(13) <= VN819_sign_out(5);
    CN330_data_in(14) <= VN917_data_out(5);
    CN330_sign_in(14) <= VN917_sign_out(5);
    CN330_data_in(15) <= VN944_data_out(5);
    CN330_sign_in(15) <= VN944_sign_out(5);
    CN330_data_in(16) <= VN1022_data_out(5);
    CN330_sign_in(16) <= VN1022_sign_out(5);
    CN330_data_in(17) <= VN1138_data_out(5);
    CN330_sign_in(17) <= VN1138_sign_out(5);
    CN330_data_in(18) <= VN1208_data_out(5);
    CN330_sign_in(18) <= VN1208_sign_out(5);
    CN330_data_in(19) <= VN1240_data_out(5);
    CN330_sign_in(19) <= VN1240_sign_out(5);
    CN330_data_in(20) <= VN1384_data_out(5);
    CN330_sign_in(20) <= VN1384_sign_out(5);
    CN330_data_in(21) <= VN1425_data_out(5);
    CN330_sign_in(21) <= VN1425_sign_out(5);
    CN330_data_in(22) <= VN1483_data_out(5);
    CN330_sign_in(22) <= VN1483_sign_out(5);
    CN330_data_in(23) <= VN1508_data_out(5);
    CN330_sign_in(23) <= VN1508_sign_out(5);
    CN330_data_in(24) <= VN1532_data_out(5);
    CN330_sign_in(24) <= VN1532_sign_out(5);
    CN330_data_in(25) <= VN1684_data_out(5);
    CN330_sign_in(25) <= VN1684_sign_out(5);
    CN330_data_in(26) <= VN1747_data_out(5);
    CN330_sign_in(26) <= VN1747_sign_out(5);
    CN330_data_in(27) <= VN1795_data_out(5);
    CN330_sign_in(27) <= VN1795_sign_out(5);
    CN330_data_in(28) <= VN1823_data_out(5);
    CN330_sign_in(28) <= VN1823_sign_out(5);
    CN330_data_in(29) <= VN1865_data_out(5);
    CN330_sign_in(29) <= VN1865_sign_out(5);
    CN330_data_in(30) <= VN1867_data_out(5);
    CN330_sign_in(30) <= VN1867_sign_out(5);
    CN330_data_in(31) <= VN1897_data_out(5);
    CN330_sign_in(31) <= VN1897_sign_out(5);
    CN331_data_in(0) <= VN42_data_out(5);
    CN331_sign_in(0) <= VN42_sign_out(5);
    CN331_data_in(1) <= VN92_data_out(5);
    CN331_sign_in(1) <= VN92_sign_out(5);
    CN331_data_in(2) <= VN167_data_out(5);
    CN331_sign_in(2) <= VN167_sign_out(5);
    CN331_data_in(3) <= VN172_data_out(5);
    CN331_sign_in(3) <= VN172_sign_out(5);
    CN331_data_in(4) <= VN350_data_out(5);
    CN331_sign_in(4) <= VN350_sign_out(5);
    CN331_data_in(5) <= VN406_data_out(5);
    CN331_sign_in(5) <= VN406_sign_out(5);
    CN331_data_in(6) <= VN534_data_out(5);
    CN331_sign_in(6) <= VN534_sign_out(5);
    CN331_data_in(7) <= VN604_data_out(5);
    CN331_sign_in(7) <= VN604_sign_out(5);
    CN331_data_in(8) <= VN646_data_out(5);
    CN331_sign_in(8) <= VN646_sign_out(5);
    CN331_data_in(9) <= VN720_data_out(5);
    CN331_sign_in(9) <= VN720_sign_out(5);
    CN331_data_in(10) <= VN736_data_out(5);
    CN331_sign_in(10) <= VN736_sign_out(5);
    CN331_data_in(11) <= VN826_data_out(5);
    CN331_sign_in(11) <= VN826_sign_out(5);
    CN331_data_in(12) <= VN879_data_out(5);
    CN331_sign_in(12) <= VN879_sign_out(5);
    CN331_data_in(13) <= VN943_data_out(5);
    CN331_sign_in(13) <= VN943_sign_out(5);
    CN331_data_in(14) <= VN961_data_out(5);
    CN331_sign_in(14) <= VN961_sign_out(5);
    CN331_data_in(15) <= VN1031_data_out(5);
    CN331_sign_in(15) <= VN1031_sign_out(5);
    CN331_data_in(16) <= VN1117_data_out(5);
    CN331_sign_in(16) <= VN1117_sign_out(5);
    CN331_data_in(17) <= VN1194_data_out(5);
    CN331_sign_in(17) <= VN1194_sign_out(5);
    CN331_data_in(18) <= VN1229_data_out(5);
    CN331_sign_in(18) <= VN1229_sign_out(5);
    CN331_data_in(19) <= VN1428_data_out(5);
    CN331_sign_in(19) <= VN1428_sign_out(5);
    CN331_data_in(20) <= VN1449_data_out(5);
    CN331_sign_in(20) <= VN1449_sign_out(5);
    CN331_data_in(21) <= VN1477_data_out(5);
    CN331_sign_in(21) <= VN1477_sign_out(5);
    CN331_data_in(22) <= VN1529_data_out(5);
    CN331_sign_in(22) <= VN1529_sign_out(5);
    CN331_data_in(23) <= VN1533_data_out(5);
    CN331_sign_in(23) <= VN1533_sign_out(5);
    CN331_data_in(24) <= VN1634_data_out(5);
    CN331_sign_in(24) <= VN1634_sign_out(5);
    CN331_data_in(25) <= VN1650_data_out(5);
    CN331_sign_in(25) <= VN1650_sign_out(5);
    CN331_data_in(26) <= VN1706_data_out(5);
    CN331_sign_in(26) <= VN1706_sign_out(5);
    CN331_data_in(27) <= VN1753_data_out(5);
    CN331_sign_in(27) <= VN1753_sign_out(5);
    CN331_data_in(28) <= VN1862_data_out(5);
    CN331_sign_in(28) <= VN1862_sign_out(5);
    CN331_data_in(29) <= VN1963_data_out(5);
    CN331_sign_in(29) <= VN1963_sign_out(5);
    CN331_data_in(30) <= VN1991_data_out(5);
    CN331_sign_in(30) <= VN1991_sign_out(5);
    CN331_data_in(31) <= VN1993_data_out(5);
    CN331_sign_in(31) <= VN1993_sign_out(5);
    CN332_data_in(0) <= VN41_data_out(5);
    CN332_sign_in(0) <= VN41_sign_out(5);
    CN332_data_in(1) <= VN71_data_out(5);
    CN332_sign_in(1) <= VN71_sign_out(5);
    CN332_data_in(2) <= VN158_data_out(5);
    CN332_sign_in(2) <= VN158_sign_out(5);
    CN332_data_in(3) <= VN179_data_out(5);
    CN332_sign_in(3) <= VN179_sign_out(5);
    CN332_data_in(4) <= VN240_data_out(5);
    CN332_sign_in(4) <= VN240_sign_out(5);
    CN332_data_in(5) <= VN363_data_out(5);
    CN332_sign_in(5) <= VN363_sign_out(5);
    CN332_data_in(6) <= VN431_data_out(5);
    CN332_sign_in(6) <= VN431_sign_out(5);
    CN332_data_in(7) <= VN489_data_out(5);
    CN332_sign_in(7) <= VN489_sign_out(5);
    CN332_data_in(8) <= VN548_data_out(5);
    CN332_sign_in(8) <= VN548_sign_out(5);
    CN332_data_in(9) <= VN561_data_out(5);
    CN332_sign_in(9) <= VN561_sign_out(5);
    CN332_data_in(10) <= VN772_data_out(5);
    CN332_sign_in(10) <= VN772_sign_out(5);
    CN332_data_in(11) <= VN793_data_out(5);
    CN332_sign_in(11) <= VN793_sign_out(5);
    CN332_data_in(12) <= VN865_data_out(5);
    CN332_sign_in(12) <= VN865_sign_out(5);
    CN332_data_in(13) <= VN931_data_out(5);
    CN332_sign_in(13) <= VN931_sign_out(5);
    CN332_data_in(14) <= VN953_data_out(5);
    CN332_sign_in(14) <= VN953_sign_out(5);
    CN332_data_in(15) <= VN1025_data_out(5);
    CN332_sign_in(15) <= VN1025_sign_out(5);
    CN332_data_in(16) <= VN1157_data_out(5);
    CN332_sign_in(16) <= VN1157_sign_out(5);
    CN332_data_in(17) <= VN1211_data_out(5);
    CN332_sign_in(17) <= VN1211_sign_out(5);
    CN332_data_in(18) <= VN1271_data_out(5);
    CN332_sign_in(18) <= VN1271_sign_out(5);
    CN332_data_in(19) <= VN1326_data_out(5);
    CN332_sign_in(19) <= VN1326_sign_out(5);
    CN332_data_in(20) <= VN1338_data_out(5);
    CN332_sign_in(20) <= VN1338_sign_out(5);
    CN332_data_in(21) <= VN1389_data_out(5);
    CN332_sign_in(21) <= VN1389_sign_out(5);
    CN332_data_in(22) <= VN1420_data_out(5);
    CN332_sign_in(22) <= VN1420_sign_out(5);
    CN332_data_in(23) <= VN1600_data_out(5);
    CN332_sign_in(23) <= VN1600_sign_out(5);
    CN332_data_in(24) <= VN1627_data_out(5);
    CN332_sign_in(24) <= VN1627_sign_out(5);
    CN332_data_in(25) <= VN1676_data_out(5);
    CN332_sign_in(25) <= VN1676_sign_out(5);
    CN332_data_in(26) <= VN1724_data_out(5);
    CN332_sign_in(26) <= VN1724_sign_out(5);
    CN332_data_in(27) <= VN1782_data_out(5);
    CN332_sign_in(27) <= VN1782_sign_out(5);
    CN332_data_in(28) <= VN1885_data_out(5);
    CN332_sign_in(28) <= VN1885_sign_out(5);
    CN332_data_in(29) <= VN1925_data_out(5);
    CN332_sign_in(29) <= VN1925_sign_out(5);
    CN332_data_in(30) <= VN2022_data_out(5);
    CN332_sign_in(30) <= VN2022_sign_out(5);
    CN332_data_in(31) <= VN2029_data_out(5);
    CN332_sign_in(31) <= VN2029_sign_out(5);
    CN333_data_in(0) <= VN108_data_out(5);
    CN333_sign_in(0) <= VN108_sign_out(5);
    CN333_data_in(1) <= VN117_data_out(5);
    CN333_sign_in(1) <= VN117_sign_out(5);
    CN333_data_in(2) <= VN215_data_out(5);
    CN333_sign_in(2) <= VN215_sign_out(5);
    CN333_data_in(3) <= VN265_data_out(5);
    CN333_sign_in(3) <= VN265_sign_out(5);
    CN333_data_in(4) <= VN324_data_out(5);
    CN333_sign_in(4) <= VN324_sign_out(5);
    CN333_data_in(5) <= VN359_data_out(5);
    CN333_sign_in(5) <= VN359_sign_out(5);
    CN333_data_in(6) <= VN411_data_out(5);
    CN333_sign_in(6) <= VN411_sign_out(5);
    CN333_data_in(7) <= VN651_data_out(5);
    CN333_sign_in(7) <= VN651_sign_out(5);
    CN333_data_in(8) <= VN774_data_out(5);
    CN333_sign_in(8) <= VN774_sign_out(5);
    CN333_data_in(9) <= VN835_data_out(5);
    CN333_sign_in(9) <= VN835_sign_out(5);
    CN333_data_in(10) <= VN920_data_out(5);
    CN333_sign_in(10) <= VN920_sign_out(5);
    CN333_data_in(11) <= VN986_data_out(5);
    CN333_sign_in(11) <= VN986_sign_out(5);
    CN333_data_in(12) <= VN1071_data_out(5);
    CN333_sign_in(12) <= VN1071_sign_out(5);
    CN333_data_in(13) <= VN1175_data_out(5);
    CN333_sign_in(13) <= VN1175_sign_out(5);
    CN333_data_in(14) <= VN1232_data_out(5);
    CN333_sign_in(14) <= VN1232_sign_out(5);
    CN333_data_in(15) <= VN1308_data_out(5);
    CN333_sign_in(15) <= VN1308_sign_out(5);
    CN333_data_in(16) <= VN1429_data_out(5);
    CN333_sign_in(16) <= VN1429_sign_out(5);
    CN333_data_in(17) <= VN1448_data_out(5);
    CN333_sign_in(17) <= VN1448_sign_out(5);
    CN333_data_in(18) <= VN1458_data_out(5);
    CN333_sign_in(18) <= VN1458_sign_out(5);
    CN333_data_in(19) <= VN1551_data_out(5);
    CN333_sign_in(19) <= VN1551_sign_out(5);
    CN333_data_in(20) <= VN1615_data_out(5);
    CN333_sign_in(20) <= VN1615_sign_out(5);
    CN333_data_in(21) <= VN1726_data_out(5);
    CN333_sign_in(21) <= VN1726_sign_out(5);
    CN333_data_in(22) <= VN1776_data_out(5);
    CN333_sign_in(22) <= VN1776_sign_out(5);
    CN333_data_in(23) <= VN1810_data_out(5);
    CN333_sign_in(23) <= VN1810_sign_out(5);
    CN333_data_in(24) <= VN1820_data_out(5);
    CN333_sign_in(24) <= VN1820_sign_out(5);
    CN333_data_in(25) <= VN1888_data_out(5);
    CN333_sign_in(25) <= VN1888_sign_out(5);
    CN333_data_in(26) <= VN1961_data_out(5);
    CN333_sign_in(26) <= VN1961_sign_out(5);
    CN333_data_in(27) <= VN1980_data_out(5);
    CN333_sign_in(27) <= VN1980_sign_out(5);
    CN333_data_in(28) <= VN2018_data_out(5);
    CN333_sign_in(28) <= VN2018_sign_out(5);
    CN333_data_in(29) <= VN2019_data_out(5);
    CN333_sign_in(29) <= VN2019_sign_out(5);
    CN333_data_in(30) <= VN2020_data_out(5);
    CN333_sign_in(30) <= VN2020_sign_out(5);
    CN333_data_in(31) <= VN2034_data_out(5);
    CN333_sign_in(31) <= VN2034_sign_out(5);
    CN334_data_in(0) <= VN40_data_out(5);
    CN334_sign_in(0) <= VN40_sign_out(5);
    CN334_data_in(1) <= VN66_data_out(5);
    CN334_sign_in(1) <= VN66_sign_out(5);
    CN334_data_in(2) <= VN217_data_out(5);
    CN334_sign_in(2) <= VN217_sign_out(5);
    CN334_data_in(3) <= VN286_data_out(5);
    CN334_sign_in(3) <= VN286_sign_out(5);
    CN334_data_in(4) <= VN380_data_out(5);
    CN334_sign_in(4) <= VN380_sign_out(5);
    CN334_data_in(5) <= VN497_data_out(5);
    CN334_sign_in(5) <= VN497_sign_out(5);
    CN334_data_in(6) <= VN528_data_out(5);
    CN334_sign_in(6) <= VN528_sign_out(5);
    CN334_data_in(7) <= VN598_data_out(5);
    CN334_sign_in(7) <= VN598_sign_out(5);
    CN334_data_in(8) <= VN654_data_out(5);
    CN334_sign_in(8) <= VN654_sign_out(5);
    CN334_data_in(9) <= VN692_data_out(5);
    CN334_sign_in(9) <= VN692_sign_out(5);
    CN334_data_in(10) <= VN761_data_out(5);
    CN334_sign_in(10) <= VN761_sign_out(5);
    CN334_data_in(11) <= VN824_data_out(5);
    CN334_sign_in(11) <= VN824_sign_out(5);
    CN334_data_in(12) <= VN881_data_out(5);
    CN334_sign_in(12) <= VN881_sign_out(5);
    CN334_data_in(13) <= VN934_data_out(5);
    CN334_sign_in(13) <= VN934_sign_out(5);
    CN334_data_in(14) <= VN996_data_out(5);
    CN334_sign_in(14) <= VN996_sign_out(5);
    CN334_data_in(15) <= VN1020_data_out(5);
    CN334_sign_in(15) <= VN1020_sign_out(5);
    CN334_data_in(16) <= VN1069_data_out(5);
    CN334_sign_in(16) <= VN1069_sign_out(5);
    CN334_data_in(17) <= VN1123_data_out(5);
    CN334_sign_in(17) <= VN1123_sign_out(5);
    CN334_data_in(18) <= VN1184_data_out(5);
    CN334_sign_in(18) <= VN1184_sign_out(5);
    CN334_data_in(19) <= VN1250_data_out(5);
    CN334_sign_in(19) <= VN1250_sign_out(5);
    CN334_data_in(20) <= VN1314_data_out(5);
    CN334_sign_in(20) <= VN1314_sign_out(5);
    CN334_data_in(21) <= VN1336_data_out(5);
    CN334_sign_in(21) <= VN1336_sign_out(5);
    CN334_data_in(22) <= VN1394_data_out(5);
    CN334_sign_in(22) <= VN1394_sign_out(5);
    CN334_data_in(23) <= VN1443_data_out(5);
    CN334_sign_in(23) <= VN1443_sign_out(5);
    CN334_data_in(24) <= VN1630_data_out(5);
    CN334_sign_in(24) <= VN1630_sign_out(5);
    CN334_data_in(25) <= VN1712_data_out(5);
    CN334_sign_in(25) <= VN1712_sign_out(5);
    CN334_data_in(26) <= VN1755_data_out(5);
    CN334_sign_in(26) <= VN1755_sign_out(5);
    CN334_data_in(27) <= VN1852_data_out(5);
    CN334_sign_in(27) <= VN1852_sign_out(5);
    CN334_data_in(28) <= VN1913_data_out(5);
    CN334_sign_in(28) <= VN1913_sign_out(5);
    CN334_data_in(29) <= VN1997_data_out(5);
    CN334_sign_in(29) <= VN1997_sign_out(5);
    CN334_data_in(30) <= VN2021_data_out(5);
    CN334_sign_in(30) <= VN2021_sign_out(5);
    CN334_data_in(31) <= VN2026_data_out(5);
    CN334_sign_in(31) <= VN2026_sign_out(5);
    CN335_data_in(0) <= VN39_data_out(5);
    CN335_sign_in(0) <= VN39_sign_out(5);
    CN335_data_in(1) <= VN78_data_out(5);
    CN335_sign_in(1) <= VN78_sign_out(5);
    CN335_data_in(2) <= VN170_data_out(5);
    CN335_sign_in(2) <= VN170_sign_out(5);
    CN335_data_in(3) <= VN189_data_out(5);
    CN335_sign_in(3) <= VN189_sign_out(5);
    CN335_data_in(4) <= VN274_data_out(5);
    CN335_sign_in(4) <= VN274_sign_out(5);
    CN335_data_in(5) <= VN291_data_out(5);
    CN335_sign_in(5) <= VN291_sign_out(5);
    CN335_data_in(6) <= VN343_data_out(5);
    CN335_sign_in(6) <= VN343_sign_out(5);
    CN335_data_in(7) <= VN432_data_out(5);
    CN335_sign_in(7) <= VN432_sign_out(5);
    CN335_data_in(8) <= VN465_data_out(5);
    CN335_sign_in(8) <= VN465_sign_out(5);
    CN335_data_in(9) <= VN517_data_out(5);
    CN335_sign_in(9) <= VN517_sign_out(5);
    CN335_data_in(10) <= VN611_data_out(5);
    CN335_sign_in(10) <= VN611_sign_out(5);
    CN335_data_in(11) <= VN645_data_out(5);
    CN335_sign_in(11) <= VN645_sign_out(5);
    CN335_data_in(12) <= VN679_data_out(5);
    CN335_sign_in(12) <= VN679_sign_out(5);
    CN335_data_in(13) <= VN804_data_out(5);
    CN335_sign_in(13) <= VN804_sign_out(5);
    CN335_data_in(14) <= VN868_data_out(5);
    CN335_sign_in(14) <= VN868_sign_out(5);
    CN335_data_in(15) <= VN899_data_out(5);
    CN335_sign_in(15) <= VN899_sign_out(5);
    CN335_data_in(16) <= VN990_data_out(5);
    CN335_sign_in(16) <= VN990_sign_out(5);
    CN335_data_in(17) <= VN1056_data_out(5);
    CN335_sign_in(17) <= VN1056_sign_out(5);
    CN335_data_in(18) <= VN1099_data_out(5);
    CN335_sign_in(18) <= VN1099_sign_out(5);
    CN335_data_in(19) <= VN1152_data_out(5);
    CN335_sign_in(19) <= VN1152_sign_out(5);
    CN335_data_in(20) <= VN1179_data_out(5);
    CN335_sign_in(20) <= VN1179_sign_out(5);
    CN335_data_in(21) <= VN1258_data_out(5);
    CN335_sign_in(21) <= VN1258_sign_out(5);
    CN335_data_in(22) <= VN1276_data_out(5);
    CN335_sign_in(22) <= VN1276_sign_out(5);
    CN335_data_in(23) <= VN1285_data_out(5);
    CN335_sign_in(23) <= VN1285_sign_out(5);
    CN335_data_in(24) <= VN1382_data_out(5);
    CN335_sign_in(24) <= VN1382_sign_out(5);
    CN335_data_in(25) <= VN1441_data_out(5);
    CN335_sign_in(25) <= VN1441_sign_out(5);
    CN335_data_in(26) <= VN1541_data_out(5);
    CN335_sign_in(26) <= VN1541_sign_out(5);
    CN335_data_in(27) <= VN1578_data_out(5);
    CN335_sign_in(27) <= VN1578_sign_out(5);
    CN335_data_in(28) <= VN1682_data_out(5);
    CN335_sign_in(28) <= VN1682_sign_out(5);
    CN335_data_in(29) <= VN1845_data_out(5);
    CN335_sign_in(29) <= VN1845_sign_out(5);
    CN335_data_in(30) <= VN1872_data_out(5);
    CN335_sign_in(30) <= VN1872_sign_out(5);
    CN335_data_in(31) <= VN1898_data_out(5);
    CN335_sign_in(31) <= VN1898_sign_out(5);
    CN336_data_in(0) <= VN38_data_out(5);
    CN336_sign_in(0) <= VN38_sign_out(5);
    CN336_data_in(1) <= VN104_data_out(5);
    CN336_sign_in(1) <= VN104_sign_out(5);
    CN336_data_in(2) <= VN121_data_out(5);
    CN336_sign_in(2) <= VN121_sign_out(5);
    CN336_data_in(3) <= VN267_data_out(5);
    CN336_sign_in(3) <= VN267_sign_out(5);
    CN336_data_in(4) <= VN332_data_out(5);
    CN336_sign_in(4) <= VN332_sign_out(5);
    CN336_data_in(5) <= VN344_data_out(5);
    CN336_sign_in(5) <= VN344_sign_out(5);
    CN336_data_in(6) <= VN405_data_out(5);
    CN336_sign_in(6) <= VN405_sign_out(5);
    CN336_data_in(7) <= VN477_data_out(5);
    CN336_sign_in(7) <= VN477_sign_out(5);
    CN336_data_in(8) <= VN506_data_out(5);
    CN336_sign_in(8) <= VN506_sign_out(5);
    CN336_data_in(9) <= VN585_data_out(5);
    CN336_sign_in(9) <= VN585_sign_out(5);
    CN336_data_in(10) <= VN695_data_out(5);
    CN336_sign_in(10) <= VN695_sign_out(5);
    CN336_data_in(11) <= VN757_data_out(5);
    CN336_sign_in(11) <= VN757_sign_out(5);
    CN336_data_in(12) <= VN806_data_out(5);
    CN336_sign_in(12) <= VN806_sign_out(5);
    CN336_data_in(13) <= VN831_data_out(5);
    CN336_sign_in(13) <= VN831_sign_out(5);
    CN336_data_in(14) <= VN909_data_out(5);
    CN336_sign_in(14) <= VN909_sign_out(5);
    CN336_data_in(15) <= VN993_data_out(5);
    CN336_sign_in(15) <= VN993_sign_out(5);
    CN336_data_in(16) <= VN1037_data_out(5);
    CN336_sign_in(16) <= VN1037_sign_out(5);
    CN336_data_in(17) <= VN1082_data_out(5);
    CN336_sign_in(17) <= VN1082_sign_out(5);
    CN336_data_in(18) <= VN1139_data_out(5);
    CN336_sign_in(18) <= VN1139_sign_out(5);
    CN336_data_in(19) <= VN1185_data_out(5);
    CN336_sign_in(19) <= VN1185_sign_out(5);
    CN336_data_in(20) <= VN1329_data_out(5);
    CN336_sign_in(20) <= VN1329_sign_out(5);
    CN336_data_in(21) <= VN1362_data_out(5);
    CN336_sign_in(21) <= VN1362_sign_out(5);
    CN336_data_in(22) <= VN1471_data_out(5);
    CN336_sign_in(22) <= VN1471_sign_out(5);
    CN336_data_in(23) <= VN1543_data_out(5);
    CN336_sign_in(23) <= VN1543_sign_out(5);
    CN336_data_in(24) <= VN1605_data_out(5);
    CN336_sign_in(24) <= VN1605_sign_out(5);
    CN336_data_in(25) <= VN1651_data_out(5);
    CN336_sign_in(25) <= VN1651_sign_out(5);
    CN336_data_in(26) <= VN1692_data_out(5);
    CN336_sign_in(26) <= VN1692_sign_out(5);
    CN336_data_in(27) <= VN1740_data_out(5);
    CN336_sign_in(27) <= VN1740_sign_out(5);
    CN336_data_in(28) <= VN1850_data_out(5);
    CN336_sign_in(28) <= VN1850_sign_out(5);
    CN336_data_in(29) <= VN1935_data_out(5);
    CN336_sign_in(29) <= VN1935_sign_out(5);
    CN336_data_in(30) <= VN1951_data_out(5);
    CN336_sign_in(30) <= VN1951_sign_out(5);
    CN336_data_in(31) <= VN1970_data_out(5);
    CN336_sign_in(31) <= VN1970_sign_out(5);
    CN337_data_in(0) <= VN37_data_out(5);
    CN337_sign_in(0) <= VN37_sign_out(5);
    CN337_data_in(1) <= VN93_data_out(5);
    CN337_sign_in(1) <= VN93_sign_out(5);
    CN337_data_in(2) <= VN115_data_out(5);
    CN337_sign_in(2) <= VN115_sign_out(5);
    CN337_data_in(3) <= VN183_data_out(5);
    CN337_sign_in(3) <= VN183_sign_out(5);
    CN337_data_in(4) <= VN253_data_out(5);
    CN337_sign_in(4) <= VN253_sign_out(5);
    CN337_data_in(5) <= VN290_data_out(5);
    CN337_sign_in(5) <= VN290_sign_out(5);
    CN337_data_in(6) <= VN379_data_out(5);
    CN337_sign_in(6) <= VN379_sign_out(5);
    CN337_data_in(7) <= VN419_data_out(5);
    CN337_sign_in(7) <= VN419_sign_out(5);
    CN337_data_in(8) <= VN475_data_out(5);
    CN337_sign_in(8) <= VN475_sign_out(5);
    CN337_data_in(9) <= VN519_data_out(5);
    CN337_sign_in(9) <= VN519_sign_out(5);
    CN337_data_in(10) <= VN564_data_out(5);
    CN337_sign_in(10) <= VN564_sign_out(5);
    CN337_data_in(11) <= VN714_data_out(5);
    CN337_sign_in(11) <= VN714_sign_out(5);
    CN337_data_in(12) <= VN728_data_out(5);
    CN337_sign_in(12) <= VN728_sign_out(5);
    CN337_data_in(13) <= VN794_data_out(5);
    CN337_sign_in(13) <= VN794_sign_out(5);
    CN337_data_in(14) <= VN862_data_out(5);
    CN337_sign_in(14) <= VN862_sign_out(5);
    CN337_data_in(15) <= VN904_data_out(5);
    CN337_sign_in(15) <= VN904_sign_out(5);
    CN337_data_in(16) <= VN983_data_out(5);
    CN337_sign_in(16) <= VN983_sign_out(5);
    CN337_data_in(17) <= VN1051_data_out(5);
    CN337_sign_in(17) <= VN1051_sign_out(5);
    CN337_data_in(18) <= VN1085_data_out(5);
    CN337_sign_in(18) <= VN1085_sign_out(5);
    CN337_data_in(19) <= VN1126_data_out(5);
    CN337_sign_in(19) <= VN1126_sign_out(5);
    CN337_data_in(20) <= VN1259_data_out(5);
    CN337_sign_in(20) <= VN1259_sign_out(5);
    CN337_data_in(21) <= VN1345_data_out(5);
    CN337_sign_in(21) <= VN1345_sign_out(5);
    CN337_data_in(22) <= VN1405_data_out(5);
    CN337_sign_in(22) <= VN1405_sign_out(5);
    CN337_data_in(23) <= VN1432_data_out(5);
    CN337_sign_in(23) <= VN1432_sign_out(5);
    CN337_data_in(24) <= VN1454_data_out(5);
    CN337_sign_in(24) <= VN1454_sign_out(5);
    CN337_data_in(25) <= VN1590_data_out(5);
    CN337_sign_in(25) <= VN1590_sign_out(5);
    CN337_data_in(26) <= VN1620_data_out(5);
    CN337_sign_in(26) <= VN1620_sign_out(5);
    CN337_data_in(27) <= VN1656_data_out(5);
    CN337_sign_in(27) <= VN1656_sign_out(5);
    CN337_data_in(28) <= VN1705_data_out(5);
    CN337_sign_in(28) <= VN1705_sign_out(5);
    CN337_data_in(29) <= VN1927_data_out(5);
    CN337_sign_in(29) <= VN1927_sign_out(5);
    CN337_data_in(30) <= VN1947_data_out(5);
    CN337_sign_in(30) <= VN1947_sign_out(5);
    CN337_data_in(31) <= VN1958_data_out(5);
    CN337_sign_in(31) <= VN1958_sign_out(5);
    CN338_data_in(0) <= VN36_data_out(5);
    CN338_sign_in(0) <= VN36_sign_out(5);
    CN338_data_in(1) <= VN80_data_out(5);
    CN338_sign_in(1) <= VN80_sign_out(5);
    CN338_data_in(2) <= VN155_data_out(5);
    CN338_sign_in(2) <= VN155_sign_out(5);
    CN338_data_in(3) <= VN190_data_out(5);
    CN338_sign_in(3) <= VN190_sign_out(5);
    CN338_data_in(4) <= VN370_data_out(5);
    CN338_sign_in(4) <= VN370_sign_out(5);
    CN338_data_in(5) <= VN492_data_out(5);
    CN338_sign_in(5) <= VN492_sign_out(5);
    CN338_data_in(6) <= VN540_data_out(5);
    CN338_sign_in(6) <= VN540_sign_out(5);
    CN338_data_in(7) <= VN587_data_out(5);
    CN338_sign_in(7) <= VN587_sign_out(5);
    CN338_data_in(8) <= VN658_data_out(5);
    CN338_sign_in(8) <= VN658_sign_out(5);
    CN338_data_in(9) <= VN669_data_out(5);
    CN338_sign_in(9) <= VN669_sign_out(5);
    CN338_data_in(10) <= VN825_data_out(5);
    CN338_sign_in(10) <= VN825_sign_out(5);
    CN338_data_in(11) <= VN859_data_out(5);
    CN338_sign_in(11) <= VN859_sign_out(5);
    CN338_data_in(12) <= VN962_data_out(5);
    CN338_sign_in(12) <= VN962_sign_out(5);
    CN338_data_in(13) <= VN1006_data_out(5);
    CN338_sign_in(13) <= VN1006_sign_out(5);
    CN338_data_in(14) <= VN1072_data_out(5);
    CN338_sign_in(14) <= VN1072_sign_out(5);
    CN338_data_in(15) <= VN1142_data_out(5);
    CN338_sign_in(15) <= VN1142_sign_out(5);
    CN338_data_in(16) <= VN1197_data_out(5);
    CN338_sign_in(16) <= VN1197_sign_out(5);
    CN338_data_in(17) <= VN1249_data_out(5);
    CN338_sign_in(17) <= VN1249_sign_out(5);
    CN338_data_in(18) <= VN1434_data_out(5);
    CN338_sign_in(18) <= VN1434_sign_out(5);
    CN338_data_in(19) <= VN1452_data_out(5);
    CN338_sign_in(19) <= VN1452_sign_out(5);
    CN338_data_in(20) <= VN1549_data_out(5);
    CN338_sign_in(20) <= VN1549_sign_out(5);
    CN338_data_in(21) <= VN1613_data_out(5);
    CN338_sign_in(21) <= VN1613_sign_out(5);
    CN338_data_in(22) <= VN1677_data_out(5);
    CN338_sign_in(22) <= VN1677_sign_out(5);
    CN338_data_in(23) <= VN1717_data_out(5);
    CN338_sign_in(23) <= VN1717_sign_out(5);
    CN338_data_in(24) <= VN1732_data_out(5);
    CN338_sign_in(24) <= VN1732_sign_out(5);
    CN338_data_in(25) <= VN1770_data_out(5);
    CN338_sign_in(25) <= VN1770_sign_out(5);
    CN338_data_in(26) <= VN1797_data_out(5);
    CN338_sign_in(26) <= VN1797_sign_out(5);
    CN338_data_in(27) <= VN1819_data_out(5);
    CN338_sign_in(27) <= VN1819_sign_out(5);
    CN338_data_in(28) <= VN1822_data_out(5);
    CN338_sign_in(28) <= VN1822_sign_out(5);
    CN338_data_in(29) <= VN1870_data_out(5);
    CN338_sign_in(29) <= VN1870_sign_out(5);
    CN338_data_in(30) <= VN1933_data_out(5);
    CN338_sign_in(30) <= VN1933_sign_out(5);
    CN338_data_in(31) <= VN1941_data_out(5);
    CN338_sign_in(31) <= VN1941_sign_out(5);
    CN339_data_in(0) <= VN35_data_out(5);
    CN339_sign_in(0) <= VN35_sign_out(5);
    CN339_data_in(1) <= VN96_data_out(5);
    CN339_sign_in(1) <= VN96_sign_out(5);
    CN339_data_in(2) <= VN163_data_out(5);
    CN339_sign_in(2) <= VN163_sign_out(5);
    CN339_data_in(3) <= VN216_data_out(5);
    CN339_sign_in(3) <= VN216_sign_out(5);
    CN339_data_in(4) <= VN247_data_out(5);
    CN339_sign_in(4) <= VN247_sign_out(5);
    CN339_data_in(5) <= VN322_data_out(5);
    CN339_sign_in(5) <= VN322_sign_out(5);
    CN339_data_in(6) <= VN389_data_out(5);
    CN339_sign_in(6) <= VN389_sign_out(5);
    CN339_data_in(7) <= VN426_data_out(5);
    CN339_sign_in(7) <= VN426_sign_out(5);
    CN339_data_in(8) <= VN459_data_out(5);
    CN339_sign_in(8) <= VN459_sign_out(5);
    CN339_data_in(9) <= VN550_data_out(5);
    CN339_sign_in(9) <= VN550_sign_out(5);
    CN339_data_in(10) <= VN600_data_out(5);
    CN339_sign_in(10) <= VN600_sign_out(5);
    CN339_data_in(11) <= VN660_data_out(5);
    CN339_sign_in(11) <= VN660_sign_out(5);
    CN339_data_in(12) <= VN718_data_out(5);
    CN339_sign_in(12) <= VN718_sign_out(5);
    CN339_data_in(13) <= VN738_data_out(5);
    CN339_sign_in(13) <= VN738_sign_out(5);
    CN339_data_in(14) <= VN791_data_out(5);
    CN339_sign_in(14) <= VN791_sign_out(5);
    CN339_data_in(15) <= VN873_data_out(5);
    CN339_sign_in(15) <= VN873_sign_out(5);
    CN339_data_in(16) <= VN898_data_out(5);
    CN339_sign_in(16) <= VN898_sign_out(5);
    CN339_data_in(17) <= VN1002_data_out(5);
    CN339_sign_in(17) <= VN1002_sign_out(5);
    CN339_data_in(18) <= VN1032_data_out(5);
    CN339_sign_in(18) <= VN1032_sign_out(5);
    CN339_data_in(19) <= VN1100_data_out(5);
    CN339_sign_in(19) <= VN1100_sign_out(5);
    CN339_data_in(20) <= VN1163_data_out(5);
    CN339_sign_in(20) <= VN1163_sign_out(5);
    CN339_data_in(21) <= VN1203_data_out(5);
    CN339_sign_in(21) <= VN1203_sign_out(5);
    CN339_data_in(22) <= VN1274_data_out(5);
    CN339_sign_in(22) <= VN1274_sign_out(5);
    CN339_data_in(23) <= VN1281_data_out(5);
    CN339_sign_in(23) <= VN1281_sign_out(5);
    CN339_data_in(24) <= VN1299_data_out(5);
    CN339_sign_in(24) <= VN1299_sign_out(5);
    CN339_data_in(25) <= VN1368_data_out(5);
    CN339_sign_in(25) <= VN1368_sign_out(5);
    CN339_data_in(26) <= VN1397_data_out(5);
    CN339_sign_in(26) <= VN1397_sign_out(5);
    CN339_data_in(27) <= VN1563_data_out(5);
    CN339_sign_in(27) <= VN1563_sign_out(5);
    CN339_data_in(28) <= VN1580_data_out(5);
    CN339_sign_in(28) <= VN1580_sign_out(5);
    CN339_data_in(29) <= VN1640_data_out(5);
    CN339_sign_in(29) <= VN1640_sign_out(5);
    CN339_data_in(30) <= VN1649_data_out(5);
    CN339_sign_in(30) <= VN1649_sign_out(5);
    CN339_data_in(31) <= VN1804_data_out(5);
    CN339_sign_in(31) <= VN1804_sign_out(5);
    CN340_data_in(0) <= VN34_data_out(5);
    CN340_sign_in(0) <= VN34_sign_out(5);
    CN340_data_in(1) <= VN58_data_out(5);
    CN340_sign_in(1) <= VN58_sign_out(5);
    CN340_data_in(2) <= VN127_data_out(5);
    CN340_sign_in(2) <= VN127_sign_out(5);
    CN340_data_in(3) <= VN178_data_out(5);
    CN340_sign_in(3) <= VN178_sign_out(5);
    CN340_data_in(4) <= VN245_data_out(5);
    CN340_sign_in(4) <= VN245_sign_out(5);
    CN340_data_in(5) <= VN334_data_out(5);
    CN340_sign_in(5) <= VN334_sign_out(5);
    CN340_data_in(6) <= VN393_data_out(5);
    CN340_sign_in(6) <= VN393_sign_out(5);
    CN340_data_in(7) <= VN460_data_out(5);
    CN340_sign_in(7) <= VN460_sign_out(5);
    CN340_data_in(8) <= VN545_data_out(5);
    CN340_sign_in(8) <= VN545_sign_out(5);
    CN340_data_in(9) <= VN596_data_out(5);
    CN340_sign_in(9) <= VN596_sign_out(5);
    CN340_data_in(10) <= VN629_data_out(5);
    CN340_sign_in(10) <= VN629_sign_out(5);
    CN340_data_in(11) <= VN670_data_out(5);
    CN340_sign_in(11) <= VN670_sign_out(5);
    CN340_data_in(12) <= VN730_data_out(5);
    CN340_sign_in(12) <= VN730_sign_out(5);
    CN340_data_in(13) <= VN816_data_out(5);
    CN340_sign_in(13) <= VN816_sign_out(5);
    CN340_data_in(14) <= VN922_data_out(5);
    CN340_sign_in(14) <= VN922_sign_out(5);
    CN340_data_in(15) <= VN957_data_out(5);
    CN340_sign_in(15) <= VN957_sign_out(5);
    CN340_data_in(16) <= VN1021_data_out(5);
    CN340_sign_in(16) <= VN1021_sign_out(5);
    CN340_data_in(17) <= VN1112_data_out(5);
    CN340_sign_in(17) <= VN1112_sign_out(5);
    CN340_data_in(18) <= VN1188_data_out(5);
    CN340_sign_in(18) <= VN1188_sign_out(5);
    CN340_data_in(19) <= VN1339_data_out(5);
    CN340_sign_in(19) <= VN1339_sign_out(5);
    CN340_data_in(20) <= VN1406_data_out(5);
    CN340_sign_in(20) <= VN1406_sign_out(5);
    CN340_data_in(21) <= VN1489_data_out(5);
    CN340_sign_in(21) <= VN1489_sign_out(5);
    CN340_data_in(22) <= VN1524_data_out(5);
    CN340_sign_in(22) <= VN1524_sign_out(5);
    CN340_data_in(23) <= VN1606_data_out(5);
    CN340_sign_in(23) <= VN1606_sign_out(5);
    CN340_data_in(24) <= VN1693_data_out(5);
    CN340_sign_in(24) <= VN1693_sign_out(5);
    CN340_data_in(25) <= VN1765_data_out(5);
    CN340_sign_in(25) <= VN1765_sign_out(5);
    CN340_data_in(26) <= VN1788_data_out(5);
    CN340_sign_in(26) <= VN1788_sign_out(5);
    CN340_data_in(27) <= VN1828_data_out(5);
    CN340_sign_in(27) <= VN1828_sign_out(5);
    CN340_data_in(28) <= VN1887_data_out(5);
    CN340_sign_in(28) <= VN1887_sign_out(5);
    CN340_data_in(29) <= VN1974_data_out(5);
    CN340_sign_in(29) <= VN1974_sign_out(5);
    CN340_data_in(30) <= VN1978_data_out(5);
    CN340_sign_in(30) <= VN1978_sign_out(5);
    CN340_data_in(31) <= VN1982_data_out(5);
    CN340_sign_in(31) <= VN1982_sign_out(5);
    CN341_data_in(0) <= VN33_data_out(5);
    CN341_sign_in(0) <= VN33_sign_out(5);
    CN341_data_in(1) <= VN68_data_out(5);
    CN341_sign_in(1) <= VN68_sign_out(5);
    CN341_data_in(2) <= VN125_data_out(5);
    CN341_sign_in(2) <= VN125_sign_out(5);
    CN341_data_in(3) <= VN204_data_out(5);
    CN341_sign_in(3) <= VN204_sign_out(5);
    CN341_data_in(4) <= VN258_data_out(5);
    CN341_sign_in(4) <= VN258_sign_out(5);
    CN341_data_in(5) <= VN296_data_out(5);
    CN341_sign_in(5) <= VN296_sign_out(5);
    CN341_data_in(6) <= VN491_data_out(5);
    CN341_sign_in(6) <= VN491_sign_out(5);
    CN341_data_in(7) <= VN551_data_out(5);
    CN341_sign_in(7) <= VN551_sign_out(5);
    CN341_data_in(8) <= VN614_data_out(5);
    CN341_sign_in(8) <= VN614_sign_out(5);
    CN341_data_in(9) <= VN666_data_out(5);
    CN341_sign_in(9) <= VN666_sign_out(5);
    CN341_data_in(10) <= VN842_data_out(5);
    CN341_sign_in(10) <= VN842_sign_out(5);
    CN341_data_in(11) <= VN928_data_out(5);
    CN341_sign_in(11) <= VN928_sign_out(5);
    CN341_data_in(12) <= VN968_data_out(5);
    CN341_sign_in(12) <= VN968_sign_out(5);
    CN341_data_in(13) <= VN1008_data_out(5);
    CN341_sign_in(13) <= VN1008_sign_out(5);
    CN341_data_in(14) <= VN1092_data_out(5);
    CN341_sign_in(14) <= VN1092_sign_out(5);
    CN341_data_in(15) <= VN1165_data_out(5);
    CN341_sign_in(15) <= VN1165_sign_out(5);
    CN341_data_in(16) <= VN1190_data_out(5);
    CN341_sign_in(16) <= VN1190_sign_out(5);
    CN341_data_in(17) <= VN1263_data_out(5);
    CN341_sign_in(17) <= VN1263_sign_out(5);
    CN341_data_in(18) <= VN1313_data_out(5);
    CN341_sign_in(18) <= VN1313_sign_out(5);
    CN341_data_in(19) <= VN1475_data_out(5);
    CN341_sign_in(19) <= VN1475_sign_out(5);
    CN341_data_in(20) <= VN1496_data_out(5);
    CN341_sign_in(20) <= VN1496_sign_out(5);
    CN341_data_in(21) <= VN1542_data_out(5);
    CN341_sign_in(21) <= VN1542_sign_out(5);
    CN341_data_in(22) <= VN1577_data_out(5);
    CN341_sign_in(22) <= VN1577_sign_out(5);
    CN341_data_in(23) <= VN1727_data_out(5);
    CN341_sign_in(23) <= VN1727_sign_out(5);
    CN341_data_in(24) <= VN1767_data_out(5);
    CN341_sign_in(24) <= VN1767_sign_out(5);
    CN341_data_in(25) <= VN1824_data_out(5);
    CN341_sign_in(25) <= VN1824_sign_out(5);
    CN341_data_in(26) <= VN1864_data_out(5);
    CN341_sign_in(26) <= VN1864_sign_out(5);
    CN341_data_in(27) <= VN1879_data_out(5);
    CN341_sign_in(27) <= VN1879_sign_out(5);
    CN341_data_in(28) <= VN1943_data_out(5);
    CN341_sign_in(28) <= VN1943_sign_out(5);
    CN341_data_in(29) <= VN1976_data_out(5);
    CN341_sign_in(29) <= VN1976_sign_out(5);
    CN341_data_in(30) <= VN1977_data_out(5);
    CN341_sign_in(30) <= VN1977_sign_out(5);
    CN341_data_in(31) <= VN1983_data_out(5);
    CN341_sign_in(31) <= VN1983_sign_out(5);
    CN342_data_in(0) <= VN32_data_out(5);
    CN342_sign_in(0) <= VN32_sign_out(5);
    CN342_data_in(1) <= VN63_data_out(5);
    CN342_sign_in(1) <= VN63_sign_out(5);
    CN342_data_in(2) <= VN161_data_out(5);
    CN342_sign_in(2) <= VN161_sign_out(5);
    CN342_data_in(3) <= VN251_data_out(5);
    CN342_sign_in(3) <= VN251_sign_out(5);
    CN342_data_in(4) <= VN294_data_out(5);
    CN342_sign_in(4) <= VN294_sign_out(5);
    CN342_data_in(5) <= VN403_data_out(5);
    CN342_sign_in(5) <= VN403_sign_out(5);
    CN342_data_in(6) <= VN539_data_out(5);
    CN342_sign_in(6) <= VN539_sign_out(5);
    CN342_data_in(7) <= VN581_data_out(5);
    CN342_sign_in(7) <= VN581_sign_out(5);
    CN342_data_in(8) <= VN624_data_out(5);
    CN342_sign_in(8) <= VN624_sign_out(5);
    CN342_data_in(9) <= VN681_data_out(5);
    CN342_sign_in(9) <= VN681_sign_out(5);
    CN342_data_in(10) <= VN735_data_out(5);
    CN342_sign_in(10) <= VN735_sign_out(5);
    CN342_data_in(11) <= VN853_data_out(5);
    CN342_sign_in(11) <= VN853_sign_out(5);
    CN342_data_in(12) <= VN913_data_out(5);
    CN342_sign_in(12) <= VN913_sign_out(5);
    CN342_data_in(13) <= VN997_data_out(5);
    CN342_sign_in(13) <= VN997_sign_out(5);
    CN342_data_in(14) <= VN1024_data_out(5);
    CN342_sign_in(14) <= VN1024_sign_out(5);
    CN342_data_in(15) <= VN1115_data_out(5);
    CN342_sign_in(15) <= VN1115_sign_out(5);
    CN342_data_in(16) <= VN1214_data_out(5);
    CN342_sign_in(16) <= VN1214_sign_out(5);
    CN342_data_in(17) <= VN1265_data_out(5);
    CN342_sign_in(17) <= VN1265_sign_out(5);
    CN342_data_in(18) <= VN1284_data_out(5);
    CN342_sign_in(18) <= VN1284_sign_out(5);
    CN342_data_in(19) <= VN1370_data_out(5);
    CN342_sign_in(19) <= VN1370_sign_out(5);
    CN342_data_in(20) <= VN1455_data_out(5);
    CN342_sign_in(20) <= VN1455_sign_out(5);
    CN342_data_in(21) <= VN1564_data_out(5);
    CN342_sign_in(21) <= VN1564_sign_out(5);
    CN342_data_in(22) <= VN1598_data_out(5);
    CN342_sign_in(22) <= VN1598_sign_out(5);
    CN342_data_in(23) <= VN1647_data_out(5);
    CN342_sign_in(23) <= VN1647_sign_out(5);
    CN342_data_in(24) <= VN1711_data_out(5);
    CN342_sign_in(24) <= VN1711_sign_out(5);
    CN342_data_in(25) <= VN1769_data_out(5);
    CN342_sign_in(25) <= VN1769_sign_out(5);
    CN342_data_in(26) <= VN1773_data_out(5);
    CN342_sign_in(26) <= VN1773_sign_out(5);
    CN342_data_in(27) <= VN1798_data_out(5);
    CN342_sign_in(27) <= VN1798_sign_out(5);
    CN342_data_in(28) <= VN1815_data_out(5);
    CN342_sign_in(28) <= VN1815_sign_out(5);
    CN342_data_in(29) <= VN1840_data_out(5);
    CN342_sign_in(29) <= VN1840_sign_out(5);
    CN342_data_in(30) <= VN1853_data_out(5);
    CN342_sign_in(30) <= VN1853_sign_out(5);
    CN342_data_in(31) <= VN1899_data_out(5);
    CN342_sign_in(31) <= VN1899_sign_out(5);
    CN343_data_in(0) <= VN31_data_out(5);
    CN343_sign_in(0) <= VN31_sign_out(5);
    CN343_data_in(1) <= VN69_data_out(5);
    CN343_sign_in(1) <= VN69_sign_out(5);
    CN343_data_in(2) <= VN140_data_out(5);
    CN343_sign_in(2) <= VN140_sign_out(5);
    CN343_data_in(3) <= VN206_data_out(5);
    CN343_sign_in(3) <= VN206_sign_out(5);
    CN343_data_in(4) <= VN228_data_out(5);
    CN343_sign_in(4) <= VN228_sign_out(5);
    CN343_data_in(5) <= VN327_data_out(5);
    CN343_sign_in(5) <= VN327_sign_out(5);
    CN343_data_in(6) <= VN387_data_out(5);
    CN343_sign_in(6) <= VN387_sign_out(5);
    CN343_data_in(7) <= VN422_data_out(5);
    CN343_sign_in(7) <= VN422_sign_out(5);
    CN343_data_in(8) <= VN501_data_out(5);
    CN343_sign_in(8) <= VN501_sign_out(5);
    CN343_data_in(9) <= VN508_data_out(5);
    CN343_sign_in(9) <= VN508_sign_out(5);
    CN343_data_in(10) <= VN582_data_out(5);
    CN343_sign_in(10) <= VN582_sign_out(5);
    CN343_data_in(11) <= VN688_data_out(5);
    CN343_sign_in(11) <= VN688_sign_out(5);
    CN343_data_in(12) <= VN765_data_out(5);
    CN343_sign_in(12) <= VN765_sign_out(5);
    CN343_data_in(13) <= VN818_data_out(5);
    CN343_sign_in(13) <= VN818_sign_out(5);
    CN343_data_in(14) <= VN846_data_out(5);
    CN343_sign_in(14) <= VN846_sign_out(5);
    CN343_data_in(15) <= VN985_data_out(5);
    CN343_sign_in(15) <= VN985_sign_out(5);
    CN343_data_in(16) <= VN1043_data_out(5);
    CN343_sign_in(16) <= VN1043_sign_out(5);
    CN343_data_in(17) <= VN1101_data_out(5);
    CN343_sign_in(17) <= VN1101_sign_out(5);
    CN343_data_in(18) <= VN1162_data_out(5);
    CN343_sign_in(18) <= VN1162_sign_out(5);
    CN343_data_in(19) <= VN1195_data_out(5);
    CN343_sign_in(19) <= VN1195_sign_out(5);
    CN343_data_in(20) <= VN1235_data_out(5);
    CN343_sign_in(20) <= VN1235_sign_out(5);
    CN343_data_in(21) <= VN1282_data_out(5);
    CN343_sign_in(21) <= VN1282_sign_out(5);
    CN343_data_in(22) <= VN1305_data_out(5);
    CN343_sign_in(22) <= VN1305_sign_out(5);
    CN343_data_in(23) <= VN1433_data_out(5);
    CN343_sign_in(23) <= VN1433_sign_out(5);
    CN343_data_in(24) <= VN1535_data_out(5);
    CN343_sign_in(24) <= VN1535_sign_out(5);
    CN343_data_in(25) <= VN1637_data_out(5);
    CN343_sign_in(25) <= VN1637_sign_out(5);
    CN343_data_in(26) <= VN1678_data_out(5);
    CN343_sign_in(26) <= VN1678_sign_out(5);
    CN343_data_in(27) <= VN1691_data_out(5);
    CN343_sign_in(27) <= VN1691_sign_out(5);
    CN343_data_in(28) <= VN1799_data_out(5);
    CN343_sign_in(28) <= VN1799_sign_out(5);
    CN343_data_in(29) <= VN1825_data_out(5);
    CN343_sign_in(29) <= VN1825_sign_out(5);
    CN343_data_in(30) <= VN1841_data_out(5);
    CN343_sign_in(30) <= VN1841_sign_out(5);
    CN343_data_in(31) <= VN1900_data_out(5);
    CN343_sign_in(31) <= VN1900_sign_out(5);
    CN344_data_in(0) <= VN30_data_out(5);
    CN344_sign_in(0) <= VN30_sign_out(5);
    CN344_data_in(1) <= VN57_data_out(5);
    CN344_sign_in(1) <= VN57_sign_out(5);
    CN344_data_in(2) <= VN143_data_out(5);
    CN344_sign_in(2) <= VN143_sign_out(5);
    CN344_data_in(3) <= VN218_data_out(5);
    CN344_sign_in(3) <= VN218_sign_out(5);
    CN344_data_in(4) <= VN238_data_out(5);
    CN344_sign_in(4) <= VN238_sign_out(5);
    CN344_data_in(5) <= VN307_data_out(5);
    CN344_sign_in(5) <= VN307_sign_out(5);
    CN344_data_in(6) <= VN367_data_out(5);
    CN344_sign_in(6) <= VN367_sign_out(5);
    CN344_data_in(7) <= VN443_data_out(5);
    CN344_sign_in(7) <= VN443_sign_out(5);
    CN344_data_in(8) <= VN449_data_out(5);
    CN344_sign_in(8) <= VN449_sign_out(5);
    CN344_data_in(9) <= VN514_data_out(5);
    CN344_sign_in(9) <= VN514_sign_out(5);
    CN344_data_in(10) <= VN613_data_out(5);
    CN344_sign_in(10) <= VN613_sign_out(5);
    CN344_data_in(11) <= VN659_data_out(5);
    CN344_sign_in(11) <= VN659_sign_out(5);
    CN344_data_in(12) <= VN673_data_out(5);
    CN344_sign_in(12) <= VN673_sign_out(5);
    CN344_data_in(13) <= VN763_data_out(5);
    CN344_sign_in(13) <= VN763_sign_out(5);
    CN344_data_in(14) <= VN805_data_out(5);
    CN344_sign_in(14) <= VN805_sign_out(5);
    CN344_data_in(15) <= VN850_data_out(5);
    CN344_sign_in(15) <= VN850_sign_out(5);
    CN344_data_in(16) <= VN938_data_out(5);
    CN344_sign_in(16) <= VN938_sign_out(5);
    CN344_data_in(17) <= VN971_data_out(5);
    CN344_sign_in(17) <= VN971_sign_out(5);
    CN344_data_in(18) <= VN1053_data_out(5);
    CN344_sign_in(18) <= VN1053_sign_out(5);
    CN344_data_in(19) <= VN1094_data_out(5);
    CN344_sign_in(19) <= VN1094_sign_out(5);
    CN344_data_in(20) <= VN1129_data_out(5);
    CN344_sign_in(20) <= VN1129_sign_out(5);
    CN344_data_in(21) <= VN1207_data_out(5);
    CN344_sign_in(21) <= VN1207_sign_out(5);
    CN344_data_in(22) <= VN1272_data_out(5);
    CN344_sign_in(22) <= VN1272_sign_out(5);
    CN344_data_in(23) <= VN1293_data_out(5);
    CN344_sign_in(23) <= VN1293_sign_out(5);
    CN344_data_in(24) <= VN1351_data_out(5);
    CN344_sign_in(24) <= VN1351_sign_out(5);
    CN344_data_in(25) <= VN1400_data_out(5);
    CN344_sign_in(25) <= VN1400_sign_out(5);
    CN344_data_in(26) <= VN1451_data_out(5);
    CN344_sign_in(26) <= VN1451_sign_out(5);
    CN344_data_in(27) <= VN1459_data_out(5);
    CN344_sign_in(27) <= VN1459_sign_out(5);
    CN344_data_in(28) <= VN1470_data_out(5);
    CN344_sign_in(28) <= VN1470_sign_out(5);
    CN344_data_in(29) <= VN1621_data_out(5);
    CN344_sign_in(29) <= VN1621_sign_out(5);
    CN344_data_in(30) <= VN1675_data_out(5);
    CN344_sign_in(30) <= VN1675_sign_out(5);
    CN344_data_in(31) <= VN1805_data_out(5);
    CN344_sign_in(31) <= VN1805_sign_out(5);
    CN345_data_in(0) <= VN29_data_out(5);
    CN345_sign_in(0) <= VN29_sign_out(5);
    CN345_data_in(1) <= VN83_data_out(5);
    CN345_sign_in(1) <= VN83_sign_out(5);
    CN345_data_in(2) <= VN128_data_out(5);
    CN345_sign_in(2) <= VN128_sign_out(5);
    CN345_data_in(3) <= VN232_data_out(5);
    CN345_sign_in(3) <= VN232_sign_out(5);
    CN345_data_in(4) <= VN309_data_out(5);
    CN345_sign_in(4) <= VN309_sign_out(5);
    CN345_data_in(5) <= VN375_data_out(5);
    CN345_sign_in(5) <= VN375_sign_out(5);
    CN345_data_in(6) <= VN444_data_out(5);
    CN345_sign_in(6) <= VN444_sign_out(5);
    CN345_data_in(7) <= VN505_data_out(5);
    CN345_sign_in(7) <= VN505_sign_out(5);
    CN345_data_in(8) <= VN554_data_out(5);
    CN345_sign_in(8) <= VN554_sign_out(5);
    CN345_data_in(9) <= VN605_data_out(5);
    CN345_sign_in(9) <= VN605_sign_out(5);
    CN345_data_in(10) <= VN674_data_out(5);
    CN345_sign_in(10) <= VN674_sign_out(5);
    CN345_data_in(11) <= VN776_data_out(5);
    CN345_sign_in(11) <= VN776_sign_out(5);
    CN345_data_in(12) <= VN823_data_out(5);
    CN345_sign_in(12) <= VN823_sign_out(5);
    CN345_data_in(13) <= VN839_data_out(5);
    CN345_sign_in(13) <= VN839_sign_out(5);
    CN345_data_in(14) <= VN921_data_out(5);
    CN345_sign_in(14) <= VN921_sign_out(5);
    CN345_data_in(15) <= VN988_data_out(5);
    CN345_sign_in(15) <= VN988_sign_out(5);
    CN345_data_in(16) <= VN1048_data_out(5);
    CN345_sign_in(16) <= VN1048_sign_out(5);
    CN345_data_in(17) <= VN1083_data_out(5);
    CN345_sign_in(17) <= VN1083_sign_out(5);
    CN345_data_in(18) <= VN1135_data_out(5);
    CN345_sign_in(18) <= VN1135_sign_out(5);
    CN345_data_in(19) <= VN1222_data_out(5);
    CN345_sign_in(19) <= VN1222_sign_out(5);
    CN345_data_in(20) <= VN1228_data_out(5);
    CN345_sign_in(20) <= VN1228_sign_out(5);
    CN345_data_in(21) <= VN1315_data_out(5);
    CN345_sign_in(21) <= VN1315_sign_out(5);
    CN345_data_in(22) <= VN1359_data_out(5);
    CN345_sign_in(22) <= VN1359_sign_out(5);
    CN345_data_in(23) <= VN1385_data_out(5);
    CN345_sign_in(23) <= VN1385_sign_out(5);
    CN345_data_in(24) <= VN1423_data_out(5);
    CN345_sign_in(24) <= VN1423_sign_out(5);
    CN345_data_in(25) <= VN1493_data_out(5);
    CN345_sign_in(25) <= VN1493_sign_out(5);
    CN345_data_in(26) <= VN1737_data_out(5);
    CN345_sign_in(26) <= VN1737_sign_out(5);
    CN345_data_in(27) <= VN1835_data_out(5);
    CN345_sign_in(27) <= VN1835_sign_out(5);
    CN345_data_in(28) <= VN1966_data_out(5);
    CN345_sign_in(28) <= VN1966_sign_out(5);
    CN345_data_in(29) <= VN1994_data_out(5);
    CN345_sign_in(29) <= VN1994_sign_out(5);
    CN345_data_in(30) <= VN2004_data_out(5);
    CN345_sign_in(30) <= VN2004_sign_out(5);
    CN345_data_in(31) <= VN2014_data_out(5);
    CN345_sign_in(31) <= VN2014_sign_out(5);
    CN346_data_in(0) <= VN28_data_out(5);
    CN346_sign_in(0) <= VN28_sign_out(5);
    CN346_data_in(1) <= VN89_data_out(5);
    CN346_sign_in(1) <= VN89_sign_out(5);
    CN346_data_in(2) <= VN162_data_out(5);
    CN346_sign_in(2) <= VN162_sign_out(5);
    CN346_data_in(3) <= VN181_data_out(5);
    CN346_sign_in(3) <= VN181_sign_out(5);
    CN346_data_in(4) <= VN235_data_out(5);
    CN346_sign_in(4) <= VN235_sign_out(5);
    CN346_data_in(5) <= VN297_data_out(5);
    CN346_sign_in(5) <= VN297_sign_out(5);
    CN346_data_in(6) <= VN339_data_out(5);
    CN346_sign_in(6) <= VN339_sign_out(5);
    CN346_data_in(7) <= VN421_data_out(5);
    CN346_sign_in(7) <= VN421_sign_out(5);
    CN346_data_in(8) <= VN448_data_out(5);
    CN346_sign_in(8) <= VN448_sign_out(5);
    CN346_data_in(9) <= VN556_data_out(5);
    CN346_sign_in(9) <= VN556_sign_out(5);
    CN346_data_in(10) <= VN568_data_out(5);
    CN346_sign_in(10) <= VN568_sign_out(5);
    CN346_data_in(11) <= VN647_data_out(5);
    CN346_sign_in(11) <= VN647_sign_out(5);
    CN346_data_in(12) <= VN699_data_out(5);
    CN346_sign_in(12) <= VN699_sign_out(5);
    CN346_data_in(13) <= VN770_data_out(5);
    CN346_sign_in(13) <= VN770_sign_out(5);
    CN346_data_in(14) <= VN798_data_out(5);
    CN346_sign_in(14) <= VN798_sign_out(5);
    CN346_data_in(15) <= VN874_data_out(5);
    CN346_sign_in(15) <= VN874_sign_out(5);
    CN346_data_in(16) <= VN949_data_out(5);
    CN346_sign_in(16) <= VN949_sign_out(5);
    CN346_data_in(17) <= VN1054_data_out(5);
    CN346_sign_in(17) <= VN1054_sign_out(5);
    CN346_data_in(18) <= VN1059_data_out(5);
    CN346_sign_in(18) <= VN1059_sign_out(5);
    CN346_data_in(19) <= VN1098_data_out(5);
    CN346_sign_in(19) <= VN1098_sign_out(5);
    CN346_data_in(20) <= VN1119_data_out(5);
    CN346_sign_in(20) <= VN1119_sign_out(5);
    CN346_data_in(21) <= VN1189_data_out(5);
    CN346_sign_in(21) <= VN1189_sign_out(5);
    CN346_data_in(22) <= VN1236_data_out(5);
    CN346_sign_in(22) <= VN1236_sign_out(5);
    CN346_data_in(23) <= VN1307_data_out(5);
    CN346_sign_in(23) <= VN1307_sign_out(5);
    CN346_data_in(24) <= VN1355_data_out(5);
    CN346_sign_in(24) <= VN1355_sign_out(5);
    CN346_data_in(25) <= VN1457_data_out(5);
    CN346_sign_in(25) <= VN1457_sign_out(5);
    CN346_data_in(26) <= VN1544_data_out(5);
    CN346_sign_in(26) <= VN1544_sign_out(5);
    CN346_data_in(27) <= VN1616_data_out(5);
    CN346_sign_in(27) <= VN1616_sign_out(5);
    CN346_data_in(28) <= VN1665_data_out(5);
    CN346_sign_in(28) <= VN1665_sign_out(5);
    CN346_data_in(29) <= VN1746_data_out(5);
    CN346_sign_in(29) <= VN1746_sign_out(5);
    CN346_data_in(30) <= VN1789_data_out(5);
    CN346_sign_in(30) <= VN1789_sign_out(5);
    CN346_data_in(31) <= VN1874_data_out(5);
    CN346_sign_in(31) <= VN1874_sign_out(5);
    CN347_data_in(0) <= VN27_data_out(5);
    CN347_sign_in(0) <= VN27_sign_out(5);
    CN347_data_in(1) <= VN73_data_out(5);
    CN347_sign_in(1) <= VN73_sign_out(5);
    CN347_data_in(2) <= VN124_data_out(5);
    CN347_sign_in(2) <= VN124_sign_out(5);
    CN347_data_in(3) <= VN199_data_out(5);
    CN347_sign_in(3) <= VN199_sign_out(5);
    CN347_data_in(4) <= VN225_data_out(5);
    CN347_sign_in(4) <= VN225_sign_out(5);
    CN347_data_in(5) <= VN328_data_out(5);
    CN347_sign_in(5) <= VN328_sign_out(5);
    CN347_data_in(6) <= VN337_data_out(5);
    CN347_sign_in(6) <= VN337_sign_out(5);
    CN347_data_in(7) <= VN412_data_out(5);
    CN347_sign_in(7) <= VN412_sign_out(5);
    CN347_data_in(8) <= VN499_data_out(5);
    CN347_sign_in(8) <= VN499_sign_out(5);
    CN347_data_in(9) <= VN523_data_out(5);
    CN347_sign_in(9) <= VN523_sign_out(5);
    CN347_data_in(10) <= VN572_data_out(5);
    CN347_sign_in(10) <= VN572_sign_out(5);
    CN347_data_in(11) <= VN625_data_out(5);
    CN347_sign_in(11) <= VN625_sign_out(5);
    CN347_data_in(12) <= VN680_data_out(5);
    CN347_sign_in(12) <= VN680_sign_out(5);
    CN347_data_in(13) <= VN745_data_out(5);
    CN347_sign_in(13) <= VN745_sign_out(5);
    CN347_data_in(14) <= VN796_data_out(5);
    CN347_sign_in(14) <= VN796_sign_out(5);
    CN347_data_in(15) <= VN858_data_out(5);
    CN347_sign_in(15) <= VN858_sign_out(5);
    CN347_data_in(16) <= VN939_data_out(5);
    CN347_sign_in(16) <= VN939_sign_out(5);
    CN347_data_in(17) <= VN959_data_out(5);
    CN347_sign_in(17) <= VN959_sign_out(5);
    CN347_data_in(18) <= VN1042_data_out(5);
    CN347_sign_in(18) <= VN1042_sign_out(5);
    CN347_data_in(19) <= VN1077_data_out(5);
    CN347_sign_in(19) <= VN1077_sign_out(5);
    CN347_data_in(20) <= VN1121_data_out(5);
    CN347_sign_in(20) <= VN1121_sign_out(5);
    CN347_data_in(21) <= VN1202_data_out(5);
    CN347_sign_in(21) <= VN1202_sign_out(5);
    CN347_data_in(22) <= VN1264_data_out(5);
    CN347_sign_in(22) <= VN1264_sign_out(5);
    CN347_data_in(23) <= VN1297_data_out(5);
    CN347_sign_in(23) <= VN1297_sign_out(5);
    CN347_data_in(24) <= VN1330_data_out(5);
    CN347_sign_in(24) <= VN1330_sign_out(5);
    CN347_data_in(25) <= VN1360_data_out(5);
    CN347_sign_in(25) <= VN1360_sign_out(5);
    CN347_data_in(26) <= VN1387_data_out(5);
    CN347_sign_in(26) <= VN1387_sign_out(5);
    CN347_data_in(27) <= VN1540_data_out(5);
    CN347_sign_in(27) <= VN1540_sign_out(5);
    CN347_data_in(28) <= VN1604_data_out(5);
    CN347_sign_in(28) <= VN1604_sign_out(5);
    CN347_data_in(29) <= VN1666_data_out(5);
    CN347_sign_in(29) <= VN1666_sign_out(5);
    CN347_data_in(30) <= VN1710_data_out(5);
    CN347_sign_in(30) <= VN1710_sign_out(5);
    CN347_data_in(31) <= VN1806_data_out(5);
    CN347_sign_in(31) <= VN1806_sign_out(5);
    CN348_data_in(0) <= VN26_data_out(5);
    CN348_sign_in(0) <= VN26_sign_out(5);
    CN348_data_in(1) <= VN75_data_out(5);
    CN348_sign_in(1) <= VN75_sign_out(5);
    CN348_data_in(2) <= VN152_data_out(5);
    CN348_sign_in(2) <= VN152_sign_out(5);
    CN348_data_in(3) <= VN200_data_out(5);
    CN348_sign_in(3) <= VN200_sign_out(5);
    CN348_data_in(4) <= VN259_data_out(5);
    CN348_sign_in(4) <= VN259_sign_out(5);
    CN348_data_in(5) <= VN293_data_out(5);
    CN348_sign_in(5) <= VN293_sign_out(5);
    CN348_data_in(6) <= VN373_data_out(5);
    CN348_sign_in(6) <= VN373_sign_out(5);
    CN348_data_in(7) <= VN430_data_out(5);
    CN348_sign_in(7) <= VN430_sign_out(5);
    CN348_data_in(8) <= VN481_data_out(5);
    CN348_sign_in(8) <= VN481_sign_out(5);
    CN348_data_in(9) <= VN507_data_out(5);
    CN348_sign_in(9) <= VN507_sign_out(5);
    CN348_data_in(10) <= VN616_data_out(5);
    CN348_sign_in(10) <= VN616_sign_out(5);
    CN348_data_in(11) <= VN649_data_out(5);
    CN348_sign_in(11) <= VN649_sign_out(5);
    CN348_data_in(12) <= VN691_data_out(5);
    CN348_sign_in(12) <= VN691_sign_out(5);
    CN348_data_in(13) <= VN755_data_out(5);
    CN348_sign_in(13) <= VN755_sign_out(5);
    CN348_data_in(14) <= VN809_data_out(5);
    CN348_sign_in(14) <= VN809_sign_out(5);
    CN348_data_in(15) <= VN869_data_out(5);
    CN348_sign_in(15) <= VN869_sign_out(5);
    CN348_data_in(16) <= VN914_data_out(5);
    CN348_sign_in(16) <= VN914_sign_out(5);
    CN348_data_in(17) <= VN954_data_out(5);
    CN348_sign_in(17) <= VN954_sign_out(5);
    CN348_data_in(18) <= VN1011_data_out(5);
    CN348_sign_in(18) <= VN1011_sign_out(5);
    CN348_data_in(19) <= VN1074_data_out(5);
    CN348_sign_in(19) <= VN1074_sign_out(5);
    CN348_data_in(20) <= VN1146_data_out(5);
    CN348_sign_in(20) <= VN1146_sign_out(5);
    CN348_data_in(21) <= VN1176_data_out(5);
    CN348_sign_in(21) <= VN1176_sign_out(5);
    CN348_data_in(22) <= VN1224_data_out(5);
    CN348_sign_in(22) <= VN1224_sign_out(5);
    CN348_data_in(23) <= VN1312_data_out(5);
    CN348_sign_in(23) <= VN1312_sign_out(5);
    CN348_data_in(24) <= VN1350_data_out(5);
    CN348_sign_in(24) <= VN1350_sign_out(5);
    CN348_data_in(25) <= VN1490_data_out(5);
    CN348_sign_in(25) <= VN1490_sign_out(5);
    CN348_data_in(26) <= VN1523_data_out(5);
    CN348_sign_in(26) <= VN1523_sign_out(5);
    CN348_data_in(27) <= VN1584_data_out(5);
    CN348_sign_in(27) <= VN1584_sign_out(5);
    CN348_data_in(28) <= VN1696_data_out(5);
    CN348_sign_in(28) <= VN1696_sign_out(5);
    CN348_data_in(29) <= VN1752_data_out(5);
    CN348_sign_in(29) <= VN1752_sign_out(5);
    CN348_data_in(30) <= VN1908_data_out(5);
    CN348_sign_in(30) <= VN1908_sign_out(5);
    CN348_data_in(31) <= VN1918_data_out(5);
    CN348_sign_in(31) <= VN1918_sign_out(5);
    CN349_data_in(0) <= VN25_data_out(5);
    CN349_sign_in(0) <= VN25_sign_out(5);
    CN349_data_in(1) <= VN99_data_out(5);
    CN349_sign_in(1) <= VN99_sign_out(5);
    CN349_data_in(2) <= VN180_data_out(5);
    CN349_sign_in(2) <= VN180_sign_out(5);
    CN349_data_in(3) <= VN244_data_out(5);
    CN349_sign_in(3) <= VN244_sign_out(5);
    CN349_data_in(4) <= VN319_data_out(5);
    CN349_sign_in(4) <= VN319_sign_out(5);
    CN349_data_in(5) <= VN352_data_out(5);
    CN349_sign_in(5) <= VN352_sign_out(5);
    CN349_data_in(6) <= VN435_data_out(5);
    CN349_sign_in(6) <= VN435_sign_out(5);
    CN349_data_in(7) <= VN487_data_out(5);
    CN349_sign_in(7) <= VN487_sign_out(5);
    CN349_data_in(8) <= VN571_data_out(5);
    CN349_sign_in(8) <= VN571_sign_out(5);
    CN349_data_in(9) <= VN661_data_out(5);
    CN349_sign_in(9) <= VN661_sign_out(5);
    CN349_data_in(10) <= VN700_data_out(5);
    CN349_sign_in(10) <= VN700_sign_out(5);
    CN349_data_in(11) <= VN802_data_out(5);
    CN349_sign_in(11) <= VN802_sign_out(5);
    CN349_data_in(12) <= VN880_data_out(5);
    CN349_sign_in(12) <= VN880_sign_out(5);
    CN349_data_in(13) <= VN927_data_out(5);
    CN349_sign_in(13) <= VN927_sign_out(5);
    CN349_data_in(14) <= VN960_data_out(5);
    CN349_sign_in(14) <= VN960_sign_out(5);
    CN349_data_in(15) <= VN1017_data_out(5);
    CN349_sign_in(15) <= VN1017_sign_out(5);
    CN349_data_in(16) <= VN1113_data_out(5);
    CN349_sign_in(16) <= VN1113_sign_out(5);
    CN349_data_in(17) <= VN1127_data_out(5);
    CN349_sign_in(17) <= VN1127_sign_out(5);
    CN349_data_in(18) <= VN1210_data_out(5);
    CN349_sign_in(18) <= VN1210_sign_out(5);
    CN349_data_in(19) <= VN1251_data_out(5);
    CN349_sign_in(19) <= VN1251_sign_out(5);
    CN349_data_in(20) <= VN1290_data_out(5);
    CN349_sign_in(20) <= VN1290_sign_out(5);
    CN349_data_in(21) <= VN1373_data_out(5);
    CN349_sign_in(21) <= VN1373_sign_out(5);
    CN349_data_in(22) <= VN1417_data_out(5);
    CN349_sign_in(22) <= VN1417_sign_out(5);
    CN349_data_in(23) <= VN1431_data_out(5);
    CN349_sign_in(23) <= VN1431_sign_out(5);
    CN349_data_in(24) <= VN1582_data_out(5);
    CN349_sign_in(24) <= VN1582_sign_out(5);
    CN349_data_in(25) <= VN1639_data_out(5);
    CN349_sign_in(25) <= VN1639_sign_out(5);
    CN349_data_in(26) <= VN1683_data_out(5);
    CN349_sign_in(26) <= VN1683_sign_out(5);
    CN349_data_in(27) <= VN1728_data_out(5);
    CN349_sign_in(27) <= VN1728_sign_out(5);
    CN349_data_in(28) <= VN1818_data_out(5);
    CN349_sign_in(28) <= VN1818_sign_out(5);
    CN349_data_in(29) <= VN1842_data_out(5);
    CN349_sign_in(29) <= VN1842_sign_out(5);
    CN349_data_in(30) <= VN1863_data_out(5);
    CN349_sign_in(30) <= VN1863_sign_out(5);
    CN349_data_in(31) <= VN1901_data_out(5);
    CN349_sign_in(31) <= VN1901_sign_out(5);
    CN350_data_in(0) <= VN24_data_out(5);
    CN350_sign_in(0) <= VN24_sign_out(5);
    CN350_data_in(1) <= VN81_data_out(5);
    CN350_sign_in(1) <= VN81_sign_out(5);
    CN350_data_in(2) <= VN164_data_out(5);
    CN350_sign_in(2) <= VN164_sign_out(5);
    CN350_data_in(3) <= VN171_data_out(5);
    CN350_sign_in(3) <= VN171_sign_out(5);
    CN350_data_in(4) <= VN254_data_out(5);
    CN350_sign_in(4) <= VN254_sign_out(5);
    CN350_data_in(5) <= VN303_data_out(5);
    CN350_sign_in(5) <= VN303_sign_out(5);
    CN350_data_in(6) <= VN447_data_out(5);
    CN350_sign_in(6) <= VN447_sign_out(5);
    CN350_data_in(7) <= VN455_data_out(5);
    CN350_sign_in(7) <= VN455_sign_out(5);
    CN350_data_in(8) <= VN566_data_out(5);
    CN350_sign_in(8) <= VN566_sign_out(5);
    CN350_data_in(9) <= VN657_data_out(5);
    CN350_sign_in(9) <= VN657_sign_out(5);
    CN350_data_in(10) <= VN752_data_out(5);
    CN350_sign_in(10) <= VN752_sign_out(5);
    CN350_data_in(11) <= VN854_data_out(5);
    CN350_sign_in(11) <= VN854_sign_out(5);
    CN350_data_in(12) <= VN900_data_out(5);
    CN350_sign_in(12) <= VN900_sign_out(5);
    CN350_data_in(13) <= VN948_data_out(5);
    CN350_sign_in(13) <= VN948_sign_out(5);
    CN350_data_in(14) <= VN1058_data_out(5);
    CN350_sign_in(14) <= VN1058_sign_out(5);
    CN350_data_in(15) <= VN1080_data_out(5);
    CN350_sign_in(15) <= VN1080_sign_out(5);
    CN350_data_in(16) <= VN1177_data_out(5);
    CN350_sign_in(16) <= VN1177_sign_out(5);
    CN350_data_in(17) <= VN1231_data_out(5);
    CN350_sign_in(17) <= VN1231_sign_out(5);
    CN350_data_in(18) <= VN1280_data_out(5);
    CN350_sign_in(18) <= VN1280_sign_out(5);
    CN350_data_in(19) <= VN1287_data_out(5);
    CN350_sign_in(19) <= VN1287_sign_out(5);
    CN350_data_in(20) <= VN1379_data_out(5);
    CN350_sign_in(20) <= VN1379_sign_out(5);
    CN350_data_in(21) <= VN1418_data_out(5);
    CN350_sign_in(21) <= VN1418_sign_out(5);
    CN350_data_in(22) <= VN1473_data_out(5);
    CN350_sign_in(22) <= VN1473_sign_out(5);
    CN350_data_in(23) <= VN1592_data_out(5);
    CN350_sign_in(23) <= VN1592_sign_out(5);
    CN350_data_in(24) <= VN1655_data_out(5);
    CN350_sign_in(24) <= VN1655_sign_out(5);
    CN350_data_in(25) <= VN1700_data_out(5);
    CN350_sign_in(25) <= VN1700_sign_out(5);
    CN350_data_in(26) <= VN1839_data_out(5);
    CN350_sign_in(26) <= VN1839_sign_out(5);
    CN350_data_in(27) <= VN1942_data_out(5);
    CN350_sign_in(27) <= VN1942_sign_out(5);
    CN350_data_in(28) <= VN1964_data_out(5);
    CN350_sign_in(28) <= VN1964_sign_out(5);
    CN350_data_in(29) <= VN1987_data_out(5);
    CN350_sign_in(29) <= VN1987_sign_out(5);
    CN350_data_in(30) <= VN2043_data_out(5);
    CN350_sign_in(30) <= VN2043_sign_out(5);
    CN350_data_in(31) <= VN2047_data_out(5);
    CN350_sign_in(31) <= VN2047_sign_out(5);
    CN351_data_in(0) <= VN23_data_out(5);
    CN351_sign_in(0) <= VN23_sign_out(5);
    CN351_data_in(1) <= VN154_data_out(5);
    CN351_sign_in(1) <= VN154_sign_out(5);
    CN351_data_in(2) <= VN188_data_out(5);
    CN351_sign_in(2) <= VN188_sign_out(5);
    CN351_data_in(3) <= VN266_data_out(5);
    CN351_sign_in(3) <= VN266_sign_out(5);
    CN351_data_in(4) <= VN329_data_out(5);
    CN351_sign_in(4) <= VN329_sign_out(5);
    CN351_data_in(5) <= VN340_data_out(5);
    CN351_sign_in(5) <= VN340_sign_out(5);
    CN351_data_in(6) <= VN434_data_out(5);
    CN351_sign_in(6) <= VN434_sign_out(5);
    CN351_data_in(7) <= VN453_data_out(5);
    CN351_sign_in(7) <= VN453_sign_out(5);
    CN351_data_in(8) <= VN555_data_out(5);
    CN351_sign_in(8) <= VN555_sign_out(5);
    CN351_data_in(9) <= VN622_data_out(5);
    CN351_sign_in(9) <= VN622_sign_out(5);
    CN351_data_in(10) <= VN687_data_out(5);
    CN351_sign_in(10) <= VN687_sign_out(5);
    CN351_data_in(11) <= VN743_data_out(5);
    CN351_sign_in(11) <= VN743_sign_out(5);
    CN351_data_in(12) <= VN789_data_out(5);
    CN351_sign_in(12) <= VN789_sign_out(5);
    CN351_data_in(13) <= VN830_data_out(5);
    CN351_sign_in(13) <= VN830_sign_out(5);
    CN351_data_in(14) <= VN841_data_out(5);
    CN351_sign_in(14) <= VN841_sign_out(5);
    CN351_data_in(15) <= VN933_data_out(5);
    CN351_sign_in(15) <= VN933_sign_out(5);
    CN351_data_in(16) <= VN974_data_out(5);
    CN351_sign_in(16) <= VN974_sign_out(5);
    CN351_data_in(17) <= VN1004_data_out(5);
    CN351_sign_in(17) <= VN1004_sign_out(5);
    CN351_data_in(18) <= VN1109_data_out(5);
    CN351_sign_in(18) <= VN1109_sign_out(5);
    CN351_data_in(19) <= VN1147_data_out(5);
    CN351_sign_in(19) <= VN1147_sign_out(5);
    CN351_data_in(20) <= VN1191_data_out(5);
    CN351_sign_in(20) <= VN1191_sign_out(5);
    CN351_data_in(21) <= VN1253_data_out(5);
    CN351_sign_in(21) <= VN1253_sign_out(5);
    CN351_data_in(22) <= VN1301_data_out(5);
    CN351_sign_in(22) <= VN1301_sign_out(5);
    CN351_data_in(23) <= VN1395_data_out(5);
    CN351_sign_in(23) <= VN1395_sign_out(5);
    CN351_data_in(24) <= VN1642_data_out(5);
    CN351_sign_in(24) <= VN1642_sign_out(5);
    CN351_data_in(25) <= VN1658_data_out(5);
    CN351_sign_in(25) <= VN1658_sign_out(5);
    CN351_data_in(26) <= VN1703_data_out(5);
    CN351_sign_in(26) <= VN1703_sign_out(5);
    CN351_data_in(27) <= VN1869_data_out(5);
    CN351_sign_in(27) <= VN1869_sign_out(5);
    CN351_data_in(28) <= VN1883_data_out(5);
    CN351_sign_in(28) <= VN1883_sign_out(5);
    CN351_data_in(29) <= VN1996_data_out(5);
    CN351_sign_in(29) <= VN1996_sign_out(5);
    CN351_data_in(30) <= VN2012_data_out(5);
    CN351_sign_in(30) <= VN2012_sign_out(5);
    CN351_data_in(31) <= VN2027_data_out(5);
    CN351_sign_in(31) <= VN2027_sign_out(5);
    CN352_data_in(0) <= VN22_data_out(5);
    CN352_sign_in(0) <= VN22_sign_out(5);
    CN352_data_in(1) <= VN100_data_out(5);
    CN352_sign_in(1) <= VN100_sign_out(5);
    CN352_data_in(2) <= VN141_data_out(5);
    CN352_sign_in(2) <= VN141_sign_out(5);
    CN352_data_in(3) <= VN192_data_out(5);
    CN352_sign_in(3) <= VN192_sign_out(5);
    CN352_data_in(4) <= VN239_data_out(5);
    CN352_sign_in(4) <= VN239_sign_out(5);
    CN352_data_in(5) <= VN321_data_out(5);
    CN352_sign_in(5) <= VN321_sign_out(5);
    CN352_data_in(6) <= VN374_data_out(5);
    CN352_sign_in(6) <= VN374_sign_out(5);
    CN352_data_in(7) <= VN428_data_out(5);
    CN352_sign_in(7) <= VN428_sign_out(5);
    CN352_data_in(8) <= VN485_data_out(5);
    CN352_sign_in(8) <= VN485_sign_out(5);
    CN352_data_in(9) <= VN513_data_out(5);
    CN352_sign_in(9) <= VN513_sign_out(5);
    CN352_data_in(10) <= VN609_data_out(5);
    CN352_sign_in(10) <= VN609_sign_out(5);
    CN352_data_in(11) <= VN642_data_out(5);
    CN352_sign_in(11) <= VN642_sign_out(5);
    CN352_data_in(12) <= VN715_data_out(5);
    CN352_sign_in(12) <= VN715_sign_out(5);
    CN352_data_in(13) <= VN723_data_out(5);
    CN352_sign_in(13) <= VN723_sign_out(5);
    CN352_data_in(14) <= VN783_data_out(5);
    CN352_sign_in(14) <= VN783_sign_out(5);
    CN352_data_in(15) <= VN883_data_out(5);
    CN352_sign_in(15) <= VN883_sign_out(5);
    CN352_data_in(16) <= VN902_data_out(5);
    CN352_sign_in(16) <= VN902_sign_out(5);
    CN352_data_in(17) <= VN1027_data_out(5);
    CN352_sign_in(17) <= VN1027_sign_out(5);
    CN352_data_in(18) <= VN1067_data_out(5);
    CN352_sign_in(18) <= VN1067_sign_out(5);
    CN352_data_in(19) <= VN1120_data_out(5);
    CN352_sign_in(19) <= VN1120_sign_out(5);
    CN352_data_in(20) <= VN1187_data_out(5);
    CN352_sign_in(20) <= VN1187_sign_out(5);
    CN352_data_in(21) <= VN1266_data_out(5);
    CN352_sign_in(21) <= VN1266_sign_out(5);
    CN352_data_in(22) <= VN1295_data_out(5);
    CN352_sign_in(22) <= VN1295_sign_out(5);
    CN352_data_in(23) <= VN1333_data_out(5);
    CN352_sign_in(23) <= VN1333_sign_out(5);
    CN352_data_in(24) <= VN1365_data_out(5);
    CN352_sign_in(24) <= VN1365_sign_out(5);
    CN352_data_in(25) <= VN1550_data_out(5);
    CN352_sign_in(25) <= VN1550_sign_out(5);
    CN352_data_in(26) <= VN1610_data_out(5);
    CN352_sign_in(26) <= VN1610_sign_out(5);
    CN352_data_in(27) <= VN1687_data_out(5);
    CN352_sign_in(27) <= VN1687_sign_out(5);
    CN352_data_in(28) <= VN1754_data_out(5);
    CN352_sign_in(28) <= VN1754_sign_out(5);
    CN352_data_in(29) <= VN1784_data_out(5);
    CN352_sign_in(29) <= VN1784_sign_out(5);
    CN352_data_in(30) <= VN1843_data_out(5);
    CN352_sign_in(30) <= VN1843_sign_out(5);
    CN352_data_in(31) <= VN1902_data_out(5);
    CN352_sign_in(31) <= VN1902_sign_out(5);
    CN353_data_in(0) <= VN21_data_out(5);
    CN353_sign_in(0) <= VN21_sign_out(5);
    CN353_data_in(1) <= VN74_data_out(5);
    CN353_sign_in(1) <= VN74_sign_out(5);
    CN353_data_in(2) <= VN160_data_out(5);
    CN353_sign_in(2) <= VN160_sign_out(5);
    CN353_data_in(3) <= VN224_data_out(5);
    CN353_sign_in(3) <= VN224_sign_out(5);
    CN353_data_in(4) <= VN227_data_out(5);
    CN353_sign_in(4) <= VN227_sign_out(5);
    CN353_data_in(5) <= VN336_data_out(5);
    CN353_sign_in(5) <= VN336_sign_out(5);
    CN353_data_in(6) <= VN409_data_out(5);
    CN353_sign_in(6) <= VN409_sign_out(5);
    CN353_data_in(7) <= VN467_data_out(5);
    CN353_sign_in(7) <= VN467_sign_out(5);
    CN353_data_in(8) <= VN541_data_out(5);
    CN353_sign_in(8) <= VN541_sign_out(5);
    CN353_data_in(9) <= VN643_data_out(5);
    CN353_sign_in(9) <= VN643_sign_out(5);
    CN353_data_in(10) <= VN694_data_out(5);
    CN353_sign_in(10) <= VN694_sign_out(5);
    CN353_data_in(11) <= VN762_data_out(5);
    CN353_sign_in(11) <= VN762_sign_out(5);
    CN353_data_in(12) <= VN786_data_out(5);
    CN353_sign_in(12) <= VN786_sign_out(5);
    CN353_data_in(13) <= VN844_data_out(5);
    CN353_sign_in(13) <= VN844_sign_out(5);
    CN353_data_in(14) <= VN915_data_out(5);
    CN353_sign_in(14) <= VN915_sign_out(5);
    CN353_data_in(15) <= VN1009_data_out(5);
    CN353_sign_in(15) <= VN1009_sign_out(5);
    CN353_data_in(16) <= VN1134_data_out(5);
    CN353_sign_in(16) <= VN1134_sign_out(5);
    CN353_data_in(17) <= VN1205_data_out(5);
    CN353_sign_in(17) <= VN1205_sign_out(5);
    CN353_data_in(18) <= VN1262_data_out(5);
    CN353_sign_in(18) <= VN1262_sign_out(5);
    CN353_data_in(19) <= VN1323_data_out(5);
    CN353_sign_in(19) <= VN1323_sign_out(5);
    CN353_data_in(20) <= VN1404_data_out(5);
    CN353_sign_in(20) <= VN1404_sign_out(5);
    CN353_data_in(21) <= VN1472_data_out(5);
    CN353_sign_in(21) <= VN1472_sign_out(5);
    CN353_data_in(22) <= VN1576_data_out(5);
    CN353_sign_in(22) <= VN1576_sign_out(5);
    CN353_data_in(23) <= VN1618_data_out(5);
    CN353_sign_in(23) <= VN1618_sign_out(5);
    CN353_data_in(24) <= VN1780_data_out(5);
    CN353_sign_in(24) <= VN1780_sign_out(5);
    CN353_data_in(25) <= VN1791_data_out(5);
    CN353_sign_in(25) <= VN1791_sign_out(5);
    CN353_data_in(26) <= VN1871_data_out(5);
    CN353_sign_in(26) <= VN1871_sign_out(5);
    CN353_data_in(27) <= VN1881_data_out(5);
    CN353_sign_in(27) <= VN1881_sign_out(5);
    CN353_data_in(28) <= VN1890_data_out(5);
    CN353_sign_in(28) <= VN1890_sign_out(5);
    CN353_data_in(29) <= VN1894_data_out(5);
    CN353_sign_in(29) <= VN1894_sign_out(5);
    CN353_data_in(30) <= VN2011_data_out(5);
    CN353_sign_in(30) <= VN2011_sign_out(5);
    CN353_data_in(31) <= VN2028_data_out(5);
    CN353_sign_in(31) <= VN2028_sign_out(5);
    CN354_data_in(0) <= VN20_data_out(5);
    CN354_sign_in(0) <= VN20_sign_out(5);
    CN354_data_in(1) <= VN88_data_out(5);
    CN354_sign_in(1) <= VN88_sign_out(5);
    CN354_data_in(2) <= VN133_data_out(5);
    CN354_sign_in(2) <= VN133_sign_out(5);
    CN354_data_in(3) <= VN191_data_out(5);
    CN354_sign_in(3) <= VN191_sign_out(5);
    CN354_data_in(4) <= VN326_data_out(5);
    CN354_sign_in(4) <= VN326_sign_out(5);
    CN354_data_in(5) <= VN364_data_out(5);
    CN354_sign_in(5) <= VN364_sign_out(5);
    CN354_data_in(6) <= VN417_data_out(5);
    CN354_sign_in(6) <= VN417_sign_out(5);
    CN354_data_in(7) <= VN470_data_out(5);
    CN354_sign_in(7) <= VN470_sign_out(5);
    CN354_data_in(8) <= VN576_data_out(5);
    CN354_sign_in(8) <= VN576_sign_out(5);
    CN354_data_in(9) <= VN621_data_out(5);
    CN354_sign_in(9) <= VN621_sign_out(5);
    CN354_data_in(10) <= VN773_data_out(5);
    CN354_sign_in(10) <= VN773_sign_out(5);
    CN354_data_in(11) <= VN864_data_out(5);
    CN354_sign_in(11) <= VN864_sign_out(5);
    CN354_data_in(12) <= VN912_data_out(5);
    CN354_sign_in(12) <= VN912_sign_out(5);
    CN354_data_in(13) <= VN965_data_out(5);
    CN354_sign_in(13) <= VN965_sign_out(5);
    CN354_data_in(14) <= VN1064_data_out(5);
    CN354_sign_in(14) <= VN1064_sign_out(5);
    CN354_data_in(15) <= VN1108_data_out(5);
    CN354_sign_in(15) <= VN1108_sign_out(5);
    CN354_data_in(16) <= VN1172_data_out(5);
    CN354_sign_in(16) <= VN1172_sign_out(5);
    CN354_data_in(17) <= VN1226_data_out(5);
    CN354_sign_in(17) <= VN1226_sign_out(5);
    CN354_data_in(18) <= VN1371_data_out(5);
    CN354_sign_in(18) <= VN1371_sign_out(5);
    CN354_data_in(19) <= VN1409_data_out(5);
    CN354_sign_in(19) <= VN1409_sign_out(5);
    CN354_data_in(20) <= VN1440_data_out(5);
    CN354_sign_in(20) <= VN1440_sign_out(5);
    CN354_data_in(21) <= VN1478_data_out(5);
    CN354_sign_in(21) <= VN1478_sign_out(5);
    CN354_data_in(22) <= VN1531_data_out(5);
    CN354_sign_in(22) <= VN1531_sign_out(5);
    CN354_data_in(23) <= VN1707_data_out(5);
    CN354_sign_in(23) <= VN1707_sign_out(5);
    CN354_data_in(24) <= VN1738_data_out(5);
    CN354_sign_in(24) <= VN1738_sign_out(5);
    CN354_data_in(25) <= VN1817_data_out(5);
    CN354_sign_in(25) <= VN1817_sign_out(5);
    CN354_data_in(26) <= VN1877_data_out(5);
    CN354_sign_in(26) <= VN1877_sign_out(5);
    CN354_data_in(27) <= VN1892_data_out(5);
    CN354_sign_in(27) <= VN1892_sign_out(5);
    CN354_data_in(28) <= VN1921_data_out(5);
    CN354_sign_in(28) <= VN1921_sign_out(5);
    CN354_data_in(29) <= VN1973_data_out(5);
    CN354_sign_in(29) <= VN1973_sign_out(5);
    CN354_data_in(30) <= VN2002_data_out(5);
    CN354_sign_in(30) <= VN2002_sign_out(5);
    CN354_data_in(31) <= VN2015_data_out(5);
    CN354_sign_in(31) <= VN2015_sign_out(5);
    CN355_data_in(0) <= VN19_data_out(5);
    CN355_sign_in(0) <= VN19_sign_out(5);
    CN355_data_in(1) <= VN59_data_out(5);
    CN355_sign_in(1) <= VN59_sign_out(5);
    CN355_data_in(2) <= VN130_data_out(5);
    CN355_sign_in(2) <= VN130_sign_out(5);
    CN355_data_in(3) <= VN186_data_out(5);
    CN355_sign_in(3) <= VN186_sign_out(5);
    CN355_data_in(4) <= VN230_data_out(5);
    CN355_sign_in(4) <= VN230_sign_out(5);
    CN355_data_in(5) <= VN300_data_out(5);
    CN355_sign_in(5) <= VN300_sign_out(5);
    CN355_data_in(6) <= VN349_data_out(5);
    CN355_sign_in(6) <= VN349_sign_out(5);
    CN355_data_in(7) <= VN456_data_out(5);
    CN355_sign_in(7) <= VN456_sign_out(5);
    CN355_data_in(8) <= VN543_data_out(5);
    CN355_sign_in(8) <= VN543_sign_out(5);
    CN355_data_in(9) <= VN667_data_out(5);
    CN355_sign_in(9) <= VN667_sign_out(5);
    CN355_data_in(10) <= VN675_data_out(5);
    CN355_sign_in(10) <= VN675_sign_out(5);
    CN355_data_in(11) <= VN729_data_out(5);
    CN355_sign_in(11) <= VN729_sign_out(5);
    CN355_data_in(12) <= VN810_data_out(5);
    CN355_sign_in(12) <= VN810_sign_out(5);
    CN355_data_in(13) <= VN871_data_out(5);
    CN355_sign_in(13) <= VN871_sign_out(5);
    CN355_data_in(14) <= VN930_data_out(5);
    CN355_sign_in(14) <= VN930_sign_out(5);
    CN355_data_in(15) <= VN1028_data_out(5);
    CN355_sign_in(15) <= VN1028_sign_out(5);
    CN355_data_in(16) <= VN1106_data_out(5);
    CN355_sign_in(16) <= VN1106_sign_out(5);
    CN355_data_in(17) <= VN1141_data_out(5);
    CN355_sign_in(17) <= VN1141_sign_out(5);
    CN355_data_in(18) <= VN1173_data_out(5);
    CN355_sign_in(18) <= VN1173_sign_out(5);
    CN355_data_in(19) <= VN1246_data_out(5);
    CN355_sign_in(19) <= VN1246_sign_out(5);
    CN355_data_in(20) <= VN1327_data_out(5);
    CN355_sign_in(20) <= VN1327_sign_out(5);
    CN355_data_in(21) <= VN1383_data_out(5);
    CN355_sign_in(21) <= VN1383_sign_out(5);
    CN355_data_in(22) <= VN1482_data_out(5);
    CN355_sign_in(22) <= VN1482_sign_out(5);
    CN355_data_in(23) <= VN1552_data_out(5);
    CN355_sign_in(23) <= VN1552_sign_out(5);
    CN355_data_in(24) <= VN1557_data_out(5);
    CN355_sign_in(24) <= VN1557_sign_out(5);
    CN355_data_in(25) <= VN1619_data_out(5);
    CN355_sign_in(25) <= VN1619_sign_out(5);
    CN355_data_in(26) <= VN1681_data_out(5);
    CN355_sign_in(26) <= VN1681_sign_out(5);
    CN355_data_in(27) <= VN1847_data_out(5);
    CN355_sign_in(27) <= VN1847_sign_out(5);
    CN355_data_in(28) <= VN1990_data_out(5);
    CN355_sign_in(28) <= VN1990_sign_out(5);
    CN355_data_in(29) <= VN2000_data_out(5);
    CN355_sign_in(29) <= VN2000_sign_out(5);
    CN355_data_in(30) <= VN2001_data_out(5);
    CN355_sign_in(30) <= VN2001_sign_out(5);
    CN355_data_in(31) <= VN2016_data_out(5);
    CN355_sign_in(31) <= VN2016_sign_out(5);
    CN356_data_in(0) <= VN18_data_out(5);
    CN356_sign_in(0) <= VN18_sign_out(5);
    CN356_data_in(1) <= VN95_data_out(5);
    CN356_sign_in(1) <= VN95_sign_out(5);
    CN356_data_in(2) <= VN146_data_out(5);
    CN356_sign_in(2) <= VN146_sign_out(5);
    CN356_data_in(3) <= VN222_data_out(5);
    CN356_sign_in(3) <= VN222_sign_out(5);
    CN356_data_in(4) <= VN299_data_out(5);
    CN356_sign_in(4) <= VN299_sign_out(5);
    CN356_data_in(5) <= VN376_data_out(5);
    CN356_sign_in(5) <= VN376_sign_out(5);
    CN356_data_in(6) <= VN438_data_out(5);
    CN356_sign_in(6) <= VN438_sign_out(5);
    CN356_data_in(7) <= VN486_data_out(5);
    CN356_sign_in(7) <= VN486_sign_out(5);
    CN356_data_in(8) <= VN557_data_out(5);
    CN356_sign_in(8) <= VN557_sign_out(5);
    CN356_data_in(9) <= VN589_data_out(5);
    CN356_sign_in(9) <= VN589_sign_out(5);
    CN356_data_in(10) <= VN672_data_out(5);
    CN356_sign_in(10) <= VN672_sign_out(5);
    CN356_data_in(11) <= VN756_data_out(5);
    CN356_sign_in(11) <= VN756_sign_out(5);
    CN356_data_in(12) <= VN795_data_out(5);
    CN356_sign_in(12) <= VN795_sign_out(5);
    CN356_data_in(13) <= VN895_data_out(5);
    CN356_sign_in(13) <= VN895_sign_out(5);
    CN356_data_in(14) <= VN972_data_out(5);
    CN356_sign_in(14) <= VN972_sign_out(5);
    CN356_data_in(15) <= VN1088_data_out(5);
    CN356_sign_in(15) <= VN1088_sign_out(5);
    CN356_data_in(16) <= VN1204_data_out(5);
    CN356_sign_in(16) <= VN1204_sign_out(5);
    CN356_data_in(17) <= VN1247_data_out(5);
    CN356_sign_in(17) <= VN1247_sign_out(5);
    CN356_data_in(18) <= VN1408_data_out(5);
    CN356_sign_in(18) <= VN1408_sign_out(5);
    CN356_data_in(19) <= VN1464_data_out(5);
    CN356_sign_in(19) <= VN1464_sign_out(5);
    CN356_data_in(20) <= VN1495_data_out(5);
    CN356_sign_in(20) <= VN1495_sign_out(5);
    CN356_data_in(21) <= VN1504_data_out(5);
    CN356_sign_in(21) <= VN1504_sign_out(5);
    CN356_data_in(22) <= VN1511_data_out(5);
    CN356_sign_in(22) <= VN1511_sign_out(5);
    CN356_data_in(23) <= VN1528_data_out(5);
    CN356_sign_in(23) <= VN1528_sign_out(5);
    CN356_data_in(24) <= VN1567_data_out(5);
    CN356_sign_in(24) <= VN1567_sign_out(5);
    CN356_data_in(25) <= VN1609_data_out(5);
    CN356_sign_in(25) <= VN1609_sign_out(5);
    CN356_data_in(26) <= VN1736_data_out(5);
    CN356_sign_in(26) <= VN1736_sign_out(5);
    CN356_data_in(27) <= VN1794_data_out(5);
    CN356_sign_in(27) <= VN1794_sign_out(5);
    CN356_data_in(28) <= VN1893_data_out(5);
    CN356_sign_in(28) <= VN1893_sign_out(5);
    CN356_data_in(29) <= VN1931_data_out(5);
    CN356_sign_in(29) <= VN1931_sign_out(5);
    CN356_data_in(30) <= VN2005_data_out(5);
    CN356_sign_in(30) <= VN2005_sign_out(5);
    CN356_data_in(31) <= VN2006_data_out(5);
    CN356_sign_in(31) <= VN2006_sign_out(5);
    CN357_data_in(0) <= VN17_data_out(5);
    CN357_sign_in(0) <= VN17_sign_out(5);
    CN357_data_in(1) <= VN61_data_out(5);
    CN357_sign_in(1) <= VN61_sign_out(5);
    CN357_data_in(2) <= VN138_data_out(5);
    CN357_sign_in(2) <= VN138_sign_out(5);
    CN357_data_in(3) <= VN176_data_out(5);
    CN357_sign_in(3) <= VN176_sign_out(5);
    CN357_data_in(4) <= VN256_data_out(5);
    CN357_sign_in(4) <= VN256_sign_out(5);
    CN357_data_in(5) <= VN312_data_out(5);
    CN357_sign_in(5) <= VN312_sign_out(5);
    CN357_data_in(6) <= VN366_data_out(5);
    CN357_sign_in(6) <= VN366_sign_out(5);
    CN357_data_in(7) <= VN415_data_out(5);
    CN357_sign_in(7) <= VN415_sign_out(5);
    CN357_data_in(8) <= VN452_data_out(5);
    CN357_sign_in(8) <= VN452_sign_out(5);
    CN357_data_in(9) <= VN632_data_out(5);
    CN357_sign_in(9) <= VN632_sign_out(5);
    CN357_data_in(10) <= VN872_data_out(5);
    CN357_sign_in(10) <= VN872_sign_out(5);
    CN357_data_in(11) <= VN896_data_out(5);
    CN357_sign_in(11) <= VN896_sign_out(5);
    CN357_data_in(12) <= VN984_data_out(5);
    CN357_sign_in(12) <= VN984_sign_out(5);
    CN357_data_in(13) <= VN1016_data_out(5);
    CN357_sign_in(13) <= VN1016_sign_out(5);
    CN357_data_in(14) <= VN1073_data_out(5);
    CN357_sign_in(14) <= VN1073_sign_out(5);
    CN357_data_in(15) <= VN1196_data_out(5);
    CN357_sign_in(15) <= VN1196_sign_out(5);
    CN357_data_in(16) <= VN1225_data_out(5);
    CN357_sign_in(16) <= VN1225_sign_out(5);
    CN357_data_in(17) <= VN1320_data_out(5);
    CN357_sign_in(17) <= VN1320_sign_out(5);
    CN357_data_in(18) <= VN1364_data_out(5);
    CN357_sign_in(18) <= VN1364_sign_out(5);
    CN357_data_in(19) <= VN1402_data_out(5);
    CN357_sign_in(19) <= VN1402_sign_out(5);
    CN357_data_in(20) <= VN1444_data_out(5);
    CN357_sign_in(20) <= VN1444_sign_out(5);
    CN357_data_in(21) <= VN1575_data_out(5);
    CN357_sign_in(21) <= VN1575_sign_out(5);
    CN357_data_in(22) <= VN1593_data_out(5);
    CN357_sign_in(22) <= VN1593_sign_out(5);
    CN357_data_in(23) <= VN1760_data_out(5);
    CN357_sign_in(23) <= VN1760_sign_out(5);
    CN357_data_in(24) <= VN1792_data_out(5);
    CN357_sign_in(24) <= VN1792_sign_out(5);
    CN357_data_in(25) <= VN1830_data_out(5);
    CN357_sign_in(25) <= VN1830_sign_out(5);
    CN357_data_in(26) <= VN1876_data_out(5);
    CN357_sign_in(26) <= VN1876_sign_out(5);
    CN357_data_in(27) <= VN1962_data_out(5);
    CN357_sign_in(27) <= VN1962_sign_out(5);
    CN357_data_in(28) <= VN1975_data_out(5);
    CN357_sign_in(28) <= VN1975_sign_out(5);
    CN357_data_in(29) <= VN2025_data_out(5);
    CN357_sign_in(29) <= VN2025_sign_out(5);
    CN357_data_in(30) <= VN2032_data_out(5);
    CN357_sign_in(30) <= VN2032_sign_out(5);
    CN357_data_in(31) <= VN2041_data_out(5);
    CN357_sign_in(31) <= VN2041_sign_out(5);
    CN358_data_in(0) <= VN16_data_out(5);
    CN358_sign_in(0) <= VN16_sign_out(5);
    CN358_data_in(1) <= VN76_data_out(5);
    CN358_sign_in(1) <= VN76_sign_out(5);
    CN358_data_in(2) <= VN112_data_out(5);
    CN358_sign_in(2) <= VN112_sign_out(5);
    CN358_data_in(3) <= VN252_data_out(5);
    CN358_sign_in(3) <= VN252_sign_out(5);
    CN358_data_in(4) <= VN305_data_out(5);
    CN358_sign_in(4) <= VN305_sign_out(5);
    CN358_data_in(5) <= VN353_data_out(5);
    CN358_sign_in(5) <= VN353_sign_out(5);
    CN358_data_in(6) <= VN396_data_out(5);
    CN358_sign_in(6) <= VN396_sign_out(5);
    CN358_data_in(7) <= VN478_data_out(5);
    CN358_sign_in(7) <= VN478_sign_out(5);
    CN358_data_in(8) <= VN515_data_out(5);
    CN358_sign_in(8) <= VN515_sign_out(5);
    CN358_data_in(9) <= VN578_data_out(5);
    CN358_sign_in(9) <= VN578_sign_out(5);
    CN358_data_in(10) <= VN668_data_out(5);
    CN358_sign_in(10) <= VN668_sign_out(5);
    CN358_data_in(11) <= VN711_data_out(5);
    CN358_sign_in(11) <= VN711_sign_out(5);
    CN358_data_in(12) <= VN731_data_out(5);
    CN358_sign_in(12) <= VN731_sign_out(5);
    CN358_data_in(13) <= VN817_data_out(5);
    CN358_sign_in(13) <= VN817_sign_out(5);
    CN358_data_in(14) <= VN863_data_out(5);
    CN358_sign_in(14) <= VN863_sign_out(5);
    CN358_data_in(15) <= VN929_data_out(5);
    CN358_sign_in(15) <= VN929_sign_out(5);
    CN358_data_in(16) <= VN992_data_out(5);
    CN358_sign_in(16) <= VN992_sign_out(5);
    CN358_data_in(17) <= VN1044_data_out(5);
    CN358_sign_in(17) <= VN1044_sign_out(5);
    CN358_data_in(18) <= VN1084_data_out(5);
    CN358_sign_in(18) <= VN1084_sign_out(5);
    CN358_data_in(19) <= VN1118_data_out(5);
    CN358_sign_in(19) <= VN1118_sign_out(5);
    CN358_data_in(20) <= VN1213_data_out(5);
    CN358_sign_in(20) <= VN1213_sign_out(5);
    CN358_data_in(21) <= VN1273_data_out(5);
    CN358_sign_in(21) <= VN1273_sign_out(5);
    CN358_data_in(22) <= VN1378_data_out(5);
    CN358_sign_in(22) <= VN1378_sign_out(5);
    CN358_data_in(23) <= VN1447_data_out(5);
    CN358_sign_in(23) <= VN1447_sign_out(5);
    CN358_data_in(24) <= VN1566_data_out(5);
    CN358_sign_in(24) <= VN1566_sign_out(5);
    CN358_data_in(25) <= VN1581_data_out(5);
    CN358_sign_in(25) <= VN1581_sign_out(5);
    CN358_data_in(26) <= VN1733_data_out(5);
    CN358_sign_in(26) <= VN1733_sign_out(5);
    CN358_data_in(27) <= VN1812_data_out(5);
    CN358_sign_in(27) <= VN1812_sign_out(5);
    CN358_data_in(28) <= VN1866_data_out(5);
    CN358_sign_in(28) <= VN1866_sign_out(5);
    CN358_data_in(29) <= VN1932_data_out(5);
    CN358_sign_in(29) <= VN1932_sign_out(5);
    CN358_data_in(30) <= VN1944_data_out(5);
    CN358_sign_in(30) <= VN1944_sign_out(5);
    CN358_data_in(31) <= VN1959_data_out(5);
    CN358_sign_in(31) <= VN1959_sign_out(5);
    CN359_data_in(0) <= VN15_data_out(5);
    CN359_sign_in(0) <= VN15_sign_out(5);
    CN359_data_in(1) <= VN72_data_out(5);
    CN359_sign_in(1) <= VN72_sign_out(5);
    CN359_data_in(2) <= VN122_data_out(5);
    CN359_sign_in(2) <= VN122_sign_out(5);
    CN359_data_in(3) <= VN195_data_out(5);
    CN359_sign_in(3) <= VN195_sign_out(5);
    CN359_data_in(4) <= VN257_data_out(5);
    CN359_sign_in(4) <= VN257_sign_out(5);
    CN359_data_in(5) <= VN283_data_out(5);
    CN359_sign_in(5) <= VN283_sign_out(5);
    CN359_data_in(6) <= VN372_data_out(5);
    CN359_sign_in(6) <= VN372_sign_out(5);
    CN359_data_in(7) <= VN399_data_out(5);
    CN359_sign_in(7) <= VN399_sign_out(5);
    CN359_data_in(8) <= VN464_data_out(5);
    CN359_sign_in(8) <= VN464_sign_out(5);
    CN359_data_in(9) <= VN536_data_out(5);
    CN359_sign_in(9) <= VN536_sign_out(5);
    CN359_data_in(10) <= VN608_data_out(5);
    CN359_sign_in(10) <= VN608_sign_out(5);
    CN359_data_in(11) <= VN631_data_out(5);
    CN359_sign_in(11) <= VN631_sign_out(5);
    CN359_data_in(12) <= VN712_data_out(5);
    CN359_sign_in(12) <= VN712_sign_out(5);
    CN359_data_in(13) <= VN747_data_out(5);
    CN359_sign_in(13) <= VN747_sign_out(5);
    CN359_data_in(14) <= VN790_data_out(5);
    CN359_sign_in(14) <= VN790_sign_out(5);
    CN359_data_in(15) <= VN886_data_out(5);
    CN359_sign_in(15) <= VN886_sign_out(5);
    CN359_data_in(16) <= VN964_data_out(5);
    CN359_sign_in(16) <= VN964_sign_out(5);
    CN359_data_in(17) <= VN1023_data_out(5);
    CN359_sign_in(17) <= VN1023_sign_out(5);
    CN359_data_in(18) <= VN1093_data_out(5);
    CN359_sign_in(18) <= VN1093_sign_out(5);
    CN359_data_in(19) <= VN1137_data_out(5);
    CN359_sign_in(19) <= VN1137_sign_out(5);
    CN359_data_in(20) <= VN1216_data_out(5);
    CN359_sign_in(20) <= VN1216_sign_out(5);
    CN359_data_in(21) <= VN1286_data_out(5);
    CN359_sign_in(21) <= VN1286_sign_out(5);
    CN359_data_in(22) <= VN1352_data_out(5);
    CN359_sign_in(22) <= VN1352_sign_out(5);
    CN359_data_in(23) <= VN1561_data_out(5);
    CN359_sign_in(23) <= VN1561_sign_out(5);
    CN359_data_in(24) <= VN1591_data_out(5);
    CN359_sign_in(24) <= VN1591_sign_out(5);
    CN359_data_in(25) <= VN1623_data_out(5);
    CN359_sign_in(25) <= VN1623_sign_out(5);
    CN359_data_in(26) <= VN1685_data_out(5);
    CN359_sign_in(26) <= VN1685_sign_out(5);
    CN359_data_in(27) <= VN1743_data_out(5);
    CN359_sign_in(27) <= VN1743_sign_out(5);
    CN359_data_in(28) <= VN1771_data_out(5);
    CN359_sign_in(28) <= VN1771_sign_out(5);
    CN359_data_in(29) <= VN1834_data_out(5);
    CN359_sign_in(29) <= VN1834_sign_out(5);
    CN359_data_in(30) <= VN1920_data_out(5);
    CN359_sign_in(30) <= VN1920_sign_out(5);
    CN359_data_in(31) <= VN1924_data_out(5);
    CN359_sign_in(31) <= VN1924_sign_out(5);
    CN360_data_in(0) <= VN14_data_out(5);
    CN360_sign_in(0) <= VN14_sign_out(5);
    CN360_data_in(1) <= VN91_data_out(5);
    CN360_sign_in(1) <= VN91_sign_out(5);
    CN360_data_in(2) <= VN116_data_out(5);
    CN360_sign_in(2) <= VN116_sign_out(5);
    CN360_data_in(3) <= VN174_data_out(5);
    CN360_sign_in(3) <= VN174_sign_out(5);
    CN360_data_in(4) <= VN248_data_out(5);
    CN360_sign_in(4) <= VN248_sign_out(5);
    CN360_data_in(5) <= VN292_data_out(5);
    CN360_sign_in(5) <= VN292_sign_out(5);
    CN360_data_in(6) <= VN345_data_out(5);
    CN360_sign_in(6) <= VN345_sign_out(5);
    CN360_data_in(7) <= VN440_data_out(5);
    CN360_sign_in(7) <= VN440_sign_out(5);
    CN360_data_in(8) <= VN488_data_out(5);
    CN360_sign_in(8) <= VN488_sign_out(5);
    CN360_data_in(9) <= VN537_data_out(5);
    CN360_sign_in(9) <= VN537_sign_out(5);
    CN360_data_in(10) <= VN575_data_out(5);
    CN360_sign_in(10) <= VN575_sign_out(5);
    CN360_data_in(11) <= VN627_data_out(5);
    CN360_sign_in(11) <= VN627_sign_out(5);
    CN360_data_in(12) <= VN689_data_out(5);
    CN360_sign_in(12) <= VN689_sign_out(5);
    CN360_data_in(13) <= VN767_data_out(5);
    CN360_sign_in(13) <= VN767_sign_out(5);
    CN360_data_in(14) <= VN779_data_out(5);
    CN360_sign_in(14) <= VN779_sign_out(5);
    CN360_data_in(15) <= VN836_data_out(5);
    CN360_sign_in(15) <= VN836_sign_out(5);
    CN360_data_in(16) <= VN937_data_out(5);
    CN360_sign_in(16) <= VN937_sign_out(5);
    CN360_data_in(17) <= VN980_data_out(5);
    CN360_sign_in(17) <= VN980_sign_out(5);
    CN360_data_in(18) <= VN1046_data_out(5);
    CN360_sign_in(18) <= VN1046_sign_out(5);
    CN360_data_in(19) <= VN1068_data_out(5);
    CN360_sign_in(19) <= VN1068_sign_out(5);
    CN360_data_in(20) <= VN1159_data_out(5);
    CN360_sign_in(20) <= VN1159_sign_out(5);
    CN360_data_in(21) <= VN1168_data_out(5);
    CN360_sign_in(21) <= VN1168_sign_out(5);
    CN360_data_in(22) <= VN1239_data_out(5);
    CN360_sign_in(22) <= VN1239_sign_out(5);
    CN360_data_in(23) <= VN1298_data_out(5);
    CN360_sign_in(23) <= VN1298_sign_out(5);
    CN360_data_in(24) <= VN1414_data_out(5);
    CN360_sign_in(24) <= VN1414_sign_out(5);
    CN360_data_in(25) <= VN1438_data_out(5);
    CN360_sign_in(25) <= VN1438_sign_out(5);
    CN360_data_in(26) <= VN1519_data_out(5);
    CN360_sign_in(26) <= VN1519_sign_out(5);
    CN360_data_in(27) <= VN1534_data_out(5);
    CN360_sign_in(27) <= VN1534_sign_out(5);
    CN360_data_in(28) <= VN1599_data_out(5);
    CN360_sign_in(28) <= VN1599_sign_out(5);
    CN360_data_in(29) <= VN1625_data_out(5);
    CN360_sign_in(29) <= VN1625_sign_out(5);
    CN360_data_in(30) <= VN1698_data_out(5);
    CN360_sign_in(30) <= VN1698_sign_out(5);
    CN360_data_in(31) <= VN1807_data_out(5);
    CN360_sign_in(31) <= VN1807_sign_out(5);
    CN361_data_in(0) <= VN13_data_out(5);
    CN361_sign_in(0) <= VN13_sign_out(5);
    CN361_data_in(1) <= VN54_data_out(5);
    CN361_sign_in(1) <= VN54_sign_out(5);
    CN361_data_in(2) <= VN120_data_out(5);
    CN361_sign_in(2) <= VN120_sign_out(5);
    CN361_data_in(3) <= VN207_data_out(5);
    CN361_sign_in(3) <= VN207_sign_out(5);
    CN361_data_in(4) <= VN271_data_out(5);
    CN361_sign_in(4) <= VN271_sign_out(5);
    CN361_data_in(5) <= VN285_data_out(5);
    CN361_sign_in(5) <= VN285_sign_out(5);
    CN361_data_in(6) <= VN342_data_out(5);
    CN361_sign_in(6) <= VN342_sign_out(5);
    CN361_data_in(7) <= VN391_data_out(5);
    CN361_sign_in(7) <= VN391_sign_out(5);
    CN361_data_in(8) <= VN416_data_out(5);
    CN361_sign_in(8) <= VN416_sign_out(5);
    CN361_data_in(9) <= VN480_data_out(5);
    CN361_sign_in(9) <= VN480_sign_out(5);
    CN361_data_in(10) <= VN601_data_out(5);
    CN361_sign_in(10) <= VN601_sign_out(5);
    CN361_data_in(11) <= VN664_data_out(5);
    CN361_sign_in(11) <= VN664_sign_out(5);
    CN361_data_in(12) <= VN775_data_out(5);
    CN361_sign_in(12) <= VN775_sign_out(5);
    CN361_data_in(13) <= VN876_data_out(5);
    CN361_sign_in(13) <= VN876_sign_out(5);
    CN361_data_in(14) <= VN942_data_out(5);
    CN361_sign_in(14) <= VN942_sign_out(5);
    CN361_data_in(15) <= VN950_data_out(5);
    CN361_sign_in(15) <= VN950_sign_out(5);
    CN361_data_in(16) <= VN1005_data_out(5);
    CN361_sign_in(16) <= VN1005_sign_out(5);
    CN361_data_in(17) <= VN1160_data_out(5);
    CN361_sign_in(17) <= VN1160_sign_out(5);
    CN361_data_in(18) <= VN1215_data_out(5);
    CN361_sign_in(18) <= VN1215_sign_out(5);
    CN361_data_in(19) <= VN1306_data_out(5);
    CN361_sign_in(19) <= VN1306_sign_out(5);
    CN361_data_in(20) <= VN1354_data_out(5);
    CN361_sign_in(20) <= VN1354_sign_out(5);
    CN361_data_in(21) <= VN1412_data_out(5);
    CN361_sign_in(21) <= VN1412_sign_out(5);
    CN361_data_in(22) <= VN1468_data_out(5);
    CN361_sign_in(22) <= VN1468_sign_out(5);
    CN361_data_in(23) <= VN1487_data_out(5);
    CN361_sign_in(23) <= VN1487_sign_out(5);
    CN361_data_in(24) <= VN1506_data_out(5);
    CN361_sign_in(24) <= VN1506_sign_out(5);
    CN361_data_in(25) <= VN1525_data_out(5);
    CN361_sign_in(25) <= VN1525_sign_out(5);
    CN361_data_in(26) <= VN1645_data_out(5);
    CN361_sign_in(26) <= VN1645_sign_out(5);
    CN361_data_in(27) <= VN1774_data_out(5);
    CN361_sign_in(27) <= VN1774_sign_out(5);
    CN361_data_in(28) <= VN1811_data_out(5);
    CN361_sign_in(28) <= VN1811_sign_out(5);
    CN361_data_in(29) <= VN1915_data_out(5);
    CN361_sign_in(29) <= VN1915_sign_out(5);
    CN361_data_in(30) <= VN2007_data_out(5);
    CN361_sign_in(30) <= VN2007_sign_out(5);
    CN361_data_in(31) <= VN2009_data_out(5);
    CN361_sign_in(31) <= VN2009_sign_out(5);
    CN362_data_in(0) <= VN12_data_out(5);
    CN362_sign_in(0) <= VN12_sign_out(5);
    CN362_data_in(1) <= VN55_data_out(5);
    CN362_sign_in(1) <= VN55_sign_out(5);
    CN362_data_in(2) <= VN169_data_out(5);
    CN362_sign_in(2) <= VN169_sign_out(5);
    CN362_data_in(3) <= VN210_data_out(5);
    CN362_sign_in(3) <= VN210_sign_out(5);
    CN362_data_in(4) <= VN276_data_out(5);
    CN362_sign_in(4) <= VN276_sign_out(5);
    CN362_data_in(5) <= VN289_data_out(5);
    CN362_sign_in(5) <= VN289_sign_out(5);
    CN362_data_in(6) <= VN357_data_out(5);
    CN362_sign_in(6) <= VN357_sign_out(5);
    CN362_data_in(7) <= VN468_data_out(5);
    CN362_sign_in(7) <= VN468_sign_out(5);
    CN362_data_in(8) <= VN586_data_out(5);
    CN362_sign_in(8) <= VN586_sign_out(5);
    CN362_data_in(9) <= VN619_data_out(5);
    CN362_sign_in(9) <= VN619_sign_out(5);
    CN362_data_in(10) <= VN698_data_out(5);
    CN362_sign_in(10) <= VN698_sign_out(5);
    CN362_data_in(11) <= VN771_data_out(5);
    CN362_sign_in(11) <= VN771_sign_out(5);
    CN362_data_in(12) <= VN781_data_out(5);
    CN362_sign_in(12) <= VN781_sign_out(5);
    CN362_data_in(13) <= VN877_data_out(5);
    CN362_sign_in(13) <= VN877_sign_out(5);
    CN362_data_in(14) <= VN987_data_out(5);
    CN362_sign_in(14) <= VN987_sign_out(5);
    CN362_data_in(15) <= VN1057_data_out(5);
    CN362_sign_in(15) <= VN1057_sign_out(5);
    CN362_data_in(16) <= VN1095_data_out(5);
    CN362_sign_in(16) <= VN1095_sign_out(5);
    CN362_data_in(17) <= VN1136_data_out(5);
    CN362_sign_in(17) <= VN1136_sign_out(5);
    CN362_data_in(18) <= VN1164_data_out(5);
    CN362_sign_in(18) <= VN1164_sign_out(5);
    CN362_data_in(19) <= VN1212_data_out(5);
    CN362_sign_in(19) <= VN1212_sign_out(5);
    CN362_data_in(20) <= VN1238_data_out(5);
    CN362_sign_in(20) <= VN1238_sign_out(5);
    CN362_data_in(21) <= VN1283_data_out(5);
    CN362_sign_in(21) <= VN1283_sign_out(5);
    CN362_data_in(22) <= VN1366_data_out(5);
    CN362_sign_in(22) <= VN1366_sign_out(5);
    CN362_data_in(23) <= VN1392_data_out(5);
    CN362_sign_in(23) <= VN1392_sign_out(5);
    CN362_data_in(24) <= VN1466_data_out(5);
    CN362_sign_in(24) <= VN1466_sign_out(5);
    CN362_data_in(25) <= VN1502_data_out(5);
    CN362_sign_in(25) <= VN1502_sign_out(5);
    CN362_data_in(26) <= VN1663_data_out(5);
    CN362_sign_in(26) <= VN1663_sign_out(5);
    CN362_data_in(27) <= VN1731_data_out(5);
    CN362_sign_in(27) <= VN1731_sign_out(5);
    CN362_data_in(28) <= VN1739_data_out(5);
    CN362_sign_in(28) <= VN1739_sign_out(5);
    CN362_data_in(29) <= VN1829_data_out(5);
    CN362_sign_in(29) <= VN1829_sign_out(5);
    CN362_data_in(30) <= VN1995_data_out(5);
    CN362_sign_in(30) <= VN1995_sign_out(5);
    CN362_data_in(31) <= VN1999_data_out(5);
    CN362_sign_in(31) <= VN1999_sign_out(5);
    CN363_data_in(0) <= VN90_data_out(5);
    CN363_sign_in(0) <= VN90_sign_out(5);
    CN363_data_in(1) <= VN147_data_out(5);
    CN363_sign_in(1) <= VN147_sign_out(5);
    CN363_data_in(2) <= VN197_data_out(5);
    CN363_sign_in(2) <= VN197_sign_out(5);
    CN363_data_in(3) <= VN261_data_out(5);
    CN363_sign_in(3) <= VN261_sign_out(5);
    CN363_data_in(4) <= VN281_data_out(5);
    CN363_sign_in(4) <= VN281_sign_out(5);
    CN363_data_in(5) <= VN407_data_out(5);
    CN363_sign_in(5) <= VN407_sign_out(5);
    CN363_data_in(6) <= VN522_data_out(5);
    CN363_sign_in(6) <= VN522_sign_out(5);
    CN363_data_in(7) <= VN610_data_out(5);
    CN363_sign_in(7) <= VN610_sign_out(5);
    CN363_data_in(8) <= VN638_data_out(5);
    CN363_sign_in(8) <= VN638_sign_out(5);
    CN363_data_in(9) <= VN703_data_out(5);
    CN363_sign_in(9) <= VN703_sign_out(5);
    CN363_data_in(10) <= VN848_data_out(5);
    CN363_sign_in(10) <= VN848_sign_out(5);
    CN363_data_in(11) <= VN941_data_out(5);
    CN363_sign_in(11) <= VN941_sign_out(5);
    CN363_data_in(12) <= VN952_data_out(5);
    CN363_sign_in(12) <= VN952_sign_out(5);
    CN363_data_in(13) <= VN1019_data_out(5);
    CN363_sign_in(13) <= VN1019_sign_out(5);
    CN363_data_in(14) <= VN1111_data_out(5);
    CN363_sign_in(14) <= VN1111_sign_out(5);
    CN363_data_in(15) <= VN1128_data_out(5);
    CN363_sign_in(15) <= VN1128_sign_out(5);
    CN363_data_in(16) <= VN1193_data_out(5);
    CN363_sign_in(16) <= VN1193_sign_out(5);
    CN363_data_in(17) <= VN1223_data_out(5);
    CN363_sign_in(17) <= VN1223_sign_out(5);
    CN363_data_in(18) <= VN1233_data_out(5);
    CN363_sign_in(18) <= VN1233_sign_out(5);
    CN363_data_in(19) <= VN1322_data_out(5);
    CN363_sign_in(19) <= VN1322_sign_out(5);
    CN363_data_in(20) <= VN1363_data_out(5);
    CN363_sign_in(20) <= VN1363_sign_out(5);
    CN363_data_in(21) <= VN1571_data_out(5);
    CN363_sign_in(21) <= VN1571_sign_out(5);
    CN363_data_in(22) <= VN1601_data_out(5);
    CN363_sign_in(22) <= VN1601_sign_out(5);
    CN363_data_in(23) <= VN1638_data_out(5);
    CN363_sign_in(23) <= VN1638_sign_out(5);
    CN363_data_in(24) <= VN1686_data_out(5);
    CN363_sign_in(24) <= VN1686_sign_out(5);
    CN363_data_in(25) <= VN1785_data_out(5);
    CN363_sign_in(25) <= VN1785_sign_out(5);
    CN363_data_in(26) <= VN1821_data_out(5);
    CN363_sign_in(26) <= VN1821_sign_out(5);
    CN363_data_in(27) <= VN1858_data_out(5);
    CN363_sign_in(27) <= VN1858_sign_out(5);
    CN363_data_in(28) <= VN1889_data_out(5);
    CN363_sign_in(28) <= VN1889_sign_out(5);
    CN363_data_in(29) <= VN1945_data_out(5);
    CN363_sign_in(29) <= VN1945_sign_out(5);
    CN363_data_in(30) <= VN1956_data_out(5);
    CN363_sign_in(30) <= VN1956_sign_out(5);
    CN363_data_in(31) <= VN1965_data_out(5);
    CN363_sign_in(31) <= VN1965_sign_out(5);
    CN364_data_in(0) <= VN11_data_out(5);
    CN364_sign_in(0) <= VN11_sign_out(5);
    CN364_data_in(1) <= VN82_data_out(5);
    CN364_sign_in(1) <= VN82_sign_out(5);
    CN364_data_in(2) <= VN129_data_out(5);
    CN364_sign_in(2) <= VN129_sign_out(5);
    CN364_data_in(3) <= VN175_data_out(5);
    CN364_sign_in(3) <= VN175_sign_out(5);
    CN364_data_in(4) <= VN263_data_out(5);
    CN364_sign_in(4) <= VN263_sign_out(5);
    CN364_data_in(5) <= VN313_data_out(5);
    CN364_sign_in(5) <= VN313_sign_out(5);
    CN364_data_in(6) <= VN384_data_out(5);
    CN364_sign_in(6) <= VN384_sign_out(5);
    CN364_data_in(7) <= VN461_data_out(5);
    CN364_sign_in(7) <= VN461_sign_out(5);
    CN364_data_in(8) <= VN526_data_out(5);
    CN364_sign_in(8) <= VN526_sign_out(5);
    CN364_data_in(9) <= VN602_data_out(5);
    CN364_sign_in(9) <= VN602_sign_out(5);
    CN364_data_in(10) <= VN636_data_out(5);
    CN364_sign_in(10) <= VN636_sign_out(5);
    CN364_data_in(11) <= VN766_data_out(5);
    CN364_sign_in(11) <= VN766_sign_out(5);
    CN364_data_in(12) <= VN807_data_out(5);
    CN364_sign_in(12) <= VN807_sign_out(5);
    CN364_data_in(13) <= VN884_data_out(5);
    CN364_sign_in(13) <= VN884_sign_out(5);
    CN364_data_in(14) <= VN935_data_out(5);
    CN364_sign_in(14) <= VN935_sign_out(5);
    CN364_data_in(15) <= VN966_data_out(5);
    CN364_sign_in(15) <= VN966_sign_out(5);
    CN364_data_in(16) <= VN1039_data_out(5);
    CN364_sign_in(16) <= VN1039_sign_out(5);
    CN364_data_in(17) <= VN1078_data_out(5);
    CN364_sign_in(17) <= VN1078_sign_out(5);
    CN364_data_in(18) <= VN1145_data_out(5);
    CN364_sign_in(18) <= VN1145_sign_out(5);
    CN364_data_in(19) <= VN1200_data_out(5);
    CN364_sign_in(19) <= VN1200_sign_out(5);
    CN364_data_in(20) <= VN1270_data_out(5);
    CN364_sign_in(20) <= VN1270_sign_out(5);
    CN364_data_in(21) <= VN1309_data_out(5);
    CN364_sign_in(21) <= VN1309_sign_out(5);
    CN364_data_in(22) <= VN1381_data_out(5);
    CN364_sign_in(22) <= VN1381_sign_out(5);
    CN364_data_in(23) <= VN1450_data_out(5);
    CN364_sign_in(23) <= VN1450_sign_out(5);
    CN364_data_in(24) <= VN1498_data_out(5);
    CN364_sign_in(24) <= VN1498_sign_out(5);
    CN364_data_in(25) <= VN1646_data_out(5);
    CN364_sign_in(25) <= VN1646_sign_out(5);
    CN364_data_in(26) <= VN1661_data_out(5);
    CN364_sign_in(26) <= VN1661_sign_out(5);
    CN364_data_in(27) <= VN1763_data_out(5);
    CN364_sign_in(27) <= VN1763_sign_out(5);
    CN364_data_in(28) <= VN1786_data_out(5);
    CN364_sign_in(28) <= VN1786_sign_out(5);
    CN364_data_in(29) <= VN1967_data_out(5);
    CN364_sign_in(29) <= VN1967_sign_out(5);
    CN364_data_in(30) <= VN2035_data_out(5);
    CN364_sign_in(30) <= VN2035_sign_out(5);
    CN364_data_in(31) <= VN2042_data_out(5);
    CN364_sign_in(31) <= VN2042_sign_out(5);
    CN365_data_in(0) <= VN10_data_out(5);
    CN365_sign_in(0) <= VN10_sign_out(5);
    CN365_data_in(1) <= VN98_data_out(5);
    CN365_sign_in(1) <= VN98_sign_out(5);
    CN365_data_in(2) <= VN142_data_out(5);
    CN365_sign_in(2) <= VN142_sign_out(5);
    CN365_data_in(3) <= VN194_data_out(5);
    CN365_sign_in(3) <= VN194_sign_out(5);
    CN365_data_in(4) <= VN234_data_out(5);
    CN365_sign_in(4) <= VN234_sign_out(5);
    CN365_data_in(5) <= VN298_data_out(5);
    CN365_sign_in(5) <= VN298_sign_out(5);
    CN365_data_in(6) <= VN418_data_out(5);
    CN365_sign_in(6) <= VN418_sign_out(5);
    CN365_data_in(7) <= VN458_data_out(5);
    CN365_sign_in(7) <= VN458_sign_out(5);
    CN365_data_in(8) <= VN590_data_out(5);
    CN365_sign_in(8) <= VN590_sign_out(5);
    CN365_data_in(9) <= VN617_data_out(5);
    CN365_sign_in(9) <= VN617_sign_out(5);
    CN365_data_in(10) <= VN702_data_out(5);
    CN365_sign_in(10) <= VN702_sign_out(5);
    CN365_data_in(11) <= VN734_data_out(5);
    CN365_sign_in(11) <= VN734_sign_out(5);
    CN365_data_in(12) <= VN803_data_out(5);
    CN365_sign_in(12) <= VN803_sign_out(5);
    CN365_data_in(13) <= VN840_data_out(5);
    CN365_sign_in(13) <= VN840_sign_out(5);
    CN365_data_in(14) <= VN919_data_out(5);
    CN365_sign_in(14) <= VN919_sign_out(5);
    CN365_data_in(15) <= VN963_data_out(5);
    CN365_sign_in(15) <= VN963_sign_out(5);
    CN365_data_in(16) <= VN1040_data_out(5);
    CN365_sign_in(16) <= VN1040_sign_out(5);
    CN365_data_in(17) <= VN1086_data_out(5);
    CN365_sign_in(17) <= VN1086_sign_out(5);
    CN365_data_in(18) <= VN1150_data_out(5);
    CN365_sign_in(18) <= VN1150_sign_out(5);
    CN365_data_in(19) <= VN1325_data_out(5);
    CN365_sign_in(19) <= VN1325_sign_out(5);
    CN365_data_in(20) <= VN1347_data_out(5);
    CN365_sign_in(20) <= VN1347_sign_out(5);
    CN365_data_in(21) <= VN1390_data_out(5);
    CN365_sign_in(21) <= VN1390_sign_out(5);
    CN365_data_in(22) <= VN1415_data_out(5);
    CN365_sign_in(22) <= VN1415_sign_out(5);
    CN365_data_in(23) <= VN1497_data_out(5);
    CN365_sign_in(23) <= VN1497_sign_out(5);
    CN365_data_in(24) <= VN1517_data_out(5);
    CN365_sign_in(24) <= VN1517_sign_out(5);
    CN365_data_in(25) <= VN1521_data_out(5);
    CN365_sign_in(25) <= VN1521_sign_out(5);
    CN365_data_in(26) <= VN1556_data_out(5);
    CN365_sign_in(26) <= VN1556_sign_out(5);
    CN365_data_in(27) <= VN1586_data_out(5);
    CN365_sign_in(27) <= VN1586_sign_out(5);
    CN365_data_in(28) <= VN1624_data_out(5);
    CN365_sign_in(28) <= VN1624_sign_out(5);
    CN365_data_in(29) <= VN1679_data_out(5);
    CN365_sign_in(29) <= VN1679_sign_out(5);
    CN365_data_in(30) <= VN1768_data_out(5);
    CN365_sign_in(30) <= VN1768_sign_out(5);
    CN365_data_in(31) <= VN1875_data_out(5);
    CN365_sign_in(31) <= VN1875_sign_out(5);
    CN366_data_in(0) <= VN9_data_out(5);
    CN366_sign_in(0) <= VN9_sign_out(5);
    CN366_data_in(1) <= VN102_data_out(5);
    CN366_sign_in(1) <= VN102_sign_out(5);
    CN366_data_in(2) <= VN153_data_out(5);
    CN366_sign_in(2) <= VN153_sign_out(5);
    CN366_data_in(3) <= VN219_data_out(5);
    CN366_sign_in(3) <= VN219_sign_out(5);
    CN366_data_in(4) <= VN269_data_out(5);
    CN366_sign_in(4) <= VN269_sign_out(5);
    CN366_data_in(5) <= VN308_data_out(5);
    CN366_sign_in(5) <= VN308_sign_out(5);
    CN366_data_in(6) <= VN388_data_out(5);
    CN366_sign_in(6) <= VN388_sign_out(5);
    CN366_data_in(7) <= VN473_data_out(5);
    CN366_sign_in(7) <= VN473_sign_out(5);
    CN366_data_in(8) <= VN525_data_out(5);
    CN366_sign_in(8) <= VN525_sign_out(5);
    CN366_data_in(9) <= VN607_data_out(5);
    CN366_sign_in(9) <= VN607_sign_out(5);
    CN366_data_in(10) <= VN652_data_out(5);
    CN366_sign_in(10) <= VN652_sign_out(5);
    CN366_data_in(11) <= VN696_data_out(5);
    CN366_sign_in(11) <= VN696_sign_out(5);
    CN366_data_in(12) <= VN740_data_out(5);
    CN366_sign_in(12) <= VN740_sign_out(5);
    CN366_data_in(13) <= VN808_data_out(5);
    CN366_sign_in(13) <= VN808_sign_out(5);
    CN366_data_in(14) <= VN849_data_out(5);
    CN366_sign_in(14) <= VN849_sign_out(5);
    CN366_data_in(15) <= VN926_data_out(5);
    CN366_sign_in(15) <= VN926_sign_out(5);
    CN366_data_in(16) <= VN982_data_out(5);
    CN366_sign_in(16) <= VN982_sign_out(5);
    CN366_data_in(17) <= VN1018_data_out(5);
    CN366_sign_in(17) <= VN1018_sign_out(5);
    CN366_data_in(18) <= VN1081_data_out(5);
    CN366_sign_in(18) <= VN1081_sign_out(5);
    CN366_data_in(19) <= VN1242_data_out(5);
    CN366_sign_in(19) <= VN1242_sign_out(5);
    CN366_data_in(20) <= VN1277_data_out(5);
    CN366_sign_in(20) <= VN1277_sign_out(5);
    CN366_data_in(21) <= VN1292_data_out(5);
    CN366_sign_in(21) <= VN1292_sign_out(5);
    CN366_data_in(22) <= VN1348_data_out(5);
    CN366_sign_in(22) <= VN1348_sign_out(5);
    CN366_data_in(23) <= VN1514_data_out(5);
    CN366_sign_in(23) <= VN1514_sign_out(5);
    CN366_data_in(24) <= VN1635_data_out(5);
    CN366_sign_in(24) <= VN1635_sign_out(5);
    CN366_data_in(25) <= VN1668_data_out(5);
    CN366_sign_in(25) <= VN1668_sign_out(5);
    CN366_data_in(26) <= VN1690_data_out(5);
    CN366_sign_in(26) <= VN1690_sign_out(5);
    CN366_data_in(27) <= VN1744_data_out(5);
    CN366_sign_in(27) <= VN1744_sign_out(5);
    CN366_data_in(28) <= VN1748_data_out(5);
    CN366_sign_in(28) <= VN1748_sign_out(5);
    CN366_data_in(29) <= VN1986_data_out(5);
    CN366_sign_in(29) <= VN1986_sign_out(5);
    CN366_data_in(30) <= VN2031_data_out(5);
    CN366_sign_in(30) <= VN2031_sign_out(5);
    CN366_data_in(31) <= VN2039_data_out(5);
    CN366_sign_in(31) <= VN2039_sign_out(5);
    CN367_data_in(0) <= VN8_data_out(5);
    CN367_sign_in(0) <= VN8_sign_out(5);
    CN367_data_in(1) <= VN110_data_out(5);
    CN367_sign_in(1) <= VN110_sign_out(5);
    CN367_data_in(2) <= VN123_data_out(5);
    CN367_sign_in(2) <= VN123_sign_out(5);
    CN367_data_in(3) <= VN205_data_out(5);
    CN367_sign_in(3) <= VN205_sign_out(5);
    CN367_data_in(4) <= VN226_data_out(5);
    CN367_sign_in(4) <= VN226_sign_out(5);
    CN367_data_in(5) <= VN320_data_out(5);
    CN367_sign_in(5) <= VN320_sign_out(5);
    CN367_data_in(6) <= VN333_data_out(5);
    CN367_sign_in(6) <= VN333_sign_out(5);
    CN367_data_in(7) <= VN397_data_out(5);
    CN367_sign_in(7) <= VN397_sign_out(5);
    CN367_data_in(8) <= VN466_data_out(5);
    CN367_sign_in(8) <= VN466_sign_out(5);
    CN367_data_in(9) <= VN520_data_out(5);
    CN367_sign_in(9) <= VN520_sign_out(5);
    CN367_data_in(10) <= VN678_data_out(5);
    CN367_sign_in(10) <= VN678_sign_out(5);
    CN367_data_in(11) <= VN799_data_out(5);
    CN367_sign_in(11) <= VN799_sign_out(5);
    CN367_data_in(12) <= VN891_data_out(5);
    CN367_sign_in(12) <= VN891_sign_out(5);
    CN367_data_in(13) <= VN945_data_out(5);
    CN367_sign_in(13) <= VN945_sign_out(5);
    CN367_data_in(14) <= VN1010_data_out(5);
    CN367_sign_in(14) <= VN1010_sign_out(5);
    CN367_data_in(15) <= VN1087_data_out(5);
    CN367_sign_in(15) <= VN1087_sign_out(5);
    CN367_data_in(16) <= VN1149_data_out(5);
    CN367_sign_in(16) <= VN1149_sign_out(5);
    CN367_data_in(17) <= VN1241_data_out(5);
    CN367_sign_in(17) <= VN1241_sign_out(5);
    CN367_data_in(18) <= VN1300_data_out(5);
    CN367_sign_in(18) <= VN1300_sign_out(5);
    CN367_data_in(19) <= VN1380_data_out(5);
    CN367_sign_in(19) <= VN1380_sign_out(5);
    CN367_data_in(20) <= VN1494_data_out(5);
    CN367_sign_in(20) <= VN1494_sign_out(5);
    CN367_data_in(21) <= VN1589_data_out(5);
    CN367_sign_in(21) <= VN1589_sign_out(5);
    CN367_data_in(22) <= VN1611_data_out(5);
    CN367_sign_in(22) <= VN1611_sign_out(5);
    CN367_data_in(23) <= VN1694_data_out(5);
    CN367_sign_in(23) <= VN1694_sign_out(5);
    CN367_data_in(24) <= VN1734_data_out(5);
    CN367_sign_in(24) <= VN1734_sign_out(5);
    CN367_data_in(25) <= VN1735_data_out(5);
    CN367_sign_in(25) <= VN1735_sign_out(5);
    CN367_data_in(26) <= VN1749_data_out(5);
    CN367_sign_in(26) <= VN1749_sign_out(5);
    CN367_data_in(27) <= VN1800_data_out(5);
    CN367_sign_in(27) <= VN1800_sign_out(5);
    CN367_data_in(28) <= VN1857_data_out(5);
    CN367_sign_in(28) <= VN1857_sign_out(5);
    CN367_data_in(29) <= VN1919_data_out(5);
    CN367_sign_in(29) <= VN1919_sign_out(5);
    CN367_data_in(30) <= VN1934_data_out(5);
    CN367_sign_in(30) <= VN1934_sign_out(5);
    CN367_data_in(31) <= VN1950_data_out(5);
    CN367_sign_in(31) <= VN1950_sign_out(5);
    CN368_data_in(0) <= VN7_data_out(5);
    CN368_sign_in(0) <= VN7_sign_out(5);
    CN368_data_in(1) <= VN177_data_out(5);
    CN368_sign_in(1) <= VN177_sign_out(5);
    CN368_data_in(2) <= VN381_data_out(5);
    CN368_sign_in(2) <= VN381_sign_out(5);
    CN368_data_in(3) <= VN414_data_out(5);
    CN368_sign_in(3) <= VN414_sign_out(5);
    CN368_data_in(4) <= VN496_data_out(5);
    CN368_sign_in(4) <= VN496_sign_out(5);
    CN368_data_in(5) <= VN560_data_out(5);
    CN368_sign_in(5) <= VN560_sign_out(5);
    CN368_data_in(6) <= VN580_data_out(5);
    CN368_sign_in(6) <= VN580_sign_out(5);
    CN368_data_in(7) <= VN639_data_out(5);
    CN368_sign_in(7) <= VN639_sign_out(5);
    CN368_data_in(8) <= VN685_data_out(5);
    CN368_sign_in(8) <= VN685_sign_out(5);
    CN368_data_in(9) <= VN726_data_out(5);
    CN368_sign_in(9) <= VN726_sign_out(5);
    CN368_data_in(10) <= VN822_data_out(5);
    CN368_sign_in(10) <= VN822_sign_out(5);
    CN368_data_in(11) <= VN889_data_out(5);
    CN368_sign_in(11) <= VN889_sign_out(5);
    CN368_data_in(12) <= VN946_data_out(5);
    CN368_sign_in(12) <= VN946_sign_out(5);
    CN368_data_in(13) <= VN1026_data_out(5);
    CN368_sign_in(13) <= VN1026_sign_out(5);
    CN368_data_in(14) <= VN1143_data_out(5);
    CN368_sign_in(14) <= VN1143_sign_out(5);
    CN368_data_in(15) <= VN1180_data_out(5);
    CN368_sign_in(15) <= VN1180_sign_out(5);
    CN368_data_in(16) <= VN1296_data_out(5);
    CN368_sign_in(16) <= VN1296_sign_out(5);
    CN368_data_in(17) <= VN1372_data_out(5);
    CN368_sign_in(17) <= VN1372_sign_out(5);
    CN368_data_in(18) <= VN1467_data_out(5);
    CN368_sign_in(18) <= VN1467_sign_out(5);
    CN368_data_in(19) <= VN1545_data_out(5);
    CN368_sign_in(19) <= VN1545_sign_out(5);
    CN368_data_in(20) <= VN1641_data_out(5);
    CN368_sign_in(20) <= VN1641_sign_out(5);
    CN368_data_in(21) <= VN1714_data_out(5);
    CN368_sign_in(21) <= VN1714_sign_out(5);
    CN368_data_in(22) <= VN1787_data_out(5);
    CN368_sign_in(22) <= VN1787_sign_out(5);
    CN368_data_in(23) <= VN1837_data_out(5);
    CN368_sign_in(23) <= VN1837_sign_out(5);
    CN368_data_in(24) <= VN1859_data_out(5);
    CN368_sign_in(24) <= VN1859_sign_out(5);
    CN368_data_in(25) <= VN1907_data_out(5);
    CN368_sign_in(25) <= VN1907_sign_out(5);
    CN368_data_in(26) <= VN1916_data_out(5);
    CN368_sign_in(26) <= VN1916_sign_out(5);
    CN368_data_in(27) <= VN1940_data_out(5);
    CN368_sign_in(27) <= VN1940_sign_out(5);
    CN368_data_in(28) <= VN1952_data_out(5);
    CN368_sign_in(28) <= VN1952_sign_out(5);
    CN368_data_in(29) <= VN1989_data_out(5);
    CN368_sign_in(29) <= VN1989_sign_out(5);
    CN368_data_in(30) <= VN2040_data_out(5);
    CN368_sign_in(30) <= VN2040_sign_out(5);
    CN368_data_in(31) <= VN2046_data_out(5);
    CN368_sign_in(31) <= VN2046_sign_out(5);
    CN369_data_in(0) <= VN6_data_out(5);
    CN369_sign_in(0) <= VN6_sign_out(5);
    CN369_data_in(1) <= VN156_data_out(5);
    CN369_sign_in(1) <= VN156_sign_out(5);
    CN369_data_in(2) <= VN221_data_out(5);
    CN369_sign_in(2) <= VN221_sign_out(5);
    CN369_data_in(3) <= VN262_data_out(5);
    CN369_sign_in(3) <= VN262_sign_out(5);
    CN369_data_in(4) <= VN358_data_out(5);
    CN369_sign_in(4) <= VN358_sign_out(5);
    CN369_data_in(5) <= VN445_data_out(5);
    CN369_sign_in(5) <= VN445_sign_out(5);
    CN369_data_in(6) <= VN450_data_out(5);
    CN369_sign_in(6) <= VN450_sign_out(5);
    CN369_data_in(7) <= VN511_data_out(5);
    CN369_sign_in(7) <= VN511_sign_out(5);
    CN369_data_in(8) <= VN594_data_out(5);
    CN369_sign_in(8) <= VN594_sign_out(5);
    CN369_data_in(9) <= VN618_data_out(5);
    CN369_sign_in(9) <= VN618_sign_out(5);
    CN369_data_in(10) <= VN708_data_out(5);
    CN369_sign_in(10) <= VN708_sign_out(5);
    CN369_data_in(11) <= VN750_data_out(5);
    CN369_sign_in(11) <= VN750_sign_out(5);
    CN369_data_in(12) <= VN827_data_out(5);
    CN369_sign_in(12) <= VN827_sign_out(5);
    CN369_data_in(13) <= VN924_data_out(5);
    CN369_sign_in(13) <= VN924_sign_out(5);
    CN369_data_in(14) <= VN981_data_out(5);
    CN369_sign_in(14) <= VN981_sign_out(5);
    CN369_data_in(15) <= VN1030_data_out(5);
    CN369_sign_in(15) <= VN1030_sign_out(5);
    CN369_data_in(16) <= VN1125_data_out(5);
    CN369_sign_in(16) <= VN1125_sign_out(5);
    CN369_data_in(17) <= VN1166_data_out(5);
    CN369_sign_in(17) <= VN1166_sign_out(5);
    CN369_data_in(18) <= VN1183_data_out(5);
    CN369_sign_in(18) <= VN1183_sign_out(5);
    CN369_data_in(19) <= VN1255_data_out(5);
    CN369_sign_in(19) <= VN1255_sign_out(5);
    CN369_data_in(20) <= VN1335_data_out(5);
    CN369_sign_in(20) <= VN1335_sign_out(5);
    CN369_data_in(21) <= VN1422_data_out(5);
    CN369_sign_in(21) <= VN1422_sign_out(5);
    CN369_data_in(22) <= VN1570_data_out(5);
    CN369_sign_in(22) <= VN1570_sign_out(5);
    CN369_data_in(23) <= VN1585_data_out(5);
    CN369_sign_in(23) <= VN1585_sign_out(5);
    CN369_data_in(24) <= VN1612_data_out(5);
    CN369_sign_in(24) <= VN1612_sign_out(5);
    CN369_data_in(25) <= VN1670_data_out(5);
    CN369_sign_in(25) <= VN1670_sign_out(5);
    CN369_data_in(26) <= VN1715_data_out(5);
    CN369_sign_in(26) <= VN1715_sign_out(5);
    CN369_data_in(27) <= VN1917_data_out(5);
    CN369_sign_in(27) <= VN1917_sign_out(5);
    CN369_data_in(28) <= VN1998_data_out(5);
    CN369_sign_in(28) <= VN1998_sign_out(5);
    CN369_data_in(29) <= VN2008_data_out(5);
    CN369_sign_in(29) <= VN2008_sign_out(5);
    CN369_data_in(30) <= VN2017_data_out(5);
    CN369_sign_in(30) <= VN2017_sign_out(5);
    CN369_data_in(31) <= VN2030_data_out(5);
    CN369_sign_in(31) <= VN2030_sign_out(5);
    CN370_data_in(0) <= VN5_data_out(5);
    CN370_sign_in(0) <= VN5_sign_out(5);
    CN370_data_in(1) <= VN114_data_out(5);
    CN370_sign_in(1) <= VN114_sign_out(5);
    CN370_data_in(2) <= VN208_data_out(5);
    CN370_sign_in(2) <= VN208_sign_out(5);
    CN370_data_in(3) <= VN275_data_out(5);
    CN370_sign_in(3) <= VN275_sign_out(5);
    CN370_data_in(4) <= VN341_data_out(5);
    CN370_sign_in(4) <= VN341_sign_out(5);
    CN370_data_in(5) <= VN442_data_out(5);
    CN370_sign_in(5) <= VN442_sign_out(5);
    CN370_data_in(6) <= VN500_data_out(5);
    CN370_sign_in(6) <= VN500_sign_out(5);
    CN370_data_in(7) <= VN532_data_out(5);
    CN370_sign_in(7) <= VN532_sign_out(5);
    CN370_data_in(8) <= VN635_data_out(5);
    CN370_sign_in(8) <= VN635_sign_out(5);
    CN370_data_in(9) <= VN706_data_out(5);
    CN370_sign_in(9) <= VN706_sign_out(5);
    CN370_data_in(10) <= VN732_data_out(5);
    CN370_sign_in(10) <= VN732_sign_out(5);
    CN370_data_in(11) <= VN812_data_out(5);
    CN370_sign_in(11) <= VN812_sign_out(5);
    CN370_data_in(12) <= VN843_data_out(5);
    CN370_sign_in(12) <= VN843_sign_out(5);
    CN370_data_in(13) <= VN905_data_out(5);
    CN370_sign_in(13) <= VN905_sign_out(5);
    CN370_data_in(14) <= VN973_data_out(5);
    CN370_sign_in(14) <= VN973_sign_out(5);
    CN370_data_in(15) <= VN1103_data_out(5);
    CN370_sign_in(15) <= VN1103_sign_out(5);
    CN370_data_in(16) <= VN1110_data_out(5);
    CN370_sign_in(16) <= VN1110_sign_out(5);
    CN370_data_in(17) <= VN1132_data_out(5);
    CN370_sign_in(17) <= VN1132_sign_out(5);
    CN370_data_in(18) <= VN1257_data_out(5);
    CN370_sign_in(18) <= VN1257_sign_out(5);
    CN370_data_in(19) <= VN1291_data_out(5);
    CN370_sign_in(19) <= VN1291_sign_out(5);
    CN370_data_in(20) <= VN1393_data_out(5);
    CN370_sign_in(20) <= VN1393_sign_out(5);
    CN370_data_in(21) <= VN1435_data_out(5);
    CN370_sign_in(21) <= VN1435_sign_out(5);
    CN370_data_in(22) <= VN1505_data_out(5);
    CN370_sign_in(22) <= VN1505_sign_out(5);
    CN370_data_in(23) <= VN1518_data_out(5);
    CN370_sign_in(23) <= VN1518_sign_out(5);
    CN370_data_in(24) <= VN1603_data_out(5);
    CN370_sign_in(24) <= VN1603_sign_out(5);
    CN370_data_in(25) <= VN1745_data_out(5);
    CN370_sign_in(25) <= VN1745_sign_out(5);
    CN370_data_in(26) <= VN1757_data_out(5);
    CN370_sign_in(26) <= VN1757_sign_out(5);
    CN370_data_in(27) <= VN1778_data_out(5);
    CN370_sign_in(27) <= VN1778_sign_out(5);
    CN370_data_in(28) <= VN1826_data_out(5);
    CN370_sign_in(28) <= VN1826_sign_out(5);
    CN370_data_in(29) <= VN1910_data_out(5);
    CN370_sign_in(29) <= VN1910_sign_out(5);
    CN370_data_in(30) <= VN2033_data_out(5);
    CN370_sign_in(30) <= VN2033_sign_out(5);
    CN370_data_in(31) <= VN2036_data_out(5);
    CN370_sign_in(31) <= VN2036_sign_out(5);
    CN371_data_in(0) <= VN4_data_out(5);
    CN371_sign_in(0) <= VN4_sign_out(5);
    CN371_data_in(1) <= VN135_data_out(5);
    CN371_sign_in(1) <= VN135_sign_out(5);
    CN371_data_in(2) <= VN173_data_out(5);
    CN371_sign_in(2) <= VN173_sign_out(5);
    CN371_data_in(3) <= VN249_data_out(5);
    CN371_sign_in(3) <= VN249_sign_out(5);
    CN371_data_in(4) <= VN354_data_out(5);
    CN371_sign_in(4) <= VN354_sign_out(5);
    CN371_data_in(5) <= VN401_data_out(5);
    CN371_sign_in(5) <= VN401_sign_out(5);
    CN371_data_in(6) <= VN504_data_out(5);
    CN371_sign_in(6) <= VN504_sign_out(5);
    CN371_data_in(7) <= VN530_data_out(5);
    CN371_sign_in(7) <= VN530_sign_out(5);
    CN371_data_in(8) <= VN563_data_out(5);
    CN371_sign_in(8) <= VN563_sign_out(5);
    CN371_data_in(9) <= VN662_data_out(5);
    CN371_sign_in(9) <= VN662_sign_out(5);
    CN371_data_in(10) <= VN683_data_out(5);
    CN371_sign_in(10) <= VN683_sign_out(5);
    CN371_data_in(11) <= VN744_data_out(5);
    CN371_sign_in(11) <= VN744_sign_out(5);
    CN371_data_in(12) <= VN814_data_out(5);
    CN371_sign_in(12) <= VN814_sign_out(5);
    CN371_data_in(13) <= VN866_data_out(5);
    CN371_sign_in(13) <= VN866_sign_out(5);
    CN371_data_in(14) <= VN908_data_out(5);
    CN371_sign_in(14) <= VN908_sign_out(5);
    CN371_data_in(15) <= VN991_data_out(5);
    CN371_sign_in(15) <= VN991_sign_out(5);
    CN371_data_in(16) <= VN1029_data_out(5);
    CN371_sign_in(16) <= VN1029_sign_out(5);
    CN371_data_in(17) <= VN1155_data_out(5);
    CN371_sign_in(17) <= VN1155_sign_out(5);
    CN371_data_in(18) <= VN1167_data_out(5);
    CN371_sign_in(18) <= VN1167_sign_out(5);
    CN371_data_in(19) <= VN1199_data_out(5);
    CN371_sign_in(19) <= VN1199_sign_out(5);
    CN371_data_in(20) <= VN1243_data_out(5);
    CN371_sign_in(20) <= VN1243_sign_out(5);
    CN371_data_in(21) <= VN1311_data_out(5);
    CN371_sign_in(21) <= VN1311_sign_out(5);
    CN371_data_in(22) <= VN1386_data_out(5);
    CN371_sign_in(22) <= VN1386_sign_out(5);
    CN371_data_in(23) <= VN1461_data_out(5);
    CN371_sign_in(23) <= VN1461_sign_out(5);
    CN371_data_in(24) <= VN1536_data_out(5);
    CN371_sign_in(24) <= VN1536_sign_out(5);
    CN371_data_in(25) <= VN1547_data_out(5);
    CN371_sign_in(25) <= VN1547_sign_out(5);
    CN371_data_in(26) <= VN1622_data_out(5);
    CN371_sign_in(26) <= VN1622_sign_out(5);
    CN371_data_in(27) <= VN1689_data_out(5);
    CN371_sign_in(27) <= VN1689_sign_out(5);
    CN371_data_in(28) <= VN1766_data_out(5);
    CN371_sign_in(28) <= VN1766_sign_out(5);
    CN371_data_in(29) <= VN1988_data_out(5);
    CN371_sign_in(29) <= VN1988_sign_out(5);
    CN371_data_in(30) <= VN2038_data_out(5);
    CN371_sign_in(30) <= VN2038_sign_out(5);
    CN371_data_in(31) <= VN2045_data_out(5);
    CN371_sign_in(31) <= VN2045_sign_out(5);
    CN372_data_in(0) <= VN106_data_out(5);
    CN372_sign_in(0) <= VN106_sign_out(5);
    CN372_data_in(1) <= VN144_data_out(5);
    CN372_sign_in(1) <= VN144_sign_out(5);
    CN372_data_in(2) <= VN201_data_out(5);
    CN372_sign_in(2) <= VN201_sign_out(5);
    CN372_data_in(3) <= VN229_data_out(5);
    CN372_sign_in(3) <= VN229_sign_out(5);
    CN372_data_in(4) <= VN301_data_out(5);
    CN372_sign_in(4) <= VN301_sign_out(5);
    CN372_data_in(5) <= VN365_data_out(5);
    CN372_sign_in(5) <= VN365_sign_out(5);
    CN372_data_in(6) <= VN394_data_out(5);
    CN372_sign_in(6) <= VN394_sign_out(5);
    CN372_data_in(7) <= VN493_data_out(5);
    CN372_sign_in(7) <= VN493_sign_out(5);
    CN372_data_in(8) <= VN573_data_out(5);
    CN372_sign_in(8) <= VN573_sign_out(5);
    CN372_data_in(9) <= VN648_data_out(5);
    CN372_sign_in(9) <= VN648_sign_out(5);
    CN372_data_in(10) <= VN751_data_out(5);
    CN372_sign_in(10) <= VN751_sign_out(5);
    CN372_data_in(11) <= VN878_data_out(5);
    CN372_sign_in(11) <= VN878_sign_out(5);
    CN372_data_in(12) <= VN887_data_out(5);
    CN372_sign_in(12) <= VN887_sign_out(5);
    CN372_data_in(13) <= VN892_data_out(5);
    CN372_sign_in(13) <= VN892_sign_out(5);
    CN372_data_in(14) <= VN995_data_out(5);
    CN372_sign_in(14) <= VN995_sign_out(5);
    CN372_data_in(15) <= VN1090_data_out(5);
    CN372_sign_in(15) <= VN1090_sign_out(5);
    CN372_data_in(16) <= VN1317_data_out(5);
    CN372_sign_in(16) <= VN1317_sign_out(5);
    CN372_data_in(17) <= VN1337_data_out(5);
    CN372_sign_in(17) <= VN1337_sign_out(5);
    CN372_data_in(18) <= VN1469_data_out(5);
    CN372_sign_in(18) <= VN1469_sign_out(5);
    CN372_data_in(19) <= VN1516_data_out(5);
    CN372_sign_in(19) <= VN1516_sign_out(5);
    CN372_data_in(20) <= VN1520_data_out(5);
    CN372_sign_in(20) <= VN1520_sign_out(5);
    CN372_data_in(21) <= VN1595_data_out(5);
    CN372_sign_in(21) <= VN1595_sign_out(5);
    CN372_data_in(22) <= VN1664_data_out(5);
    CN372_sign_in(22) <= VN1664_sign_out(5);
    CN372_data_in(23) <= VN1772_data_out(5);
    CN372_sign_in(23) <= VN1772_sign_out(5);
    CN372_data_in(24) <= VN1793_data_out(5);
    CN372_sign_in(24) <= VN1793_sign_out(5);
    CN372_data_in(25) <= VN1937_data_out(5);
    CN372_sign_in(25) <= VN1937_sign_out(5);
    CN372_data_in(26) <= VN1985_data_out(5);
    CN372_sign_in(26) <= VN1985_sign_out(5);
    CN372_data_in(27) <= VN2010_data_out(5);
    CN372_sign_in(27) <= VN2010_sign_out(5);
    CN372_data_in(28) <= VN2023_data_out(5);
    CN372_sign_in(28) <= VN2023_sign_out(5);
    CN372_data_in(29) <= VN2024_data_out(5);
    CN372_sign_in(29) <= VN2024_sign_out(5);
    CN372_data_in(30) <= VN2037_data_out(5);
    CN372_sign_in(30) <= VN2037_sign_out(5);
    CN372_data_in(31) <= VN2044_data_out(5);
    CN372_sign_in(31) <= VN2044_sign_out(5);
    CN373_data_in(0) <= VN3_data_out(5);
    CN373_sign_in(0) <= VN3_sign_out(5);
    CN373_data_in(1) <= VN139_data_out(5);
    CN373_sign_in(1) <= VN139_sign_out(5);
    CN373_data_in(2) <= VN250_data_out(5);
    CN373_sign_in(2) <= VN250_sign_out(5);
    CN373_data_in(3) <= VN310_data_out(5);
    CN373_sign_in(3) <= VN310_sign_out(5);
    CN373_data_in(4) <= VN335_data_out(5);
    CN373_sign_in(4) <= VN335_sign_out(5);
    CN373_data_in(5) <= VN425_data_out(5);
    CN373_sign_in(5) <= VN425_sign_out(5);
    CN373_data_in(6) <= VN474_data_out(5);
    CN373_sign_in(6) <= VN474_sign_out(5);
    CN373_data_in(7) <= VN546_data_out(5);
    CN373_sign_in(7) <= VN546_sign_out(5);
    CN373_data_in(8) <= VN567_data_out(5);
    CN373_sign_in(8) <= VN567_sign_out(5);
    CN373_data_in(9) <= VN620_data_out(5);
    CN373_sign_in(9) <= VN620_sign_out(5);
    CN373_data_in(10) <= VN721_data_out(5);
    CN373_sign_in(10) <= VN721_sign_out(5);
    CN373_data_in(11) <= VN725_data_out(5);
    CN373_sign_in(11) <= VN725_sign_out(5);
    CN373_data_in(12) <= VN820_data_out(5);
    CN373_sign_in(12) <= VN820_sign_out(5);
    CN373_data_in(13) <= VN875_data_out(5);
    CN373_sign_in(13) <= VN875_sign_out(5);
    CN373_data_in(14) <= VN925_data_out(5);
    CN373_sign_in(14) <= VN925_sign_out(5);
    CN373_data_in(15) <= VN1062_data_out(5);
    CN373_sign_in(15) <= VN1062_sign_out(5);
    CN373_data_in(16) <= VN1130_data_out(5);
    CN373_sign_in(16) <= VN1130_sign_out(5);
    CN373_data_in(17) <= VN1192_data_out(5);
    CN373_sign_in(17) <= VN1192_sign_out(5);
    CN373_data_in(18) <= VN1279_data_out(5);
    CN373_sign_in(18) <= VN1279_sign_out(5);
    CN373_data_in(19) <= VN1303_data_out(5);
    CN373_sign_in(19) <= VN1303_sign_out(5);
    CN373_data_in(20) <= VN1391_data_out(5);
    CN373_sign_in(20) <= VN1391_sign_out(5);
    CN373_data_in(21) <= VN1437_data_out(5);
    CN373_sign_in(21) <= VN1437_sign_out(5);
    CN373_data_in(22) <= VN1503_data_out(5);
    CN373_sign_in(22) <= VN1503_sign_out(5);
    CN373_data_in(23) <= VN1596_data_out(5);
    CN373_sign_in(23) <= VN1596_sign_out(5);
    CN373_data_in(24) <= VN1608_data_out(5);
    CN373_sign_in(24) <= VN1608_sign_out(5);
    CN373_data_in(25) <= VN1673_data_out(5);
    CN373_sign_in(25) <= VN1673_sign_out(5);
    CN373_data_in(26) <= VN1702_data_out(5);
    CN373_sign_in(26) <= VN1702_sign_out(5);
    CN373_data_in(27) <= VN1884_data_out(5);
    CN373_sign_in(27) <= VN1884_sign_out(5);
    CN373_data_in(28) <= VN1906_data_out(5);
    CN373_sign_in(28) <= VN1906_sign_out(5);
    CN373_data_in(29) <= VN1938_data_out(5);
    CN373_sign_in(29) <= VN1938_sign_out(5);
    CN373_data_in(30) <= VN1949_data_out(5);
    CN373_sign_in(30) <= VN1949_sign_out(5);
    CN373_data_in(31) <= VN1960_data_out(5);
    CN373_sign_in(31) <= VN1960_sign_out(5);
    CN374_data_in(0) <= VN2_data_out(5);
    CN374_sign_in(0) <= VN2_sign_out(5);
    CN374_data_in(1) <= VN85_data_out(5);
    CN374_sign_in(1) <= VN85_sign_out(5);
    CN374_data_in(2) <= VN145_data_out(5);
    CN374_sign_in(2) <= VN145_sign_out(5);
    CN374_data_in(3) <= VN213_data_out(5);
    CN374_sign_in(3) <= VN213_sign_out(5);
    CN374_data_in(4) <= VN264_data_out(5);
    CN374_sign_in(4) <= VN264_sign_out(5);
    CN374_data_in(5) <= VN306_data_out(5);
    CN374_sign_in(5) <= VN306_sign_out(5);
    CN374_data_in(6) <= VN383_data_out(5);
    CN374_sign_in(6) <= VN383_sign_out(5);
    CN374_data_in(7) <= VN436_data_out(5);
    CN374_sign_in(7) <= VN436_sign_out(5);
    CN374_data_in(8) <= VN457_data_out(5);
    CN374_sign_in(8) <= VN457_sign_out(5);
    CN374_data_in(9) <= VN549_data_out(5);
    CN374_sign_in(9) <= VN549_sign_out(5);
    CN374_data_in(10) <= VN570_data_out(5);
    CN374_sign_in(10) <= VN570_sign_out(5);
    CN374_data_in(11) <= VN709_data_out(5);
    CN374_sign_in(11) <= VN709_sign_out(5);
    CN374_data_in(12) <= VN739_data_out(5);
    CN374_sign_in(12) <= VN739_sign_out(5);
    CN374_data_in(13) <= VN778_data_out(5);
    CN374_sign_in(13) <= VN778_sign_out(5);
    CN374_data_in(14) <= VN838_data_out(5);
    CN374_sign_in(14) <= VN838_sign_out(5);
    CN374_data_in(15) <= VN888_data_out(5);
    CN374_sign_in(15) <= VN888_sign_out(5);
    CN374_data_in(16) <= VN994_data_out(5);
    CN374_sign_in(16) <= VN994_sign_out(5);
    CN374_data_in(17) <= VN1014_data_out(5);
    CN374_sign_in(17) <= VN1014_sign_out(5);
    CN374_data_in(18) <= VN1096_data_out(5);
    CN374_sign_in(18) <= VN1096_sign_out(5);
    CN374_data_in(19) <= VN1267_data_out(5);
    CN374_sign_in(19) <= VN1267_sign_out(5);
    CN374_data_in(20) <= VN1332_data_out(5);
    CN374_sign_in(20) <= VN1332_sign_out(5);
    CN374_data_in(21) <= VN1419_data_out(5);
    CN374_sign_in(21) <= VN1419_sign_out(5);
    CN374_data_in(22) <= VN1426_data_out(5);
    CN374_sign_in(22) <= VN1426_sign_out(5);
    CN374_data_in(23) <= VN1480_data_out(5);
    CN374_sign_in(23) <= VN1480_sign_out(5);
    CN374_data_in(24) <= VN1669_data_out(5);
    CN374_sign_in(24) <= VN1669_sign_out(5);
    CN374_data_in(25) <= VN1762_data_out(5);
    CN374_sign_in(25) <= VN1762_sign_out(5);
    CN374_data_in(26) <= VN1790_data_out(5);
    CN374_sign_in(26) <= VN1790_sign_out(5);
    CN374_data_in(27) <= VN1844_data_out(5);
    CN374_sign_in(27) <= VN1844_sign_out(5);
    CN374_data_in(28) <= VN1891_data_out(5);
    CN374_sign_in(28) <= VN1891_sign_out(5);
    CN374_data_in(29) <= VN1930_data_out(5);
    CN374_sign_in(29) <= VN1930_sign_out(5);
    CN374_data_in(30) <= VN1955_data_out(5);
    CN374_sign_in(30) <= VN1955_sign_out(5);
    CN374_data_in(31) <= VN1968_data_out(5);
    CN374_sign_in(31) <= VN1968_sign_out(5);
    CN375_data_in(0) <= VN1_data_out(5);
    CN375_sign_in(0) <= VN1_sign_out(5);
    CN375_data_in(1) <= VN64_data_out(5);
    CN375_sign_in(1) <= VN64_sign_out(5);
    CN375_data_in(2) <= VN134_data_out(5);
    CN375_sign_in(2) <= VN134_sign_out(5);
    CN375_data_in(3) <= VN260_data_out(5);
    CN375_sign_in(3) <= VN260_sign_out(5);
    CN375_data_in(4) <= VN311_data_out(5);
    CN375_sign_in(4) <= VN311_sign_out(5);
    CN375_data_in(5) <= VN368_data_out(5);
    CN375_sign_in(5) <= VN368_sign_out(5);
    CN375_data_in(6) <= VN429_data_out(5);
    CN375_sign_in(6) <= VN429_sign_out(5);
    CN375_data_in(7) <= VN469_data_out(5);
    CN375_sign_in(7) <= VN469_sign_out(5);
    CN375_data_in(8) <= VN533_data_out(5);
    CN375_sign_in(8) <= VN533_sign_out(5);
    CN375_data_in(9) <= VN615_data_out(5);
    CN375_sign_in(9) <= VN615_sign_out(5);
    CN375_data_in(10) <= VN684_data_out(5);
    CN375_sign_in(10) <= VN684_sign_out(5);
    CN375_data_in(11) <= VN768_data_out(5);
    CN375_sign_in(11) <= VN768_sign_out(5);
    CN375_data_in(12) <= VN785_data_out(5);
    CN375_sign_in(12) <= VN785_sign_out(5);
    CN375_data_in(13) <= VN860_data_out(5);
    CN375_sign_in(13) <= VN860_sign_out(5);
    CN375_data_in(14) <= VN916_data_out(5);
    CN375_sign_in(14) <= VN916_sign_out(5);
    CN375_data_in(15) <= VN989_data_out(5);
    CN375_sign_in(15) <= VN989_sign_out(5);
    CN375_data_in(16) <= VN1035_data_out(5);
    CN375_sign_in(16) <= VN1035_sign_out(5);
    CN375_data_in(17) <= VN1107_data_out(5);
    CN375_sign_in(17) <= VN1107_sign_out(5);
    CN375_data_in(18) <= VN1114_data_out(5);
    CN375_sign_in(18) <= VN1114_sign_out(5);
    CN375_data_in(19) <= VN1201_data_out(5);
    CN375_sign_in(19) <= VN1201_sign_out(5);
    CN375_data_in(20) <= VN1218_data_out(5);
    CN375_sign_in(20) <= VN1218_sign_out(5);
    CN375_data_in(21) <= VN1252_data_out(5);
    CN375_sign_in(21) <= VN1252_sign_out(5);
    CN375_data_in(22) <= VN1377_data_out(5);
    CN375_sign_in(22) <= VN1377_sign_out(5);
    CN375_data_in(23) <= VN1416_data_out(5);
    CN375_sign_in(23) <= VN1416_sign_out(5);
    CN375_data_in(24) <= VN1442_data_out(5);
    CN375_sign_in(24) <= VN1442_sign_out(5);
    CN375_data_in(25) <= VN1526_data_out(5);
    CN375_sign_in(25) <= VN1526_sign_out(5);
    CN375_data_in(26) <= VN1602_data_out(5);
    CN375_sign_in(26) <= VN1602_sign_out(5);
    CN375_data_in(27) <= VN1636_data_out(5);
    CN375_sign_in(27) <= VN1636_sign_out(5);
    CN375_data_in(28) <= VN1652_data_out(5);
    CN375_sign_in(28) <= VN1652_sign_out(5);
    CN375_data_in(29) <= VN1848_data_out(5);
    CN375_sign_in(29) <= VN1848_sign_out(5);
    CN375_data_in(30) <= VN1854_data_out(5);
    CN375_sign_in(30) <= VN1854_sign_out(5);
    CN375_data_in(31) <= VN1903_data_out(5);
    CN375_sign_in(31) <= VN1903_sign_out(5);
    CN376_data_in(0) <= VN0_data_out(5);
    CN376_sign_in(0) <= VN0_sign_out(5);
    CN376_data_in(1) <= VN67_data_out(5);
    CN376_sign_in(1) <= VN67_sign_out(5);
    CN376_data_in(2) <= VN159_data_out(5);
    CN376_sign_in(2) <= VN159_sign_out(5);
    CN376_data_in(3) <= VN278_data_out(5);
    CN376_sign_in(3) <= VN278_sign_out(5);
    CN376_data_in(4) <= VN386_data_out(5);
    CN376_sign_in(4) <= VN386_sign_out(5);
    CN376_data_in(5) <= VN433_data_out(5);
    CN376_sign_in(5) <= VN433_sign_out(5);
    CN376_data_in(6) <= VN479_data_out(5);
    CN376_sign_in(6) <= VN479_sign_out(5);
    CN376_data_in(7) <= VN510_data_out(5);
    CN376_sign_in(7) <= VN510_sign_out(5);
    CN376_data_in(8) <= VN595_data_out(5);
    CN376_sign_in(8) <= VN595_sign_out(5);
    CN376_data_in(9) <= VN705_data_out(5);
    CN376_sign_in(9) <= VN705_sign_out(5);
    CN376_data_in(10) <= VN746_data_out(5);
    CN376_sign_in(10) <= VN746_sign_out(5);
    CN376_data_in(11) <= VN813_data_out(5);
    CN376_sign_in(11) <= VN813_sign_out(5);
    CN376_data_in(12) <= VN861_data_out(5);
    CN376_sign_in(12) <= VN861_sign_out(5);
    CN376_data_in(13) <= VN901_data_out(5);
    CN376_sign_in(13) <= VN901_sign_out(5);
    CN376_data_in(14) <= VN970_data_out(5);
    CN376_sign_in(14) <= VN970_sign_out(5);
    CN376_data_in(15) <= VN1063_data_out(5);
    CN376_sign_in(15) <= VN1063_sign_out(5);
    CN376_data_in(16) <= VN1156_data_out(5);
    CN376_sign_in(16) <= VN1156_sign_out(5);
    CN376_data_in(17) <= VN1220_data_out(5);
    CN376_sign_in(17) <= VN1220_sign_out(5);
    CN376_data_in(18) <= VN1334_data_out(5);
    CN376_sign_in(18) <= VN1334_sign_out(5);
    CN376_data_in(19) <= VN1343_data_out(5);
    CN376_sign_in(19) <= VN1343_sign_out(5);
    CN376_data_in(20) <= VN1465_data_out(5);
    CN376_sign_in(20) <= VN1465_sign_out(5);
    CN376_data_in(21) <= VN1522_data_out(5);
    CN376_sign_in(21) <= VN1522_sign_out(5);
    CN376_data_in(22) <= VN1539_data_out(5);
    CN376_sign_in(22) <= VN1539_sign_out(5);
    CN376_data_in(23) <= VN1629_data_out(5);
    CN376_sign_in(23) <= VN1629_sign_out(5);
    CN376_data_in(24) <= VN1659_data_out(5);
    CN376_sign_in(24) <= VN1659_sign_out(5);
    CN376_data_in(25) <= VN1838_data_out(5);
    CN376_sign_in(25) <= VN1838_sign_out(5);
    CN376_data_in(26) <= VN1886_data_out(5);
    CN376_sign_in(26) <= VN1886_sign_out(5);
    CN376_data_in(27) <= VN1912_data_out(5);
    CN376_sign_in(27) <= VN1912_sign_out(5);
    CN376_data_in(28) <= VN1939_data_out(5);
    CN376_sign_in(28) <= VN1939_sign_out(5);
    CN376_data_in(29) <= VN1948_data_out(5);
    CN376_sign_in(29) <= VN1948_sign_out(5);
    CN376_data_in(30) <= VN1954_data_out(5);
    CN376_sign_in(30) <= VN1954_sign_out(5);
    CN376_data_in(31) <= VN1971_data_out(5);
    CN376_sign_in(31) <= VN1971_sign_out(5);
    CN377_data_in(0) <= VN107_data_out(5);
    CN377_sign_in(0) <= VN107_sign_out(5);
    CN377_data_in(1) <= VN166_data_out(5);
    CN377_sign_in(1) <= VN166_sign_out(5);
    CN377_data_in(2) <= VN193_data_out(5);
    CN377_sign_in(2) <= VN193_sign_out(5);
    CN377_data_in(3) <= VN325_data_out(5);
    CN377_sign_in(3) <= VN325_sign_out(5);
    CN377_data_in(4) <= VN347_data_out(5);
    CN377_sign_in(4) <= VN347_sign_out(5);
    CN377_data_in(5) <= VN423_data_out(5);
    CN377_sign_in(5) <= VN423_sign_out(5);
    CN377_data_in(6) <= VN451_data_out(5);
    CN377_sign_in(6) <= VN451_sign_out(5);
    CN377_data_in(7) <= VN529_data_out(5);
    CN377_sign_in(7) <= VN529_sign_out(5);
    CN377_data_in(8) <= VN579_data_out(5);
    CN377_sign_in(8) <= VN579_sign_out(5);
    CN377_data_in(9) <= VN644_data_out(5);
    CN377_sign_in(9) <= VN644_sign_out(5);
    CN377_data_in(10) <= VN676_data_out(5);
    CN377_sign_in(10) <= VN676_sign_out(5);
    CN377_data_in(11) <= VN769_data_out(5);
    CN377_sign_in(11) <= VN769_sign_out(5);
    CN377_data_in(12) <= VN837_data_out(5);
    CN377_sign_in(12) <= VN837_sign_out(5);
    CN377_data_in(13) <= VN978_data_out(5);
    CN377_sign_in(13) <= VN978_sign_out(5);
    CN377_data_in(14) <= VN1013_data_out(5);
    CN377_sign_in(14) <= VN1013_sign_out(5);
    CN377_data_in(15) <= VN1131_data_out(5);
    CN377_sign_in(15) <= VN1131_sign_out(5);
    CN377_data_in(16) <= VN1181_data_out(5);
    CN377_sign_in(16) <= VN1181_sign_out(5);
    CN377_data_in(17) <= VN1269_data_out(5);
    CN377_sign_in(17) <= VN1269_sign_out(5);
    CN377_data_in(18) <= VN1321_data_out(5);
    CN377_sign_in(18) <= VN1321_sign_out(5);
    CN377_data_in(19) <= VN1341_data_out(5);
    CN377_sign_in(19) <= VN1341_sign_out(5);
    CN377_data_in(20) <= VN1424_data_out(5);
    CN377_sign_in(20) <= VN1424_sign_out(5);
    CN377_data_in(21) <= VN1445_data_out(5);
    CN377_sign_in(21) <= VN1445_sign_out(5);
    CN377_data_in(22) <= VN1481_data_out(5);
    CN377_sign_in(22) <= VN1481_sign_out(5);
    CN377_data_in(23) <= VN1574_data_out(5);
    CN377_sign_in(23) <= VN1574_sign_out(5);
    CN377_data_in(24) <= VN1644_data_out(5);
    CN377_sign_in(24) <= VN1644_sign_out(5);
    CN377_data_in(25) <= VN1654_data_out(5);
    CN377_sign_in(25) <= VN1654_sign_out(5);
    CN377_data_in(26) <= VN1697_data_out(5);
    CN377_sign_in(26) <= VN1697_sign_out(5);
    CN377_data_in(27) <= VN1723_data_out(5);
    CN377_sign_in(27) <= VN1723_sign_out(5);
    CN377_data_in(28) <= VN1758_data_out(5);
    CN377_sign_in(28) <= VN1758_sign_out(5);
    CN377_data_in(29) <= VN1851_data_out(5);
    CN377_sign_in(29) <= VN1851_sign_out(5);
    CN377_data_in(30) <= VN1861_data_out(5);
    CN377_sign_in(30) <= VN1861_sign_out(5);
    CN377_data_in(31) <= VN1904_data_out(5);
    CN377_sign_in(31) <= VN1904_sign_out(5);
    CN378_data_in(0) <= VN86_data_out(5);
    CN378_sign_in(0) <= VN86_sign_out(5);
    CN378_data_in(1) <= VN149_data_out(5);
    CN378_sign_in(1) <= VN149_sign_out(5);
    CN378_data_in(2) <= VN187_data_out(5);
    CN378_sign_in(2) <= VN187_sign_out(5);
    CN378_data_in(3) <= VN246_data_out(5);
    CN378_sign_in(3) <= VN246_sign_out(5);
    CN378_data_in(4) <= VN331_data_out(5);
    CN378_sign_in(4) <= VN331_sign_out(5);
    CN378_data_in(5) <= VN355_data_out(5);
    CN378_sign_in(5) <= VN355_sign_out(5);
    CN378_data_in(6) <= VN402_data_out(5);
    CN378_sign_in(6) <= VN402_sign_out(5);
    CN378_data_in(7) <= VN495_data_out(5);
    CN378_sign_in(7) <= VN495_sign_out(5);
    CN378_data_in(8) <= VN558_data_out(5);
    CN378_sign_in(8) <= VN558_sign_out(5);
    CN378_data_in(9) <= VN591_data_out(5);
    CN378_sign_in(9) <= VN591_sign_out(5);
    CN378_data_in(10) <= VN641_data_out(5);
    CN378_sign_in(10) <= VN641_sign_out(5);
    CN378_data_in(11) <= VN716_data_out(5);
    CN378_sign_in(11) <= VN716_sign_out(5);
    CN378_data_in(12) <= VN727_data_out(5);
    CN378_sign_in(12) <= VN727_sign_out(5);
    CN378_data_in(13) <= VN800_data_out(5);
    CN378_sign_in(13) <= VN800_sign_out(5);
    CN378_data_in(14) <= VN885_data_out(5);
    CN378_sign_in(14) <= VN885_sign_out(5);
    CN378_data_in(15) <= VN918_data_out(5);
    CN378_sign_in(15) <= VN918_sign_out(5);
    CN378_data_in(16) <= VN1000_data_out(5);
    CN378_sign_in(16) <= VN1000_sign_out(5);
    CN378_data_in(17) <= VN1049_data_out(5);
    CN378_sign_in(17) <= VN1049_sign_out(5);
    CN378_data_in(18) <= VN1102_data_out(5);
    CN378_sign_in(18) <= VN1102_sign_out(5);
    CN378_data_in(19) <= VN1153_data_out(5);
    CN378_sign_in(19) <= VN1153_sign_out(5);
    CN378_data_in(20) <= VN1198_data_out(5);
    CN378_sign_in(20) <= VN1198_sign_out(5);
    CN378_data_in(21) <= VN1256_data_out(5);
    CN378_sign_in(21) <= VN1256_sign_out(5);
    CN378_data_in(22) <= VN1375_data_out(5);
    CN378_sign_in(22) <= VN1375_sign_out(5);
    CN378_data_in(23) <= VN1399_data_out(5);
    CN378_sign_in(23) <= VN1399_sign_out(5);
    CN378_data_in(24) <= VN1430_data_out(5);
    CN378_sign_in(24) <= VN1430_sign_out(5);
    CN378_data_in(25) <= VN1488_data_out(5);
    CN378_sign_in(25) <= VN1488_sign_out(5);
    CN378_data_in(26) <= VN1527_data_out(5);
    CN378_sign_in(26) <= VN1527_sign_out(5);
    CN378_data_in(27) <= VN1553_data_out(5);
    CN378_sign_in(27) <= VN1553_sign_out(5);
    CN378_data_in(28) <= VN1657_data_out(5);
    CN378_sign_in(28) <= VN1657_sign_out(5);
    CN378_data_in(29) <= VN1709_data_out(5);
    CN378_sign_in(29) <= VN1709_sign_out(5);
    CN378_data_in(30) <= VN1923_data_out(5);
    CN378_sign_in(30) <= VN1923_sign_out(5);
    CN378_data_in(31) <= VN1928_data_out(5);
    CN378_sign_in(31) <= VN1928_sign_out(5);
    CN379_data_in(0) <= VN105_data_out(5);
    CN379_sign_in(0) <= VN105_sign_out(5);
    CN379_data_in(1) <= VN151_data_out(5);
    CN379_sign_in(1) <= VN151_sign_out(5);
    CN379_data_in(2) <= VN277_data_out(5);
    CN379_sign_in(2) <= VN277_sign_out(5);
    CN379_data_in(3) <= VN315_data_out(5);
    CN379_sign_in(3) <= VN315_sign_out(5);
    CN379_data_in(4) <= VN351_data_out(5);
    CN379_sign_in(4) <= VN351_sign_out(5);
    CN379_data_in(5) <= VN441_data_out(5);
    CN379_sign_in(5) <= VN441_sign_out(5);
    CN379_data_in(6) <= VN482_data_out(5);
    CN379_sign_in(6) <= VN482_sign_out(5);
    CN379_data_in(7) <= VN542_data_out(5);
    CN379_sign_in(7) <= VN542_sign_out(5);
    CN379_data_in(8) <= VN655_data_out(5);
    CN379_sign_in(8) <= VN655_sign_out(5);
    CN379_data_in(9) <= VN686_data_out(5);
    CN379_sign_in(9) <= VN686_sign_out(5);
    CN379_data_in(10) <= VN724_data_out(5);
    CN379_sign_in(10) <= VN724_sign_out(5);
    CN379_data_in(11) <= VN780_data_out(5);
    CN379_sign_in(11) <= VN780_sign_out(5);
    CN379_data_in(12) <= VN847_data_out(5);
    CN379_sign_in(12) <= VN847_sign_out(5);
    CN379_data_in(13) <= VN906_data_out(5);
    CN379_sign_in(13) <= VN906_sign_out(5);
    CN379_data_in(14) <= VN999_data_out(5);
    CN379_sign_in(14) <= VN999_sign_out(5);
    CN379_data_in(15) <= VN1052_data_out(5);
    CN379_sign_in(15) <= VN1052_sign_out(5);
    CN379_data_in(16) <= VN1079_data_out(5);
    CN379_sign_in(16) <= VN1079_sign_out(5);
    CN379_data_in(17) <= VN1122_data_out(5);
    CN379_sign_in(17) <= VN1122_sign_out(5);
    CN379_data_in(18) <= VN1174_data_out(5);
    CN379_sign_in(18) <= VN1174_sign_out(5);
    CN379_data_in(19) <= VN1275_data_out(5);
    CN379_sign_in(19) <= VN1275_sign_out(5);
    CN379_data_in(20) <= VN1356_data_out(5);
    CN379_sign_in(20) <= VN1356_sign_out(5);
    CN379_data_in(21) <= VN1388_data_out(5);
    CN379_sign_in(21) <= VN1388_sign_out(5);
    CN379_data_in(22) <= VN1410_data_out(5);
    CN379_sign_in(22) <= VN1410_sign_out(5);
    CN379_data_in(23) <= VN1460_data_out(5);
    CN379_sign_in(23) <= VN1460_sign_out(5);
    CN379_data_in(24) <= VN1555_data_out(5);
    CN379_sign_in(24) <= VN1555_sign_out(5);
    CN379_data_in(25) <= VN1648_data_out(5);
    CN379_sign_in(25) <= VN1648_sign_out(5);
    CN379_data_in(26) <= VN1716_data_out(5);
    CN379_sign_in(26) <= VN1716_sign_out(5);
    CN379_data_in(27) <= VN1722_data_out(5);
    CN379_sign_in(27) <= VN1722_sign_out(5);
    CN379_data_in(28) <= VN1777_data_out(5);
    CN379_sign_in(28) <= VN1777_sign_out(5);
    CN379_data_in(29) <= VN1880_data_out(5);
    CN379_sign_in(29) <= VN1880_sign_out(5);
    CN379_data_in(30) <= VN1979_data_out(5);
    CN379_sign_in(30) <= VN1979_sign_out(5);
    CN379_data_in(31) <= VN1984_data_out(5);
    CN379_sign_in(31) <= VN1984_sign_out(5);
    CN380_data_in(0) <= VN77_data_out(5);
    CN380_sign_in(0) <= VN77_sign_out(5);
    CN380_data_in(1) <= VN118_data_out(5);
    CN380_sign_in(1) <= VN118_sign_out(5);
    CN380_data_in(2) <= VN182_data_out(5);
    CN380_sign_in(2) <= VN182_sign_out(5);
    CN380_data_in(3) <= VN270_data_out(5);
    CN380_sign_in(3) <= VN270_sign_out(5);
    CN380_data_in(4) <= VN317_data_out(5);
    CN380_sign_in(4) <= VN317_sign_out(5);
    CN380_data_in(5) <= VN356_data_out(5);
    CN380_sign_in(5) <= VN356_sign_out(5);
    CN380_data_in(6) <= VN398_data_out(5);
    CN380_sign_in(6) <= VN398_sign_out(5);
    CN380_data_in(7) <= VN498_data_out(5);
    CN380_sign_in(7) <= VN498_sign_out(5);
    CN380_data_in(8) <= VN512_data_out(5);
    CN380_sign_in(8) <= VN512_sign_out(5);
    CN380_data_in(9) <= VN574_data_out(5);
    CN380_sign_in(9) <= VN574_sign_out(5);
    CN380_data_in(10) <= VN650_data_out(5);
    CN380_sign_in(10) <= VN650_sign_out(5);
    CN380_data_in(11) <= VN677_data_out(5);
    CN380_sign_in(11) <= VN677_sign_out(5);
    CN380_data_in(12) <= VN742_data_out(5);
    CN380_sign_in(12) <= VN742_sign_out(5);
    CN380_data_in(13) <= VN801_data_out(5);
    CN380_sign_in(13) <= VN801_sign_out(5);
    CN380_data_in(14) <= VN852_data_out(5);
    CN380_sign_in(14) <= VN852_sign_out(5);
    CN380_data_in(15) <= VN923_data_out(5);
    CN380_sign_in(15) <= VN923_sign_out(5);
    CN380_data_in(16) <= VN976_data_out(5);
    CN380_sign_in(16) <= VN976_sign_out(5);
    CN380_data_in(17) <= VN1036_data_out(5);
    CN380_sign_in(17) <= VN1036_sign_out(5);
    CN380_data_in(18) <= VN1171_data_out(5);
    CN380_sign_in(18) <= VN1171_sign_out(5);
    CN380_data_in(19) <= VN1248_data_out(5);
    CN380_sign_in(19) <= VN1248_sign_out(5);
    CN380_data_in(20) <= VN1316_data_out(5);
    CN380_sign_in(20) <= VN1316_sign_out(5);
    CN380_data_in(21) <= VN1358_data_out(5);
    CN380_sign_in(21) <= VN1358_sign_out(5);
    CN380_data_in(22) <= VN1403_data_out(5);
    CN380_sign_in(22) <= VN1403_sign_out(5);
    CN380_data_in(23) <= VN1446_data_out(5);
    CN380_sign_in(23) <= VN1446_sign_out(5);
    CN380_data_in(24) <= VN1507_data_out(5);
    CN380_sign_in(24) <= VN1507_sign_out(5);
    CN380_data_in(25) <= VN1510_data_out(5);
    CN380_sign_in(25) <= VN1510_sign_out(5);
    CN380_data_in(26) <= VN1559_data_out(5);
    CN380_sign_in(26) <= VN1559_sign_out(5);
    CN380_data_in(27) <= VN1587_data_out(5);
    CN380_sign_in(27) <= VN1587_sign_out(5);
    CN380_data_in(28) <= VN1674_data_out(5);
    CN380_sign_in(28) <= VN1674_sign_out(5);
    CN380_data_in(29) <= VN1713_data_out(5);
    CN380_sign_in(29) <= VN1713_sign_out(5);
    CN380_data_in(30) <= VN1721_data_out(5);
    CN380_sign_in(30) <= VN1721_sign_out(5);
    CN380_data_in(31) <= VN1808_data_out(5);
    CN380_sign_in(31) <= VN1808_sign_out(5);
    CN381_data_in(0) <= VN60_data_out(5);
    CN381_sign_in(0) <= VN60_sign_out(5);
    CN381_data_in(1) <= VN157_data_out(5);
    CN381_sign_in(1) <= VN157_sign_out(5);
    CN381_data_in(2) <= VN214_data_out(5);
    CN381_sign_in(2) <= VN214_sign_out(5);
    CN381_data_in(3) <= VN233_data_out(5);
    CN381_sign_in(3) <= VN233_sign_out(5);
    CN381_data_in(4) <= VN287_data_out(5);
    CN381_sign_in(4) <= VN287_sign_out(5);
    CN381_data_in(5) <= VN346_data_out(5);
    CN381_sign_in(5) <= VN346_sign_out(5);
    CN381_data_in(6) <= VN408_data_out(5);
    CN381_sign_in(6) <= VN408_sign_out(5);
    CN381_data_in(7) <= VN463_data_out(5);
    CN381_sign_in(7) <= VN463_sign_out(5);
    CN381_data_in(8) <= VN559_data_out(5);
    CN381_sign_in(8) <= VN559_sign_out(5);
    CN381_data_in(9) <= VN562_data_out(5);
    CN381_sign_in(9) <= VN562_sign_out(5);
    CN381_data_in(10) <= VN719_data_out(5);
    CN381_sign_in(10) <= VN719_sign_out(5);
    CN381_data_in(11) <= VN815_data_out(5);
    CN381_sign_in(11) <= VN815_sign_out(5);
    CN381_data_in(12) <= VN897_data_out(5);
    CN381_sign_in(12) <= VN897_sign_out(5);
    CN381_data_in(13) <= VN955_data_out(5);
    CN381_sign_in(13) <= VN955_sign_out(5);
    CN381_data_in(14) <= VN1133_data_out(5);
    CN381_sign_in(14) <= VN1133_sign_out(5);
    CN381_data_in(15) <= VN1219_data_out(5);
    CN381_sign_in(15) <= VN1219_sign_out(5);
    CN381_data_in(16) <= VN1245_data_out(5);
    CN381_sign_in(16) <= VN1245_sign_out(5);
    CN381_data_in(17) <= VN1344_data_out(5);
    CN381_sign_in(17) <= VN1344_sign_out(5);
    CN381_data_in(18) <= VN1407_data_out(5);
    CN381_sign_in(18) <= VN1407_sign_out(5);
    CN381_data_in(19) <= VN1476_data_out(5);
    CN381_sign_in(19) <= VN1476_sign_out(5);
    CN381_data_in(20) <= VN1501_data_out(5);
    CN381_sign_in(20) <= VN1501_sign_out(5);
    CN381_data_in(21) <= VN1568_data_out(5);
    CN381_sign_in(21) <= VN1568_sign_out(5);
    CN381_data_in(22) <= VN1643_data_out(5);
    CN381_sign_in(22) <= VN1643_sign_out(5);
    CN381_data_in(23) <= VN1695_data_out(5);
    CN381_sign_in(23) <= VN1695_sign_out(5);
    CN381_data_in(24) <= VN1719_data_out(5);
    CN381_sign_in(24) <= VN1719_sign_out(5);
    CN381_data_in(25) <= VN1729_data_out(5);
    CN381_sign_in(25) <= VN1729_sign_out(5);
    CN381_data_in(26) <= VN1751_data_out(5);
    CN381_sign_in(26) <= VN1751_sign_out(5);
    CN381_data_in(27) <= VN1779_data_out(5);
    CN381_sign_in(27) <= VN1779_sign_out(5);
    CN381_data_in(28) <= VN1781_data_out(5);
    CN381_sign_in(28) <= VN1781_sign_out(5);
    CN381_data_in(29) <= VN1849_data_out(5);
    CN381_sign_in(29) <= VN1849_sign_out(5);
    CN381_data_in(30) <= VN1855_data_out(5);
    CN381_sign_in(30) <= VN1855_sign_out(5);
    CN381_data_in(31) <= VN1905_data_out(5);
    CN381_sign_in(31) <= VN1905_sign_out(5);
    CN382_data_in(0) <= VN87_data_out(5);
    CN382_sign_in(0) <= VN87_sign_out(5);
    CN382_data_in(1) <= VN111_data_out(5);
    CN382_sign_in(1) <= VN111_sign_out(5);
    CN382_data_in(2) <= VN198_data_out(5);
    CN382_sign_in(2) <= VN198_sign_out(5);
    CN382_data_in(3) <= VN237_data_out(5);
    CN382_sign_in(3) <= VN237_sign_out(5);
    CN382_data_in(4) <= VN323_data_out(5);
    CN382_sign_in(4) <= VN323_sign_out(5);
    CN382_data_in(5) <= VN371_data_out(5);
    CN382_sign_in(5) <= VN371_sign_out(5);
    CN382_data_in(6) <= VN437_data_out(5);
    CN382_sign_in(6) <= VN437_sign_out(5);
    CN382_data_in(7) <= VN471_data_out(5);
    CN382_sign_in(7) <= VN471_sign_out(5);
    CN382_data_in(8) <= VN547_data_out(5);
    CN382_sign_in(8) <= VN547_sign_out(5);
    CN382_data_in(9) <= VN603_data_out(5);
    CN382_sign_in(9) <= VN603_sign_out(5);
    CN382_data_in(10) <= VN633_data_out(5);
    CN382_sign_in(10) <= VN633_sign_out(5);
    CN382_data_in(11) <= VN682_data_out(5);
    CN382_sign_in(11) <= VN682_sign_out(5);
    CN382_data_in(12) <= VN764_data_out(5);
    CN382_sign_in(12) <= VN764_sign_out(5);
    CN382_data_in(13) <= VN811_data_out(5);
    CN382_sign_in(13) <= VN811_sign_out(5);
    CN382_data_in(14) <= VN851_data_out(5);
    CN382_sign_in(14) <= VN851_sign_out(5);
    CN382_data_in(15) <= VN894_data_out(5);
    CN382_sign_in(15) <= VN894_sign_out(5);
    CN382_data_in(16) <= VN958_data_out(5);
    CN382_sign_in(16) <= VN958_sign_out(5);
    CN382_data_in(17) <= VN1033_data_out(5);
    CN382_sign_in(17) <= VN1033_sign_out(5);
    CN382_data_in(18) <= VN1091_data_out(5);
    CN382_sign_in(18) <= VN1091_sign_out(5);
    CN382_data_in(19) <= VN1124_data_out(5);
    CN382_sign_in(19) <= VN1124_sign_out(5);
    CN382_data_in(20) <= VN1178_data_out(5);
    CN382_sign_in(20) <= VN1178_sign_out(5);
    CN382_data_in(21) <= VN1260_data_out(5);
    CN382_sign_in(21) <= VN1260_sign_out(5);
    CN382_data_in(22) <= VN1324_data_out(5);
    CN382_sign_in(22) <= VN1324_sign_out(5);
    CN382_data_in(23) <= VN1331_data_out(5);
    CN382_sign_in(23) <= VN1331_sign_out(5);
    CN382_data_in(24) <= VN1376_data_out(5);
    CN382_sign_in(24) <= VN1376_sign_out(5);
    CN382_data_in(25) <= VN1396_data_out(5);
    CN382_sign_in(25) <= VN1396_sign_out(5);
    CN382_data_in(26) <= VN1562_data_out(5);
    CN382_sign_in(26) <= VN1562_sign_out(5);
    CN382_data_in(27) <= VN1588_data_out(5);
    CN382_sign_in(27) <= VN1588_sign_out(5);
    CN382_data_in(28) <= VN1628_data_out(5);
    CN382_sign_in(28) <= VN1628_sign_out(5);
    CN382_data_in(29) <= VN1708_data_out(5);
    CN382_sign_in(29) <= VN1708_sign_out(5);
    CN382_data_in(30) <= VN1720_data_out(5);
    CN382_sign_in(30) <= VN1720_sign_out(5);
    CN382_data_in(31) <= VN1809_data_out(5);
    CN382_sign_in(31) <= VN1809_sign_out(5);
    CN383_data_in(0) <= VN52_data_out(5);
    CN383_sign_in(0) <= VN52_sign_out(5);
    CN383_data_in(1) <= VN79_data_out(5);
    CN383_sign_in(1) <= VN79_sign_out(5);
    CN383_data_in(2) <= VN119_data_out(5);
    CN383_sign_in(2) <= VN119_sign_out(5);
    CN383_data_in(3) <= VN209_data_out(5);
    CN383_sign_in(3) <= VN209_sign_out(5);
    CN383_data_in(4) <= VN279_data_out(5);
    CN383_sign_in(4) <= VN279_sign_out(5);
    CN383_data_in(5) <= VN282_data_out(5);
    CN383_sign_in(5) <= VN282_sign_out(5);
    CN383_data_in(6) <= VN378_data_out(5);
    CN383_sign_in(6) <= VN378_sign_out(5);
    CN383_data_in(7) <= VN424_data_out(5);
    CN383_sign_in(7) <= VN424_sign_out(5);
    CN383_data_in(8) <= VN509_data_out(5);
    CN383_sign_in(8) <= VN509_sign_out(5);
    CN383_data_in(9) <= VN565_data_out(5);
    CN383_sign_in(9) <= VN565_sign_out(5);
    CN383_data_in(10) <= VN628_data_out(5);
    CN383_sign_in(10) <= VN628_sign_out(5);
    CN383_data_in(11) <= VN713_data_out(5);
    CN383_sign_in(11) <= VN713_sign_out(5);
    CN383_data_in(12) <= VN741_data_out(5);
    CN383_sign_in(12) <= VN741_sign_out(5);
    CN383_data_in(13) <= VN829_data_out(5);
    CN383_sign_in(13) <= VN829_sign_out(5);
    CN383_data_in(14) <= VN845_data_out(5);
    CN383_sign_in(14) <= VN845_sign_out(5);
    CN383_data_in(15) <= VN910_data_out(5);
    CN383_sign_in(15) <= VN910_sign_out(5);
    CN383_data_in(16) <= VN1001_data_out(5);
    CN383_sign_in(16) <= VN1001_sign_out(5);
    CN383_data_in(17) <= VN1003_data_out(5);
    CN383_sign_in(17) <= VN1003_sign_out(5);
    CN383_data_in(18) <= VN1089_data_out(5);
    CN383_sign_in(18) <= VN1089_sign_out(5);
    CN383_data_in(19) <= VN1209_data_out(5);
    CN383_sign_in(19) <= VN1209_sign_out(5);
    CN383_data_in(20) <= VN1254_data_out(5);
    CN383_sign_in(20) <= VN1254_sign_out(5);
    CN383_data_in(21) <= VN1294_data_out(5);
    CN383_sign_in(21) <= VN1294_sign_out(5);
    CN383_data_in(22) <= VN1340_data_out(5);
    CN383_sign_in(22) <= VN1340_sign_out(5);
    CN383_data_in(23) <= VN1513_data_out(5);
    CN383_sign_in(23) <= VN1513_sign_out(5);
    CN383_data_in(24) <= VN1565_data_out(5);
    CN383_sign_in(24) <= VN1565_sign_out(5);
    CN383_data_in(25) <= VN1597_data_out(5);
    CN383_sign_in(25) <= VN1597_sign_out(5);
    CN383_data_in(26) <= VN1633_data_out(5);
    CN383_sign_in(26) <= VN1633_sign_out(5);
    CN383_data_in(27) <= VN1680_data_out(5);
    CN383_sign_in(27) <= VN1680_sign_out(5);
    CN383_data_in(28) <= VN1750_data_out(5);
    CN383_sign_in(28) <= VN1750_sign_out(5);
    CN383_data_in(29) <= VN1775_data_out(5);
    CN383_sign_in(29) <= VN1775_sign_out(5);
    CN383_data_in(30) <= VN1882_data_out(5);
    CN383_sign_in(30) <= VN1882_sign_out(5);
    CN383_data_in(31) <= VN1914_data_out(5);
    CN383_sign_in(31) <= VN1914_sign_out(5);



end architecture ; -- arch