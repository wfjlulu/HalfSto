library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_signed.all;
--use ieee.std_logic_arith.all;  -- sysnopsys package not ieee standard
use ieee.numeric_std.all;
-- all numbers used are signed ?
-- (1723,2048) (6,32) regular RS-LDPC code
entity HalfStoTop is    -- the decoder lacks of early stop
  port (
    clk      : in std_logic;
    rst_n    : in std_logic;
    New_LLR    : in std_logic;
    RandomNum : in std_logic_vector( 3 downto 0);  -- not used , but for convenience , not modified
    LLR_in   : in std_logic_vector( 12287 downto 0 );   -- 6 bits quantity  2
    Codeword : inout std_logic_vector( 0 to 2047); -- 128*6 = 768 LLRs
    DV_out   : inout std_logic;                     -- 2048/128 = 16
    DecoderOver : inout std_logic;        -- one fram has been decoded over
    DecodeState : out std_logic_vector( 1 downto 0);
    Iterations  : inout std_logic_vector( 4 downto 0 )
    ) ;
end HalfStoTop ;

architecture arch of HalfStoTop is

    
    --signal : LLR0 std_logic_vector( 767 downto 0 );
    --signal : LLR1 std_logic_vector( 767 downto 0 );
    --signal : LLR2 std_logic_vector( 767 downto 0 );
    --signal : LLR3 std_logic_vector( 767 downto 0 );
    --signal : LLR4 std_logic_vector( 767 downto 0 );
    --signal : LLR5 std_logic_vector( 767 downto 0 );
    --signal : LLR6 std_logic_vector( 767 downto 0 );
    --signal : LLR7 std_logic_vector( 767 downto 0 );
    --signal : LLR8 std_logic_vector( 767 downto 0 );
    --signal : LLR9 std_logic_vector( 767 downto 0 );
    --signal : LLR10 std_logic_vector( 767 downto 0 );
    --signal : LLR11 std_logic_vector( 767 downto 0 );
    --signal : LLR12 std_logic_vector( 767 downto 0 );
    --signal : LLR13 std_logic_vector( 767 downto 0 );
    --signal : LLR14 std_logic_vector( 767 downto 0 );
    --signal : LLR15 std_logic_vector( 767 downto 0 );

    --signal : counter unsigned( 3 downto 0 );

    --signal VN_sign_out : std_logic_vector( 12287 downto 0);
    --signal VN_data_out : std_logic_vector( 12287 downto 0);

component CN2VN_wire is
    port(
        CN_data_out : in std_logic_vector(12287 downto 0);
        CN_sign_out : in std_logic_vector(12287 downto 0);
        VN_data_in : out std_logic_vector(12287 downto 0);
        VN_sign_in : out std_logic_vector(12287 downto 0)
    );
end component;

component VNUpdate is 
    port(
        clk :         in std_logic;
        rst_n :       in std_logic;
        LLR :         in std_logic_vector(12287 downto 0);  --2048*6 = 12288
        VN_data_in :  in std_logic_vector(12287 downto 0);--2048*6 = 12288
        VN_sign_in :  in std_logic_vector(12287 downto 0);
        RandomNum :   in std_logic_vector(3 downto 0);
        New_LLR   :   in std_logic;
        DecoderOver : in std_logic;
        --DV_in :       in std_logic;
        VN_data_out : out std_logic_vector(12287 downto 0);
        VN_sign_out : out std_logic_vector(12287 downto 0);
        codeword :    out std_logic_vector(0 to 2047);
        Iterations :  inout std_logic_vector(4 downto 0);
        DV_out :      out std_logic;
        DecodeState : out std_logic_vector( 1 downto 0 )
    );
end component;

component VN2CN_wire is
    port(
        VN_data_out : in std_logic_vector(12287 downto 0);
        VN_sign_out : in std_logic_vector(12287 downto 0);
        CN_data_in : out std_logic_vector(12287 downto 0);
        CN_sign_in : out std_logic_vector(12287 downto 0)
    );
end component;

component CNUpdate is
    port(
        rst_n : in std_logic;
        clk : in std_logic;
        CN_sign_in : in std_logic_vector( 12287 downto 0 ); -- 384 * 32 = 12288
        CN_data_in : in std_logic_vector( 12287 downto 0 );
        CN_sign_out : out std_logic_vector( 12287 downto 0 );
        CN_data_out : out std_logic_vector( 12287 downto 0 )
    );
end component;

--signal DecoderOver : std_logic;
--signal Codeword    : std_logic_vector( 0 to 2047 );
--signal DV_out : std_logic;

signal CN_data_out : std_logic_vector(12287 downto 0);
signal CN_sign_out : std_logic_vector(12287 downto 0);
signal VN_data_in : std_logic_vector(12287 downto 0);
signal VN_sign_in : std_logic_vector(12287 downto 0);
signal CN_data_in : std_logic_vector(12287 downto 0);
signal CN_sign_in : std_logic_vector(12287 downto 0);
signal VN_data_out : std_logic_vector(12287 downto 0);
signal VN_sign_out : std_logic_vector( 12287 downto 0 );

--signal Iterations : std_logic_vector(4 downto 0);
signal check : std_logic;
signal check0 : std_logic;
signal check1 : std_logic;
signal check2 : std_logic;
signal check3 : std_logic;
signal check4 : std_logic;
signal check5 : std_logic;
signal check6 : std_logic;
signal check7 : std_logic;
signal check8 : std_logic;
signal check9 : std_logic;
signal check10 : std_logic;
signal check11 : std_logic;
signal check12 : std_logic;
signal check13 : std_logic;
signal check14 : std_logic;
signal check15 : std_logic;
signal check16 : std_logic;
signal check17 : std_logic;
signal check18 : std_logic;
signal check19 : std_logic;
signal check20 : std_logic;
signal check21 : std_logic;
signal check22 : std_logic;
signal check23 : std_logic;
signal check24 : std_logic;
signal check25 : std_logic;
signal check26 : std_logic;
signal check27 : std_logic;
signal check28 : std_logic;
signal check29 : std_logic;
signal check30 : std_logic;
signal check31 : std_logic;
signal check32 : std_logic;
signal check33 : std_logic;
signal check34 : std_logic;
signal check35 : std_logic;
signal check36 : std_logic;
signal check37 : std_logic;
signal check38 : std_logic;
signal check39 : std_logic;
signal check40 : std_logic;
signal check41 : std_logic;
signal check42 : std_logic;
signal check43 : std_logic;
signal check44 : std_logic;
signal check45 : std_logic;
signal check46 : std_logic;
signal check47 : std_logic;
signal check48 : std_logic;
signal check49 : std_logic;
signal check50 : std_logic;
signal check51 : std_logic;
signal check52 : std_logic;
signal check53 : std_logic;
signal check54 : std_logic;
signal check55 : std_logic;
signal check56 : std_logic;
signal check57 : std_logic;
signal check58 : std_logic;
signal check59 : std_logic;
signal check60 : std_logic;
signal check61 : std_logic;
signal check62 : std_logic;
signal check63 : std_logic;
signal check64 : std_logic;
signal check65 : std_logic;
signal check66 : std_logic;
signal check67 : std_logic;
signal check68 : std_logic;
signal check69 : std_logic;
signal check70 : std_logic;
signal check71 : std_logic;
signal check72 : std_logic;
signal check73 : std_logic;
signal check74 : std_logic;
signal check75 : std_logic;
signal check76 : std_logic;
signal check77 : std_logic;
signal check78 : std_logic;
signal check79 : std_logic;
signal check80 : std_logic;
signal check81 : std_logic;
signal check82 : std_logic;
signal check83 : std_logic;
signal check84 : std_logic;
signal check85 : std_logic;
signal check86 : std_logic;
signal check87 : std_logic;
signal check88 : std_logic;
signal check89 : std_logic;
signal check90 : std_logic;
signal check91 : std_logic;
signal check92 : std_logic;
signal check93 : std_logic;
signal check94 : std_logic;
signal check95 : std_logic;
signal check96 : std_logic;
signal check97 : std_logic;
signal check98 : std_logic;
signal check99 : std_logic;
signal check100 : std_logic;
signal check101 : std_logic;
signal check102 : std_logic;
signal check103 : std_logic;
signal check104 : std_logic;
signal check105 : std_logic;
signal check106 : std_logic;
signal check107 : std_logic;
signal check108 : std_logic;
signal check109 : std_logic;
signal check110 : std_logic;
signal check111 : std_logic;
signal check112 : std_logic;
signal check113 : std_logic;
signal check114 : std_logic;
signal check115 : std_logic;
signal check116 : std_logic;
signal check117 : std_logic;
signal check118 : std_logic;
signal check119 : std_logic;
signal check120 : std_logic;
signal check121 : std_logic;
signal check122 : std_logic;
signal check123 : std_logic;
signal check124 : std_logic;
signal check125 : std_logic;
signal check126 : std_logic;
signal check127 : std_logic;
signal check128 : std_logic;
signal check129 : std_logic;
signal check130 : std_logic;
signal check131 : std_logic;
signal check132 : std_logic;
signal check133 : std_logic;
signal check134 : std_logic;
signal check135 : std_logic;
signal check136 : std_logic;
signal check137 : std_logic;
signal check138 : std_logic;
signal check139 : std_logic;
signal check140 : std_logic;
signal check141 : std_logic;
signal check142 : std_logic;
signal check143 : std_logic;
signal check144 : std_logic;
signal check145 : std_logic;
signal check146 : std_logic;
signal check147 : std_logic;
signal check148 : std_logic;
signal check149 : std_logic;
signal check150 : std_logic;
signal check151 : std_logic;
signal check152 : std_logic;
signal check153 : std_logic;
signal check154 : std_logic;
signal check155 : std_logic;
signal check156 : std_logic;
signal check157 : std_logic;
signal check158 : std_logic;
signal check159 : std_logic;
signal check160 : std_logic;
signal check161 : std_logic;
signal check162 : std_logic;
signal check163 : std_logic;
signal check164 : std_logic;
signal check165 : std_logic;
signal check166 : std_logic;
signal check167 : std_logic;
signal check168 : std_logic;
signal check169 : std_logic;
signal check170 : std_logic;
signal check171 : std_logic;
signal check172 : std_logic;
signal check173 : std_logic;
signal check174 : std_logic;
signal check175 : std_logic;
signal check176 : std_logic;
signal check177 : std_logic;
signal check178 : std_logic;
signal check179 : std_logic;
signal check180 : std_logic;
signal check181 : std_logic;
signal check182 : std_logic;
signal check183 : std_logic;
signal check184 : std_logic;
signal check185 : std_logic;
signal check186 : std_logic;
signal check187 : std_logic;
signal check188 : std_logic;
signal check189 : std_logic;
signal check190 : std_logic;
signal check191 : std_logic;
signal check192 : std_logic;
signal check193 : std_logic;
signal check194 : std_logic;
signal check195 : std_logic;
signal check196 : std_logic;
signal check197 : std_logic;
signal check198 : std_logic;
signal check199 : std_logic;
signal check200 : std_logic;
signal check201 : std_logic;
signal check202 : std_logic;
signal check203 : std_logic;
signal check204 : std_logic;
signal check205 : std_logic;
signal check206 : std_logic;
signal check207 : std_logic;
signal check208 : std_logic;
signal check209 : std_logic;
signal check210 : std_logic;
signal check211 : std_logic;
signal check212 : std_logic;
signal check213 : std_logic;
signal check214 : std_logic;
signal check215 : std_logic;
signal check216 : std_logic;
signal check217 : std_logic;
signal check218 : std_logic;
signal check219 : std_logic;
signal check220 : std_logic;
signal check221 : std_logic;
signal check222 : std_logic;
signal check223 : std_logic;
signal check224 : std_logic;
signal check225 : std_logic;
signal check226 : std_logic;
signal check227 : std_logic;
signal check228 : std_logic;
signal check229 : std_logic;
signal check230 : std_logic;
signal check231 : std_logic;
signal check232 : std_logic;
signal check233 : std_logic;
signal check234 : std_logic;
signal check235 : std_logic;
signal check236 : std_logic;
signal check237 : std_logic;
signal check238 : std_logic;
signal check239 : std_logic;
signal check240 : std_logic;
signal check241 : std_logic;
signal check242 : std_logic;
signal check243 : std_logic;
signal check244 : std_logic;
signal check245 : std_logic;
signal check246 : std_logic;
signal check247 : std_logic;
signal check248 : std_logic;
signal check249 : std_logic;
signal check250 : std_logic;
signal check251 : std_logic;
signal check252 : std_logic;
signal check253 : std_logic;
signal check254 : std_logic;
signal check255 : std_logic;
signal check256 : std_logic;
signal check257 : std_logic;
signal check258 : std_logic;
signal check259 : std_logic;
signal check260 : std_logic;
signal check261 : std_logic;
signal check262 : std_logic;
signal check263 : std_logic;
signal check264 : std_logic;
signal check265 : std_logic;
signal check266 : std_logic;
signal check267 : std_logic;
signal check268 : std_logic;
signal check269 : std_logic;
signal check270 : std_logic;
signal check271 : std_logic;
signal check272 : std_logic;
signal check273 : std_logic;
signal check274 : std_logic;
signal check275 : std_logic;
signal check276 : std_logic;
signal check277 : std_logic;
signal check278 : std_logic;
signal check279 : std_logic;
signal check280 : std_logic;
signal check281 : std_logic;
signal check282 : std_logic;
signal check283 : std_logic;
signal check284 : std_logic;
signal check285 : std_logic;
signal check286 : std_logic;
signal check287 : std_logic;
signal check288 : std_logic;
signal check289 : std_logic;
signal check290 : std_logic;
signal check291 : std_logic;
signal check292 : std_logic;
signal check293 : std_logic;
signal check294 : std_logic;
signal check295 : std_logic;
signal check296 : std_logic;
signal check297 : std_logic;
signal check298 : std_logic;
signal check299 : std_logic;
signal check300 : std_logic;
signal check301 : std_logic;
signal check302 : std_logic;
signal check303 : std_logic;
signal check304 : std_logic;
signal check305 : std_logic;
signal check306 : std_logic;
signal check307 : std_logic;
signal check308 : std_logic;
signal check309 : std_logic;
signal check310 : std_logic;
signal check311 : std_logic;
signal check312 : std_logic;
signal check313 : std_logic;
signal check314 : std_logic;
signal check315 : std_logic;
signal check316 : std_logic;
signal check317 : std_logic;
signal check318 : std_logic;
signal check319 : std_logic;
signal check320 : std_logic;
signal check321 : std_logic;
signal check322 : std_logic;
signal check323 : std_logic;
signal check324 : std_logic;
signal check325 : std_logic;
signal check326 : std_logic;
signal check327 : std_logic;
signal check328 : std_logic;
signal check329 : std_logic;
signal check330 : std_logic;
signal check331 : std_logic;
signal check332 : std_logic;
signal check333 : std_logic;
signal check334 : std_logic;
signal check335 : std_logic;
signal check336 : std_logic;
signal check337 : std_logic;
signal check338 : std_logic;
signal check339 : std_logic;
signal check340 : std_logic;
signal check341 : std_logic;
signal check342 : std_logic;
signal check343 : std_logic;
signal check344 : std_logic;
signal check345 : std_logic;
signal check346 : std_logic;
signal check347 : std_logic;
signal check348 : std_logic;
signal check349 : std_logic;
signal check350 : std_logic;
signal check351 : std_logic;
signal check352 : std_logic;
signal check353 : std_logic;
signal check354 : std_logic;
signal check355 : std_logic;
signal check356 : std_logic;
signal check357 : std_logic;
signal check358 : std_logic;
signal check359 : std_logic;
signal check360 : std_logic;
signal check361 : std_logic;
signal check362 : std_logic;
signal check363 : std_logic;
signal check364 : std_logic;
signal check365 : std_logic;
signal check366 : std_logic;
signal check367 : std_logic;
signal check368 : std_logic;
signal check369 : std_logic;
signal check370 : std_logic;
signal check371 : std_logic;
signal check372 : std_logic;
signal check373 : std_logic;
signal check374 : std_logic;
signal check375 : std_logic;
signal check376 : std_logic;
signal check377 : std_logic;
signal check378 : std_logic;
signal check379 : std_logic;
signal check380 : std_logic;
signal check381 : std_logic;
signal check382 : std_logic;
signal check383 : std_logic;

signal counter : unsigned( 1 downto 0 );
--signal counter2 : unsigned( 1 downto 0 );
--signal DecoderOver : std_logic;




begin

    ------------------------------------------------------------
    --load the LLRs , 16 clks, one clk 128 LLRs
    --process( rst_n, clk )
    --    begin
    --        if rst_n = '0' then
    --            counter <= "0000";
    --        elsif clk'event and clk = '1' then
    --            if DV_in = '1' then
    --                counter <= counter + 1;
    --                case counter is 
    --                    when "0000" => LLR0 <= LLR_in;
    --                    when "0001" => LLR1 <= LLR_in;
    --                    when "0010" => LLR2 <= LLR_in;
    --                    when "0011" => LLR3 <= LLR_in;
    --                    when "0100" => LLR4 <= LLR_in;
    --                    when "0101" => LLR5 <= LLR_in;
    --                    when "0110" => LLR6 <= LLR_in;
    --                    when "0111" => LLR7 <= LLR_in;
    --                    when "1000" => LLR8 <= LLR_in;
    --                    when "1001" => LLR9 <= LLR_in;
    --                    when "1010" => LLR10 <= LLR_in;
    --                    when "1011" => LLR11 <= LLR_in;
    --                    when "1100" => LLR12 <= LLR_in;
    --                    when "1101" => LLR13 <= LLR_in;
    --                    when "1110" => LLR14 <= LLR_in;
    --                    when "1111" => LLR15 <= LLR_in;
    --                end case;
    --            end if;
    --        end if;
    --end process;

    -----------------------------------------------------------
    -- 形参  =》 实参
    U_CN2VN_wire : CN2VN_wire port map(
        CN_data_out => CN_data_out,
        CN_sign_out => CN_sign_out,
        VN_data_in => VN_data_in,
        VN_sign_in => VN_sign_in       
    );

    U_VNUpdata : VNUpdate port map(
        clk => clk,
        rst_n => rst_n,
        LLR => LLR_in,
        VN_data_in => VN_data_in,
        VN_sign_in => VN_sign_in,
        RandomNum => RandomNum,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        --DV_in => DV_in,
        VN_data_out => VN_data_out,
        VN_sign_out => VN_sign_out,
        codeword => Codeword,
        Iterations => Iterations,
        DV_out => DV_out,
        DecodeState => DecodeState
    );

    U_VN2CN_wire : VN2CN_wire port map(
        VN_data_out => VN_data_out,
        VN_sign_out => VN_sign_out,
        CN_data_in => CN_data_in,
        CN_sign_in => CN_sign_in
    );

    U_CNUpdate : CNUpdate port map(
        rst_n => rst_n,
        clk => clk,
        CN_sign_in => CN_sign_in,
        CN_data_in => CN_data_in,
        CN_sign_out => CN_sign_out,
        CN_data_out => CN_data_out
    );

    -- codewore check  exa
    --check0 <= Codeword(83) xor Codeword(90).......;
    process( clk, rst_n )
    begin
        if( rst_n = '0') then
            NULL;
            --check <= '1';
            --DecoderOver <= '1';
        elsif( clk'event and clk = '1' ) then
            if( DV_out = '1' ) then
                check0 <= Codeword(53) xor Codeword(110) xor Codeword(170) xor Codeword(224) xor
                Codeword(279) xor Codeword(332) xor Codeword(447) xor Codeword(505) xor
                Codeword(616) xor Codeword(668) xor Codeword(1496) xor Codeword(1497) xor
                Codeword(1498) xor Codeword(1499) xor Codeword(1500) xor Codeword(1501) xor
                Codeword(1502) xor Codeword(1503) xor Codeword(1505) xor Codeword(1509) xor
                Codeword(1514) xor Codeword(1519) xor Codeword(1525) xor Codeword(1532) xor
                Codeword(1536) xor Codeword(1552) xor Codeword(1575) xor Codeword(1607) xor
                Codeword(1648) xor Codeword(1687) xor Codeword(1718) xor Codeword(1724);
 
     check1 <= Codeword(51) xor Codeword(139) xor Codeword(223) xor Codeword(241) xor
                Codeword(307) xor Codeword(356) xor Codeword(408) xor Codeword(476) xor
                Codeword(515) xor Codeword(600) xor Codeword(617) xor Codeword(689) xor
                Codeword(762) xor Codeword(797) xor Codeword(854) xor Codeword(927) xor
                Codeword(990) xor Codeword(1023) xor Codeword(1059) xor Codeword(1077) xor
                Codeword(1138) xor Codeword(1200) xor Codeword(1292) xor Codeword(1442) xor
                Codeword(1488) xor Codeword(1522) xor Codeword(1535) xor Codeword(1550) xor
                Codeword(1585) xor Codeword(1681) xor Codeword(1994) xor Codeword(1996);
 
     check2 <= Codeword(50) xor Codeword(92) xor Codeword(138) xor Codeword(222) xor
                Codeword(240) xor Codeword(306) xor Codeword(355) xor Codeword(407) xor
                Codeword(475) xor Codeword(599) xor Codeword(688) xor Codeword(761) xor
                Codeword(853) xor Codeword(989) xor Codeword(1003) xor Codeword(1022) xor
                Codeword(1076) xor Codeword(1137) xor Codeword(1199) xor Codeword(1291) xor
                Codeword(1441) xor Codeword(1521) xor Codeword(1534) xor Codeword(1549) xor
                Codeword(1584) xor Codeword(1707) xor Codeword(1808) xor Codeword(1837) xor
                Codeword(1904) xor Codeword(1948) xor Codeword(2003) xor Codeword(2007);
 
     check3 <= Codeword(91) xor Codeword(137) xor Codeword(221) xor Codeword(239) xor
                Codeword(305) xor Codeword(474) xor Codeword(514) xor Codeword(598) xor
                Codeword(687) xor Codeword(760) xor Codeword(796) xor Codeword(852) xor
                Codeword(926) xor Codeword(988) xor Codeword(1021) xor Codeword(1075) xor
                Codeword(1136) xor Codeword(1290) xor Codeword(1440) xor Codeword(1520) xor
                Codeword(1533) xor Codeword(1548) xor Codeword(1647) xor Codeword(1680) xor
                Codeword(1801) xor Codeword(1824) xor Codeword(1833) xor Codeword(1845) xor
                Codeword(1850) xor Codeword(1919) xor Codeword(1940) xor Codeword(1942);
 
     check4 <= Codeword(49) xor Codeword(90) xor Codeword(220) xor Codeword(238) xor
                Codeword(304) xor Codeword(354) xor Codeword(406) xor Codeword(473) xor
                Codeword(513) xor Codeword(597) xor Codeword(667) xor Codeword(686) xor
                Codeword(759) xor Codeword(795) xor Codeword(851) xor Codeword(887) xor
                Codeword(925) xor Codeword(987) xor Codeword(1074) xor Codeword(1135) xor
                Codeword(1198) xor Codeword(1289) xor Codeword(1583) xor Codeword(1646) xor
                Codeword(1679) xor Codeword(1747) xor Codeword(1892) xor Codeword(1901) xor
                Codeword(1907) xor Codeword(1944) xor Codeword(1977) xor Codeword(1978);
 
     check5 <= Codeword(48) xor Codeword(89) xor Codeword(136) xor Codeword(219) xor
                Codeword(237) xor Codeword(303) xor Codeword(353) xor Codeword(405) xor
                Codeword(472) xor Codeword(512) xor Codeword(596) xor Codeword(666) xor
                Codeword(685) xor Codeword(758) xor Codeword(794) xor Codeword(830) xor
                Codeword(850) xor Codeword(924) xor Codeword(986) xor Codeword(1020) xor
                Codeword(1073) xor Codeword(1134) xor Codeword(1197) xor Codeword(1275) xor
                Codeword(1288) xor Codeword(1383) xor Codeword(1439) xor Codeword(1547) xor
                Codeword(1582) xor Codeword(1645) xor Codeword(1678) xor Codeword(1725);
 
     check6 <= Codeword(47) xor Codeword(88) xor Codeword(135) xor Codeword(218) xor
                Codeword(236) xor Codeword(302) xor Codeword(352) xor Codeword(404) xor
                Codeword(471) xor Codeword(511) xor Codeword(595) xor Codeword(665) xor
                Codeword(684) xor Codeword(757) xor Codeword(777) xor Codeword(793) xor
                Codeword(849) xor Codeword(923) xor Codeword(985) xor Codeword(1019) xor
                Codeword(1072) xor Codeword(1133) xor Codeword(1196) xor Codeword(1274) xor
                Codeword(1287) xor Codeword(1382) xor Codeword(1438) xor Codeword(1546) xor
                Codeword(1581) xor Codeword(1644) xor Codeword(1706) xor Codeword(1726);
 
     check7 <= Codeword(46) xor Codeword(87) xor Codeword(134) xor Codeword(217) xor
                Codeword(235) xor Codeword(301) xor Codeword(351) xor Codeword(403) xor
                Codeword(470) xor Codeword(510) xor Codeword(594) xor Codeword(664) xor
                Codeword(683) xor Codeword(722) xor Codeword(756) xor Codeword(792) xor
                Codeword(848) xor Codeword(922) xor Codeword(984) xor Codeword(1018) xor
                Codeword(1071) xor Codeword(1132) xor Codeword(1195) xor Codeword(1273) xor
                Codeword(1286) xor Codeword(1381) xor Codeword(1437) xor Codeword(1545) xor
                Codeword(1580) xor Codeword(1677) xor Codeword(1705) xor Codeword(1727);
 
     check8 <= Codeword(45) xor Codeword(133) xor Codeword(216) xor Codeword(402) xor
                Codeword(469) xor Codeword(593) xor Codeword(682) xor Codeword(755) xor
                Codeword(847) xor Codeword(983) xor Codeword(1017) xor Codeword(1070) xor
                Codeword(1131) xor Codeword(1194) xor Codeword(1272) xor Codeword(1380) xor
                Codeword(1436) xor Codeword(1544) xor Codeword(1643) xor Codeword(1676) xor
                Codeword(1788) xor Codeword(1792) xor Codeword(1859) xor Codeword(1886) xor
                Codeword(1891) xor Codeword(1902) xor Codeword(1924) xor Codeword(1965) xor
                Codeword(1997) xor Codeword(2019) xor Codeword(2037) xor Codeword(2038);
 
     check9 <= Codeword(44) xor Codeword(86) xor Codeword(132) xor Codeword(215) xor
                Codeword(234) xor Codeword(300) xor Codeword(350) xor Codeword(391) xor
                Codeword(401) xor Codeword(468) xor Codeword(509) xor Codeword(592) xor
                Codeword(663) xor Codeword(681) xor Codeword(754) xor Codeword(791) xor
                Codeword(846) xor Codeword(921) xor Codeword(982) xor Codeword(1016) xor
                Codeword(1069) xor Codeword(1130) xor Codeword(1193) xor Codeword(1271) xor
                Codeword(1285) xor Codeword(1379) xor Codeword(1435) xor Codeword(1543) xor
                Codeword(1579) xor Codeword(1642) xor Codeword(1675) xor Codeword(1728);
 
     check10 <= Codeword(43) xor Codeword(85) xor Codeword(131) xor Codeword(233) xor
                Codeword(349) xor Codeword(467) xor Codeword(508) xor Codeword(662) xor
                Codeword(753) xor Codeword(790) xor Codeword(845) xor Codeword(920) xor
                Codeword(981) xor Codeword(1015) xor Codeword(1270) xor Codeword(1378) xor
                Codeword(1455) xor Codeword(1542) xor Codeword(1578) xor Codeword(1641) xor
                Codeword(1674) xor Codeword(1704) xor Codeword(1830) xor Codeword(1895) xor
                Codeword(1918) xor Codeword(1971) xor Codeword(1981) xor Codeword(1982) xor
                Codeword(1993) xor Codeword(2009) xor Codeword(2013) xor Codeword(2014);
 
     check11 <= Codeword(42) xor Codeword(84) xor Codeword(130) xor Codeword(214) xor
                Codeword(232) xor Codeword(348) xor Codeword(400) xor Codeword(591) xor
                Codeword(661) xor Codeword(680) xor Codeword(752) xor Codeword(789) xor
                Codeword(844) xor Codeword(919) xor Codeword(1014) xor Codeword(1068) xor
                Codeword(1129) xor Codeword(1269) xor Codeword(1434) xor Codeword(1454) xor
                Codeword(1541) xor Codeword(1577) xor Codeword(1640) xor Codeword(1673) xor
                Codeword(1764) xor Codeword(1829) xor Codeword(1843) xor Codeword(1860) xor
                Codeword(1867) xor Codeword(1914) xor Codeword(1946) xor Codeword(1951);
 
     check12 <= Codeword(41) xor Codeword(83) xor Codeword(129) xor Codeword(213) xor
                Codeword(231) xor Codeword(299) xor Codeword(347) xor Codeword(399) xor
                Codeword(466) xor Codeword(507) xor Codeword(590) xor Codeword(660) xor
                Codeword(679) xor Codeword(751) xor Codeword(788) xor Codeword(843) xor
                Codeword(918) xor Codeword(980) xor Codeword(1067) xor Codeword(1128) xor
                Codeword(1192) xor Codeword(1268) xor Codeword(1284) xor Codeword(1377) xor
                Codeword(1433) xor Codeword(1453) xor Codeword(1487) xor Codeword(1540) xor
                Codeword(1639) xor Codeword(1672) xor Codeword(1703) xor Codeword(1729);
 
     check13 <= Codeword(82) xor Codeword(128) xor Codeword(212) xor Codeword(230) xor
                Codeword(298) xor Codeword(346) xor Codeword(398) xor Codeword(465) xor
                Codeword(506) xor Codeword(589) xor Codeword(659) xor Codeword(678) xor
                Codeword(750) xor Codeword(787) xor Codeword(842) xor Codeword(917) xor
                Codeword(979) xor Codeword(1013) xor Codeword(1066) xor Codeword(1127) xor
                Codeword(1191) xor Codeword(1267) xor Codeword(1283) xor Codeword(1376) xor
                Codeword(1432) xor Codeword(1452) xor Codeword(1576) xor Codeword(1638) xor
                Codeword(1671) xor Codeword(1702) xor Codeword(1750) xor Codeword(1810);
 
     check14 <= Codeword(40) xor Codeword(81) xor Codeword(127) xor Codeword(211) xor
                Codeword(229) xor Codeword(297) xor Codeword(345) xor Codeword(397) xor
                Codeword(464) xor Codeword(560) xor Codeword(588) xor Codeword(658) xor
                Codeword(677) xor Codeword(749) xor Codeword(786) xor Codeword(841) xor
                Codeword(916) xor Codeword(978) xor Codeword(1012) xor Codeword(1065) xor
                Codeword(1126) xor Codeword(1190) xor Codeword(1266) xor Codeword(1375) xor
                Codeword(1431) xor Codeword(1451) xor Codeword(1486) xor Codeword(1531) xor
                Codeword(1539) xor Codeword(1637) xor Codeword(1778) xor Codeword(1811);
 
     check15 <= Codeword(39) xor Codeword(80) xor Codeword(126) xor Codeword(210) xor
                Codeword(228) xor Codeword(296) xor Codeword(344) xor Codeword(396) xor
                Codeword(559) xor Codeword(657) xor Codeword(785) xor Codeword(840) xor
                Codeword(915) xor Codeword(977) xor Codeword(1011) xor Codeword(1064) xor
                Codeword(1125) xor Codeword(1189) xor Codeword(1265) xor Codeword(1374) xor
                Codeword(1450) xor Codeword(1483) xor Codeword(1530) xor Codeword(1701) xor
                Codeword(1753) xor Codeword(1809) xor Codeword(1842) xor Codeword(1910) xor
                Codeword(1925) xor Codeword(1937) xor Codeword(1953) xor Codeword(1961);
 
     check16 <= Codeword(38) xor Codeword(125) xor Codeword(209) xor Codeword(227) xor
                Codeword(295) xor Codeword(343) xor Codeword(395) xor Codeword(463) xor
                Codeword(587) xor Codeword(656) xor Codeword(676) xor Codeword(748) xor
                Codeword(839) xor Codeword(976) xor Codeword(1010) xor Codeword(1063) xor
                Codeword(1124) xor Codeword(1188) xor Codeword(1264) xor Codeword(1373) xor
                Codeword(1430) xor Codeword(1482) xor Codeword(1529) xor Codeword(1538) xor
                Codeword(1636) xor Codeword(1670) xor Codeword(1700) xor Codeword(1900) xor
                Codeword(2006) xor Codeword(2023) xor Codeword(2034) xor Codeword(2036);
 
     check17 <= Codeword(37) xor Codeword(79) xor Codeword(124) xor Codeword(208) xor
                Codeword(226) xor Codeword(294) xor Codeword(342) xor Codeword(394) xor
                Codeword(462) xor Codeword(558) xor Codeword(586) xor Codeword(655) xor
                Codeword(675) xor Codeword(747) xor Codeword(784) xor Codeword(838) xor
                Codeword(914) xor Codeword(975) xor Codeword(1009) xor Codeword(1062) xor
                Codeword(1123) xor Codeword(1187) xor Codeword(1263) xor Codeword(1372) xor
                Codeword(1429) xor Codeword(1449) xor Codeword(1481) xor Codeword(1528) xor
                Codeword(1699) xor Codeword(1786) xor Codeword(1807) xor Codeword(1812);
 
     check18 <= Codeword(36) xor Codeword(78) xor Codeword(123) xor Codeword(207) xor
                Codeword(225) xor Codeword(293) xor Codeword(341) xor Codeword(393) xor
                Codeword(461) xor Codeword(557) xor Codeword(585) xor Codeword(654) xor
                Codeword(674) xor Codeword(746) xor Codeword(783) xor Codeword(837) xor
                Codeword(913) xor Codeword(974) xor Codeword(1008) xor Codeword(1061) xor
                Codeword(1122) xor Codeword(1186) xor Codeword(1262) xor Codeword(1371) xor
                Codeword(1428) xor Codeword(1448) xor Codeword(1480) xor Codeword(1527) xor
                Codeword(1537) xor Codeword(1635) xor Codeword(1698) xor Codeword(1730);
 
     check19 <= Codeword(35) xor Codeword(77) xor Codeword(122) xor Codeword(278) xor
                Codeword(340) xor Codeword(460) xor Codeword(556) xor Codeword(584) xor
                Codeword(745) xor Codeword(782) xor Codeword(836) xor Codeword(912) xor
                Codeword(973) xor Codeword(1261) xor Codeword(1370) xor Codeword(1447) xor
                Codeword(1479) xor Codeword(1526) xor Codeword(1634) xor Codeword(1669) xor
                Codeword(1697) xor Codeword(1772) xor Codeword(1849) xor Codeword(1884) xor
                Codeword(1885) xor Codeword(1957) xor Codeword(1964) xor Codeword(1986) xor
                Codeword(1989) xor Codeword(2028) xor Codeword(2041) xor Codeword(2042);
 
     check20 <= Codeword(34) xor Codeword(76) xor Codeword(277) xor Codeword(292) xor
                Codeword(339) xor Codeword(459) xor Codeword(555) xor Codeword(583) xor
                Codeword(673) xor Codeword(781) xor Codeword(911) xor Codeword(972) xor
                Codeword(1007) xor Codeword(1121) xor Codeword(1185) xor Codeword(1260) xor
                Codeword(1328) xor Codeword(1427) xor Codeword(1446) xor Codeword(1478) xor
                Codeword(1508) xor Codeword(1633) xor Codeword(1696) xor Codeword(1770) xor
                Codeword(1773) xor Codeword(1787) xor Codeword(1844) xor Codeword(1852) xor
                Codeword(1854) xor Codeword(1857) xor Codeword(1858) xor Codeword(1876);
 
     check21 <= Codeword(33) xor Codeword(75) xor Codeword(121) xor Codeword(206) xor
                Codeword(276) xor Codeword(291) xor Codeword(338) xor Codeword(392) xor
                Codeword(458) xor Codeword(554) xor Codeword(653) xor Codeword(672) xor
                Codeword(744) xor Codeword(780) xor Codeword(835) xor Codeword(910) xor
                Codeword(971) xor Codeword(1006) xor Codeword(1111) xor Codeword(1120) xor
                Codeword(1184) xor Codeword(1259) xor Codeword(1327) xor Codeword(1369) xor
                Codeword(1425) xor Codeword(1426) xor Codeword(1445) xor Codeword(1477) xor
                Codeword(1632) xor Codeword(1668) xor Codeword(1932) xor Codeword(1934);
 
     check22 <= Codeword(32) xor Codeword(74) xor Codeword(120) xor Codeword(205) xor
                Codeword(275) xor Codeword(290) xor Codeword(337) xor Codeword(446) xor
                Codeword(457) xor Codeword(582) xor Codeword(671) xor Codeword(743) xor
                Codeword(834) xor Codeword(970) xor Codeword(1119) xor Codeword(1183) xor
                Codeword(1258) xor Codeword(1326) xor Codeword(1368) xor Codeword(1390) xor
                Codeword(1424) xor Codeword(1507) xor Codeword(1631) xor Codeword(1765) xor
                Codeword(1793) xor Codeword(1795) xor Codeword(1882) xor Codeword(1903) xor
                Codeword(1941) xor Codeword(1987) xor Codeword(2032) xor Codeword(2035);
 
     check23 <= Codeword(31) xor Codeword(73) xor Codeword(119) xor Codeword(204) xor
                Codeword(274) xor Codeword(289) xor Codeword(336) xor Codeword(445) xor
                Codeword(456) xor Codeword(553) xor Codeword(581) xor Codeword(652) xor
                Codeword(742) xor Codeword(779) xor Codeword(833) xor Codeword(909) xor
                Codeword(969) xor Codeword(1005) xor Codeword(1109) xor Codeword(1118) xor
                Codeword(1182) xor Codeword(1257) xor Codeword(1325) xor Codeword(1367) xor
                Codeword(1389) xor Codeword(1423) xor Codeword(1444) xor Codeword(1476) xor
                Codeword(1630) xor Codeword(1754) xor Codeword(1802) xor Codeword(1813);
 
     check24 <= Codeword(30) xor Codeword(72) xor Codeword(118) xor Codeword(203) xor
                Codeword(273) xor Codeword(288) xor Codeword(335) xor Codeword(444) xor
                Codeword(455) xor Codeword(552) xor Codeword(580) xor Codeword(651) xor
                Codeword(670) xor Codeword(741) xor Codeword(778) xor Codeword(832) xor
                Codeword(908) xor Codeword(968) xor Codeword(1004) xor Codeword(1117) xor
                Codeword(1181) xor Codeword(1324) xor Codeword(1366) xor Codeword(1388) xor
                Codeword(1422) xor Codeword(1443) xor Codeword(1506) xor Codeword(1667) xor
                Codeword(1695) xor Codeword(1760) xor Codeword(1784) xor Codeword(1814);
 
     check25 <= Codeword(29) xor Codeword(71) xor Codeword(117) xor Codeword(202) xor
                Codeword(287) xor Codeword(443) xor Codeword(454) xor Codeword(551) xor
                Codeword(579) xor Codeword(650) xor Codeword(669) xor Codeword(740) xor
                Codeword(831) xor Codeword(907) xor Codeword(967) xor Codeword(1107) xor
                Codeword(1116) xor Codeword(1180) xor Codeword(1256) xor Codeword(1323) xor
                Codeword(1365) xor Codeword(1387) xor Codeword(1466) xor Codeword(1504) xor
                Codeword(1629) xor Codeword(1759) xor Codeword(1766) xor Codeword(1800) xor
                Codeword(1841) xor Codeword(1862) xor Codeword(1875) xor Codeword(1877);
 
     check26 <= Codeword(28) xor Codeword(70) xor Codeword(116) xor Codeword(201) xor
                Codeword(272) xor Codeword(286) xor Codeword(334) xor Codeword(442) xor
                Codeword(453) xor Codeword(550) xor Codeword(578) xor Codeword(649) xor
                Codeword(721) xor Codeword(739) xor Codeword(829) xor Codeword(886) xor
                Codeword(906) xor Codeword(966) xor Codeword(1058) xor Codeword(1106) xor
                Codeword(1115) xor Codeword(1179) xor Codeword(1255) xor Codeword(1322) xor
                Codeword(1364) xor Codeword(1386) xor Codeword(1421) xor Codeword(1465) xor
                Codeword(1558) xor Codeword(1666) xor Codeword(1694) xor Codeword(1731);
 
     check27 <= Codeword(27) xor Codeword(69) xor Codeword(115) xor Codeword(200) xor
                Codeword(285) xor Codeword(441) xor Codeword(452) xor Codeword(549) xor
                Codeword(648) xor Codeword(720) xor Codeword(738) xor Codeword(828) xor
                Codeword(885) xor Codeword(905) xor Codeword(965) xor Codeword(1057) xor
                Codeword(1105) xor Codeword(1178) xor Codeword(1321) xor Codeword(1385) xor
                Codeword(1420) xor Codeword(1464) xor Codeword(1557) xor Codeword(1665) xor
                Codeword(1769) xor Codeword(1780) xor Codeword(1828) xor Codeword(1839) xor
                Codeword(1848) xor Codeword(1869) xor Codeword(1933) xor Codeword(1935);
 
     check28 <= Codeword(26) xor Codeword(68) xor Codeword(114) xor Codeword(199) xor
                Codeword(271) xor Codeword(333) xor Codeword(440) xor Codeword(451) xor
                Codeword(548) xor Codeword(577) xor Codeword(647) xor Codeword(719) xor
                Codeword(737) xor Codeword(827) xor Codeword(884) xor Codeword(904) xor
                Codeword(964) xor Codeword(1056) xor Codeword(1104) xor Codeword(1114) xor
                Codeword(1177) xor Codeword(1254) xor Codeword(1320) xor Codeword(1363) xor
                Codeword(1384) xor Codeword(1419) xor Codeword(1463) xor Codeword(1556) xor
                Codeword(1628) xor Codeword(1664) xor Codeword(1693) xor Codeword(1732);
 
     check29 <= Codeword(25) xor Codeword(67) xor Codeword(113) xor Codeword(270) xor
                Codeword(450) xor Codeword(547) xor Codeword(576) xor Codeword(646) xor
                Codeword(883) xor Codeword(903) xor Codeword(1055) xor Codeword(1103) xor
                Codeword(1253) xor Codeword(1319) xor Codeword(1362) xor Codeword(1418) xor
                Codeword(1462) xor Codeword(1555) xor Codeword(1627) xor Codeword(1758) xor
                Codeword(1781) xor Codeword(1803) xor Codeword(1894) xor Codeword(1898) xor
                Codeword(1913) xor Codeword(1922) xor Codeword(1955) xor Codeword(1960) xor
                Codeword(1980) xor Codeword(1985) xor Codeword(1988) xor Codeword(1990);
 
     check30 <= Codeword(24) xor Codeword(66) xor Codeword(112) xor Codeword(198) xor
                Codeword(269) xor Codeword(284) xor Codeword(390) xor Codeword(439) xor
                Codeword(449) xor Codeword(546) xor Codeword(575) xor Codeword(645) xor
                Codeword(718) xor Codeword(736) xor Codeword(882) xor Codeword(902) xor
                Codeword(963) xor Codeword(1054) xor Codeword(1102) xor Codeword(1176) xor
                Codeword(1252) xor Codeword(1318) xor Codeword(1334) xor Codeword(1361) xor
                Codeword(1417) xor Codeword(1461) xor Codeword(1513) xor Codeword(1663) xor
                Codeword(1692) xor Codeword(1771) xor Codeword(1806) xor Codeword(1815);
 
     check31 <= Codeword(23) xor Codeword(65) xor Codeword(197) xor Codeword(283) xor
                Codeword(389) xor Codeword(438) xor Codeword(448) xor Codeword(545) xor
                Codeword(574) xor Codeword(644) xor Codeword(717) xor Codeword(735) xor
                Codeword(826) xor Codeword(881) xor Codeword(901) xor Codeword(962) xor
                Codeword(1053) xor Codeword(1101) xor Codeword(1175) xor Codeword(1251) xor
                Codeword(1317) xor Codeword(1333) xor Codeword(1360) xor Codeword(1416) xor
                Codeword(1460) xor Codeword(1554) xor Codeword(1626) xor Codeword(1782) xor
                Codeword(1790) xor Codeword(1921) xor Codeword(1952) xor Codeword(1962);
 
     check32 <= Codeword(22) xor Codeword(64) xor Codeword(111) xor Codeword(268) xor
                Codeword(388) xor Codeword(504) xor Codeword(544) xor Codeword(573) xor
                Codeword(643) xor Codeword(734) xor Codeword(825) xor Codeword(880) xor
                Codeword(900) xor Codeword(961) xor Codeword(1052) xor Codeword(1250) xor
                Codeword(1316) xor Codeword(1359) xor Codeword(1459) xor Codeword(1662) xor
                Codeword(1691) xor Codeword(1742) xor Codeword(1826) xor Codeword(1831) xor
                Codeword(1943) xor Codeword(1958) xor Codeword(1959) xor Codeword(1973) xor
                Codeword(1999) xor Codeword(2008) xor Codeword(2027) xor Codeword(2029);
 
     check33 <= Codeword(21) xor Codeword(63) xor Codeword(169) xor Codeword(196) xor
                Codeword(267) xor Codeword(282) xor Codeword(387) xor Codeword(437) xor
                Codeword(503) xor Codeword(543) xor Codeword(572) xor Codeword(642) xor
                Codeword(716) xor Codeword(733) xor Codeword(824) xor Codeword(879) xor
                Codeword(899) xor Codeword(960) xor Codeword(1051) xor Codeword(1100) xor
                Codeword(1174) xor Codeword(1249) xor Codeword(1315) xor Codeword(1332) xor
                Codeword(1358) xor Codeword(1415) xor Codeword(1458) xor Codeword(1512) xor
                Codeword(1574) xor Codeword(1625) xor Codeword(1690) xor Codeword(1733);
 
     check34 <= Codeword(20) xor Codeword(62) xor Codeword(168) xor Codeword(195) xor
                Codeword(266) xor Codeword(281) xor Codeword(386) xor Codeword(436) xor
                Codeword(502) xor Codeword(542) xor Codeword(571) xor Codeword(641) xor
                Codeword(715) xor Codeword(732) xor Codeword(823) xor Codeword(878) xor
                Codeword(898) xor Codeword(959) xor Codeword(1050) xor Codeword(1099) xor
                Codeword(1173) xor Codeword(1248) xor Codeword(1314) xor Codeword(1331) xor
                Codeword(1414) xor Codeword(1511) xor Codeword(1573) xor Codeword(1606) xor
                Codeword(1624) xor Codeword(1661) xor Codeword(1822) xor Codeword(1878);
 
     check35 <= Codeword(19) xor Codeword(61) xor Codeword(167) xor Codeword(194) xor
                Codeword(265) xor Codeword(280) xor Codeword(385) xor Codeword(435) xor
                Codeword(501) xor Codeword(541) xor Codeword(570) xor Codeword(640) xor
                Codeword(714) xor Codeword(731) xor Codeword(822) xor Codeword(877) xor
                Codeword(897) xor Codeword(958) xor Codeword(1049) xor Codeword(1098) xor
                Codeword(1172) xor Codeword(1247) xor Codeword(1313) xor Codeword(1330) xor
                Codeword(1357) xor Codeword(1413) xor Codeword(1510) xor Codeword(1605) xor
                Codeword(1623) xor Codeword(1660) xor Codeword(1689) xor Codeword(1734);
 
     check36 <= Codeword(18) xor Codeword(60) xor Codeword(166) xor Codeword(264) xor
                Codeword(384) xor Codeword(434) xor Codeword(500) xor Codeword(540) xor
                Codeword(639) xor Codeword(821) xor Codeword(896) xor Codeword(957) xor
                Codeword(1048) xor Codeword(1171) xor Codeword(1246) xor Codeword(1329) xor
                Codeword(1356) xor Codeword(1412) xor Codeword(1604) xor Codeword(1622) xor
                Codeword(1659) xor Codeword(1743) xor Codeword(1873) xor Codeword(1888) xor
                Codeword(1947) xor Codeword(1950) xor Codeword(1969) xor Codeword(1976) xor
                Codeword(1995) xor Codeword(2002) xor Codeword(2022) xor Codeword(2030);
 
     check37 <= Codeword(17) xor Codeword(59) xor Codeword(165) xor Codeword(193) xor
                Codeword(263) xor Codeword(331) xor Codeword(383) xor Codeword(433) xor
                Codeword(499) xor Codeword(539) xor Codeword(569) xor Codeword(638) xor
                Codeword(713) xor Codeword(730) xor Codeword(820) xor Codeword(876) xor
                Codeword(895) xor Codeword(956) xor Codeword(1047) xor Codeword(1097) xor
                Codeword(1163) xor Codeword(1170) xor Codeword(1245) xor Codeword(1282) xor
                Codeword(1312) xor Codeword(1355) xor Codeword(1572) xor Codeword(1603) xor
                Codeword(1621) xor Codeword(1658) xor Codeword(1688) xor Codeword(1735);
 
     check38 <= Codeword(16) xor Codeword(58) xor Codeword(164) xor Codeword(192) xor
                Codeword(262) xor Codeword(330) xor Codeword(382) xor Codeword(432) xor
                Codeword(498) xor Codeword(538) xor Codeword(568) xor Codeword(637) xor
                Codeword(712) xor Codeword(729) xor Codeword(875) xor Codeword(894) xor
                Codeword(955) xor Codeword(1046) xor Codeword(1096) xor Codeword(1162) xor
                Codeword(1244) xor Codeword(1281) xor Codeword(1311) xor Codeword(1411) xor
                Codeword(1518) xor Codeword(1571) xor Codeword(1620) xor Codeword(1767) xor
                Codeword(1881) xor Codeword(1897) xor Codeword(1909) xor Codeword(1915);
 
     check39 <= Codeword(15) xor Codeword(57) xor Codeword(163) xor Codeword(191) xor
                Codeword(261) xor Codeword(329) xor Codeword(381) xor Codeword(431) xor
                Codeword(497) xor Codeword(537) xor Codeword(567) xor Codeword(636) xor
                Codeword(711) xor Codeword(728) xor Codeword(819) xor Codeword(874) xor
                Codeword(893) xor Codeword(954) xor Codeword(1045) xor Codeword(1095) xor
                Codeword(1161) xor Codeword(1243) xor Codeword(1280) xor Codeword(1310) xor
                Codeword(1354) xor Codeword(1410) xor Codeword(1517) xor Codeword(1570) xor
                Codeword(1602) xor Codeword(1619) xor Codeword(1657) xor Codeword(1736);
 
     check40 <= Codeword(14) xor Codeword(56) xor Codeword(162) xor Codeword(260) xor
                Codeword(380) xor Codeword(430) xor Codeword(496) xor Codeword(536) xor
                Codeword(566) xor Codeword(635) xor Codeword(727) xor Codeword(818) xor
                Codeword(873) xor Codeword(892) xor Codeword(953) xor Codeword(1044) xor
                Codeword(1160) xor Codeword(1242) xor Codeword(1279) xor Codeword(1353) xor
                Codeword(1409) xor Codeword(1569) xor Codeword(1601) xor Codeword(1618) xor
                Codeword(1656) xor Codeword(1717) xor Codeword(1856) xor Codeword(1912) xor
                Codeword(1974) xor Codeword(1984) xor Codeword(1991) xor Codeword(1992);
 
     check41 <= Codeword(13) xor Codeword(55) xor Codeword(161) xor Codeword(190) xor
                Codeword(259) xor Codeword(328) xor Codeword(379) xor Codeword(429) xor
                Codeword(495) xor Codeword(535) xor Codeword(565) xor Codeword(634) xor
                Codeword(710) xor Codeword(726) xor Codeword(817) xor Codeword(872) xor
                Codeword(891) xor Codeword(952) xor Codeword(1043) xor Codeword(1094) xor
                Codeword(1159) xor Codeword(1278) xor Codeword(1309) xor Codeword(1352) xor
                Codeword(1408) xor Codeword(1568) xor Codeword(1600) xor Codeword(1617) xor
                Codeword(1716) xor Codeword(1748) xor Codeword(1755) xor Codeword(1816);
 
     check42 <= Codeword(12) xor Codeword(54) xor Codeword(160) xor Codeword(189) xor
                Codeword(258) xor Codeword(327) xor Codeword(378) xor Codeword(428) xor
                Codeword(494) xor Codeword(534) xor Codeword(564) xor Codeword(633) xor
                Codeword(709) xor Codeword(725) xor Codeword(816) xor Codeword(871) xor
                Codeword(890) xor Codeword(951) xor Codeword(1042) xor Codeword(1093) xor
                Codeword(1158) xor Codeword(1241) xor Codeword(1308) xor Codeword(1351) xor
                Codeword(1407) xor Codeword(1516) xor Codeword(1553) xor Codeword(1567) xor
                Codeword(1616) xor Codeword(1655) xor Codeword(1715) xor Codeword(1737);
 
     check43 <= Codeword(109) xor Codeword(159) xor Codeword(188) xor Codeword(257) xor
                Codeword(326) xor Codeword(377) xor Codeword(427) xor Codeword(493) xor
                Codeword(533) xor Codeword(563) xor Codeword(632) xor Codeword(708) xor
                Codeword(815) xor Codeword(870) xor Codeword(889) xor Codeword(950) xor
                Codeword(1041) xor Codeword(1092) xor Codeword(1157) xor Codeword(1277) xor
                Codeword(1307) xor Codeword(1350) xor Codeword(1406) xor Codeword(1515) xor
                Codeword(1566) xor Codeword(1599) xor Codeword(1615) xor Codeword(1654) xor
                Codeword(1749) xor Codeword(1762) xor Codeword(1889) xor Codeword(1906);
 
     check44 <= Codeword(11) xor Codeword(108) xor Codeword(158) xor Codeword(187) xor
                Codeword(256) xor Codeword(325) xor Codeword(376) xor Codeword(426) xor
                Codeword(492) xor Codeword(532) xor Codeword(562) xor Codeword(631) xor
                Codeword(707) xor Codeword(724) xor Codeword(814) xor Codeword(869) xor
                Codeword(888) xor Codeword(949) xor Codeword(1040) xor Codeword(1091) xor
                Codeword(1156) xor Codeword(1217) xor Codeword(1240) xor Codeword(1276) xor
                Codeword(1306) xor Codeword(1349) xor Codeword(1405) xor Codeword(1565) xor
                Codeword(1598) xor Codeword(1614) xor Codeword(1714) xor Codeword(1738);
 
     check45 <= Codeword(10) xor Codeword(107) xor Codeword(157) xor Codeword(186) xor
                Codeword(255) xor Codeword(324) xor Codeword(375) xor Codeword(425) xor
                Codeword(491) xor Codeword(531) xor Codeword(561) xor Codeword(630) xor
                Codeword(706) xor Codeword(723) xor Codeword(813) xor Codeword(868) xor
                Codeword(943) xor Codeword(948) xor Codeword(1039) xor Codeword(1090) xor
                Codeword(1155) xor Codeword(1216) xor Codeword(1224) xor Codeword(1305) xor
                Codeword(1348) xor Codeword(1404) xor Codeword(1564) xor Codeword(1597) xor
                Codeword(1653) xor Codeword(1713) xor Codeword(1756) xor Codeword(1817);
 
     check46 <= Codeword(9) xor Codeword(106) xor Codeword(156) xor Codeword(185) xor
                Codeword(254) xor Codeword(323) xor Codeword(374) xor Codeword(424) xor
                Codeword(490) xor Codeword(530) xor Codeword(615) xor Codeword(705) xor
                Codeword(776) xor Codeword(812) xor Codeword(867) xor Codeword(947) xor
                Codeword(1038) xor Codeword(1154) xor Codeword(1215) xor Codeword(1223) xor
                Codeword(1239) xor Codeword(1304) xor Codeword(1347) xor Codeword(1403) xor
                Codeword(1563) xor Codeword(1596) xor Codeword(1613) xor Codeword(1791) xor
                Codeword(1825) xor Codeword(1832) xor Codeword(1861) xor Codeword(1879);
 
     check47 <= Codeword(8) xor Codeword(155) xor Codeword(253) xor Codeword(373) xor
                Codeword(489) xor Codeword(529) xor Codeword(614) xor Codeword(629) xor
                Codeword(811) xor Codeword(942) xor Codeword(946) xor Codeword(1037) xor
                Codeword(1222) xor Codeword(1238) xor Codeword(1346) xor Codeword(1402) xor
                Codeword(1612) xor Codeword(1652) xor Codeword(1741) xor Codeword(1746) xor
                Codeword(1893) xor Codeword(1896) xor Codeword(1899) xor Codeword(1923) xor
                Codeword(1956) xor Codeword(1968) xor Codeword(2001) xor Codeword(2020) xor
                Codeword(2021) xor Codeword(2033) xor Codeword(2044) xor Codeword(2045);
 
     check48 <= Codeword(7) xor Codeword(154) xor Codeword(322) xor Codeword(372) xor
                Codeword(423) xor Codeword(488) xor Codeword(528) xor Codeword(613) xor
                Codeword(704) xor Codeword(775) xor Codeword(810) xor Codeword(941) xor
                Codeword(945) xor Codeword(1036) xor Codeword(1089) xor Codeword(1153) xor
                Codeword(1221) xor Codeword(1237) xor Codeword(1345) xor Codeword(1401) xor
                Codeword(1562) xor Codeword(1595) xor Codeword(1763) xor Codeword(1796) xor
                Codeword(1823) xor Codeword(1887) xor Codeword(1911) xor Codeword(1938) xor
                Codeword(1954) xor Codeword(1979) xor Codeword(2004) xor Codeword(2005);
 
     check49 <= Codeword(6) xor Codeword(105) xor Codeword(153) xor Codeword(184) xor
                Codeword(252) xor Codeword(321) xor Codeword(371) xor Codeword(422) xor
                Codeword(487) xor Codeword(527) xor Codeword(612) xor Codeword(628) xor
                Codeword(703) xor Codeword(774) xor Codeword(809) xor Codeword(866) xor
                Codeword(940) xor Codeword(944) xor Codeword(1035) xor Codeword(1088) xor
                Codeword(1152) xor Codeword(1214) xor Codeword(1220) xor Codeword(1236) xor
                Codeword(1303) xor Codeword(1344) xor Codeword(1400) xor Codeword(1561) xor
                Codeword(1594) xor Codeword(1611) xor Codeword(1651) xor Codeword(1739);
 
     check50 <= Codeword(5) xor Codeword(104) xor Codeword(152) xor Codeword(183) xor
                Codeword(251) xor Codeword(320) xor Codeword(370) xor Codeword(421) xor
                Codeword(486) xor Codeword(526) xor Codeword(611) xor Codeword(627) xor
                Codeword(702) xor Codeword(773) xor Codeword(808) xor Codeword(865) xor
                Codeword(939) xor Codeword(1002) xor Codeword(1034) xor Codeword(1151) xor
                Codeword(1213) xor Codeword(1219) xor Codeword(1235) xor Codeword(1302) xor
                Codeword(1343) xor Codeword(1399) xor Codeword(1560) xor Codeword(1593) xor
                Codeword(1610) xor Codeword(1712) xor Codeword(1777) xor Codeword(1818);
 
     check51 <= Codeword(4) xor Codeword(103) xor Codeword(182) xor Codeword(250) xor
                Codeword(319) xor Codeword(369) xor Codeword(420) xor Codeword(485) xor
                Codeword(525) xor Codeword(610) xor Codeword(626) xor Codeword(701) xor
                Codeword(807) xor Codeword(938) xor Codeword(1001) xor Codeword(1087) xor
                Codeword(1150) xor Codeword(1218) xor Codeword(1342) xor Codeword(1398) xor
                Codeword(1457) xor Codeword(1592) xor Codeword(1609) xor Codeword(1834) xor
                Codeword(1835) xor Codeword(1864) xor Codeword(1866) xor Codeword(1868) xor
                Codeword(1926) xor Codeword(1939) xor Codeword(1998) xor Codeword(2000);
 
     check52 <= Codeword(102) xor Codeword(151) xor Codeword(181) xor Codeword(318) xor
                Codeword(368) xor Codeword(419) xor Codeword(524) xor Codeword(609) xor
                Codeword(625) xor Codeword(700) xor Codeword(772) xor Codeword(806) xor
                Codeword(864) xor Codeword(937) xor Codeword(1000) xor Codeword(1033) xor
                Codeword(1086) xor Codeword(1149) xor Codeword(1169) xor Codeword(1212) xor
                Codeword(1234) xor Codeword(1301) xor Codeword(1341) xor Codeword(1397) xor
                Codeword(1559) xor Codeword(1711) xor Codeword(1872) xor Codeword(1908) xor
                Codeword(1916) xor Codeword(1945) xor Codeword(2024) xor Codeword(2026);
 
     check53 <= Codeword(3) xor Codeword(150) xor Codeword(180) xor Codeword(249) xor
                Codeword(317) xor Codeword(367) xor Codeword(418) xor Codeword(484) xor
                Codeword(608) xor Codeword(699) xor Codeword(771) xor Codeword(863) xor
                Codeword(936) xor Codeword(1032) xor Codeword(1085) xor Codeword(1148) xor
                Codeword(1168) xor Codeword(1211) xor Codeword(1233) xor Codeword(1340) xor
                Codeword(1396) xor Codeword(1456) xor Codeword(1650) xor Codeword(1776) xor
                Codeword(1836) xor Codeword(1905) xor Codeword(1917) xor Codeword(1930) xor
                Codeword(2025) xor Codeword(2031) xor Codeword(2046) xor Codeword(2047);
 
     check54 <= Codeword(2) xor Codeword(101) xor Codeword(149) xor Codeword(179) xor
                Codeword(316) xor Codeword(366) xor Codeword(417) xor Codeword(523) xor
                Codeword(698) xor Codeword(770) xor Codeword(805) xor Codeword(862) xor
                Codeword(935) xor Codeword(999) xor Codeword(1031) xor Codeword(1084) xor
                Codeword(1147) xor Codeword(1210) xor Codeword(1232) xor Codeword(1300) xor
                Codeword(1339) xor Codeword(1475) xor Codeword(1608) xor Codeword(1649) xor
                Codeword(1752) xor Codeword(1785) xor Codeword(1797) xor Codeword(1840) xor
                Codeword(1847) xor Codeword(1890) xor Codeword(1931) xor Codeword(1936);
 
     check55 <= Codeword(1) xor Codeword(100) xor Codeword(148) xor Codeword(178) xor
                Codeword(248) xor Codeword(315) xor Codeword(365) xor Codeword(416) xor
                Codeword(483) xor Codeword(522) xor Codeword(607) xor Codeword(624) xor
                Codeword(697) xor Codeword(769) xor Codeword(804) xor Codeword(861) xor
                Codeword(934) xor Codeword(998) xor Codeword(1030) xor Codeword(1083) xor
                Codeword(1146) xor Codeword(1167) xor Codeword(1209) xor Codeword(1231) xor
                Codeword(1299) xor Codeword(1338) xor Codeword(1395) xor Codeword(1474) xor
                Codeword(1494) xor Codeword(1591) xor Codeword(1710) xor Codeword(1740);
 
     check56 <= Codeword(0) xor Codeword(99) xor Codeword(147) xor Codeword(177) xor
                Codeword(247) xor Codeword(314) xor Codeword(364) xor Codeword(415) xor
                Codeword(482) xor Codeword(521) xor Codeword(606) xor Codeword(623) xor
                Codeword(696) xor Codeword(803) xor Codeword(860) xor Codeword(933) xor
                Codeword(997) xor Codeword(1029) xor Codeword(1082) xor Codeword(1145) xor
                Codeword(1166) xor Codeword(1208) xor Codeword(1230) xor Codeword(1298) xor
                Codeword(1394) xor Codeword(1473) xor Codeword(1493) xor Codeword(1495) xor
                Codeword(1709) xor Codeword(1745) xor Codeword(1789) xor Codeword(1819);
 
     check57 <= Codeword(98) xor Codeword(146) xor Codeword(176) xor Codeword(246) xor
                Codeword(313) xor Codeword(363) xor Codeword(414) xor Codeword(481) xor
                Codeword(520) xor Codeword(605) xor Codeword(622) xor Codeword(695) xor
                Codeword(768) xor Codeword(802) xor Codeword(859) xor Codeword(932) xor
                Codeword(996) xor Codeword(1081) xor Codeword(1144) xor Codeword(1165) xor
                Codeword(1207) xor Codeword(1229) xor Codeword(1297) xor Codeword(1337) xor
                Codeword(1472) xor Codeword(1485) xor Codeword(1590) xor Codeword(1686) xor
                Codeword(1723) xor Codeword(1798) xor Codeword(1804) xor Codeword(1820);
 
     check58 <= Codeword(97) xor Codeword(145) xor Codeword(175) xor Codeword(312) xor
                Codeword(362) xor Codeword(413) xor Codeword(480) xor Codeword(519) xor
                Codeword(604) xor Codeword(621) xor Codeword(694) xor Codeword(767) xor
                Codeword(801) xor Codeword(858) xor Codeword(931) xor Codeword(995) xor
                Codeword(1028) xor Codeword(1080) xor Codeword(1143) xor Codeword(1164) xor
                Codeword(1206) xor Codeword(1228) xor Codeword(1336) xor Codeword(1393) xor
                Codeword(1471) xor Codeword(1589) xor Codeword(1685) xor Codeword(1838) xor
                Codeword(1851) xor Codeword(1870) xor Codeword(1928) xor Codeword(1929);
 
     check59 <= Codeword(144) xor Codeword(174) xor Codeword(245) xor Codeword(311) xor
                Codeword(361) xor Codeword(412) xor Codeword(479) xor Codeword(603) xor
                Codeword(693) xor Codeword(766) xor Codeword(857) xor Codeword(994) xor
                Codeword(1027) xor Codeword(1113) xor Codeword(1142) xor Codeword(1205) xor
                Codeword(1227) xor Codeword(1296) xor Codeword(1470) xor Codeword(1484) xor
                Codeword(1722) xor Codeword(1751) xor Codeword(1757) xor Codeword(1774) xor
                Codeword(1794) xor Codeword(1874) xor Codeword(1920) xor Codeword(1927) xor
                Codeword(1983) xor Codeword(2012) xor Codeword(2015) xor Codeword(2017);
 
     check60 <= Codeword(96) xor Codeword(143) xor Codeword(173) xor Codeword(244) xor
                Codeword(310) xor Codeword(360) xor Codeword(411) xor Codeword(478) xor
                Codeword(518) xor Codeword(692) xor Codeword(765) xor Codeword(800) xor
                Codeword(993) xor Codeword(1026) xor Codeword(1112) xor Codeword(1141) xor
                Codeword(1204) xor Codeword(1226) xor Codeword(1295) xor Codeword(1469) xor
                Codeword(1492) xor Codeword(1588) xor Codeword(1684) xor Codeword(1721) xor
                Codeword(1744) xor Codeword(1768) xor Codeword(1846) xor Codeword(1853) xor
                Codeword(1871) xor Codeword(1883) xor Codeword(1966) xor Codeword(1972);
 
     check61 <= Codeword(95) xor Codeword(142) xor Codeword(172) xor Codeword(243) xor
                Codeword(309) xor Codeword(359) xor Codeword(410) xor Codeword(477) xor
                Codeword(517) xor Codeword(602) xor Codeword(620) xor Codeword(691) xor
                Codeword(764) xor Codeword(856) xor Codeword(930) xor Codeword(992) xor
                Codeword(1025) xor Codeword(1079) xor Codeword(1110) xor Codeword(1140) xor
                Codeword(1203) xor Codeword(1225) xor Codeword(1294) xor Codeword(1335) xor
                Codeword(1392) xor Codeword(1468) xor Codeword(1491) xor Codeword(1683) xor
                Codeword(1719) xor Codeword(1799) xor Codeword(1805) xor Codeword(1821);
 
     check62 <= Codeword(94) xor Codeword(141) xor Codeword(171) xor Codeword(242) xor
                Codeword(308) xor Codeword(358) xor Codeword(409) xor Codeword(619) xor
                Codeword(690) xor Codeword(799) xor Codeword(855) xor Codeword(929) xor
                Codeword(1078) xor Codeword(1108) xor Codeword(1139) xor Codeword(1202) xor
                Codeword(1293) xor Codeword(1391) xor Codeword(1467) xor Codeword(1490) xor
                Codeword(1524) xor Codeword(1587) xor Codeword(1682) xor Codeword(1720) xor
                Codeword(1775) xor Codeword(1779) xor Codeword(1827) xor Codeword(1863) xor
                Codeword(1880) xor Codeword(2010) xor Codeword(2016) xor Codeword(2018);
 
     check63 <= Codeword(52) xor Codeword(93) xor Codeword(140) xor Codeword(357) xor
                Codeword(516) xor Codeword(601) xor Codeword(618) xor Codeword(763) xor
                Codeword(798) xor Codeword(928) xor Codeword(991) xor Codeword(1024) xor
                Codeword(1060) xor Codeword(1201) xor Codeword(1489) xor Codeword(1523) xor
                Codeword(1551) xor Codeword(1586) xor Codeword(1708) xor Codeword(1761) xor
                Codeword(1783) xor Codeword(1855) xor Codeword(1865) xor Codeword(1949) xor
                Codeword(1963) xor Codeword(1967) xor Codeword(1970) xor Codeword(1975) xor
                Codeword(2011) xor Codeword(2039) xor Codeword(2040) xor Codeword(2043);
 
     check64 <= Codeword(53) xor Codeword(109) xor Codeword(130) xor Codeword(245) xor
                Codeword(299) xor Codeword(342) xor Codeword(442) xor Codeword(458) xor
                Codeword(535) xor Codeword(580) xor Codeword(641) xor Codeword(763) xor
                Codeword(796) xor Codeword(859) xor Codeword(894) xor Codeword(944) xor
                Codeword(1038) xor Codeword(1074) xor Codeword(1158) xor Codeword(1171) xor
                Codeword(1245) xor Codeword(1287) xor Codeword(1346) xor Codeword(1416) xor
                Codeword(1574) xor Codeword(1582) xor Codeword(1664) xor Codeword(1740) xor
                Codeword(1902) xor Codeword(1960) xor Codeword(1992) xor Codeword(1994);
 
     check65 <= Codeword(51) xor Codeword(74) xor Codeword(141) xor Codeword(189) xor
                Codeword(286) xor Codeword(386) xor Codeword(399) xor Codeword(478) xor
                Codeword(521) xor Codeword(587) xor Codeword(655) xor Codeword(707) xor
                Codeword(757) xor Codeword(787) xor Codeword(943) xor Codeword(982) xor
                Codeword(1015) xor Codeword(1100) xor Codeword(1190) xor Codeword(1231) xor
                Codeword(1360) xor Codeword(1402) xor Codeword(1466) xor Codeword(1557) xor
                Codeword(1621) xor Codeword(1669) xor Codeword(1718) xor Codeword(1787) xor
                Codeword(1851) xor Codeword(1855) xor Codeword(1978) xor Codeword(1980);
 
     check66 <= Codeword(50) xor Codeword(66) xor Codeword(155) xor Codeword(244) xor
                Codeword(404) xor Codeword(480) xor Codeword(531) xor Codeword(609) xor
                Codeword(666) xor Codeword(701) xor Codeword(751) xor Codeword(871) xor
                Codeword(933) xor Codeword(973) xor Codeword(1045) xor Codeword(1065) xor
                Codeword(1144) xor Codeword(1174) xor Codeword(1265) xor Codeword(1322) xor
                Codeword(1391) xor Codeword(1606) xor Codeword(1675) xor Codeword(1705) xor
                Codeword(1854) xor Codeword(1860) xor Codeword(1875) xor Codeword(1930) xor
                Codeword(1940) xor Codeword(1995) xor Codeword(2011) xor Codeword(2019);
 
     check67 <= Codeword(97) xor Codeword(275) xor Codeword(322) xor Codeword(365) xor
                Codeword(393) xor Codeword(449) xor Codeword(524) xor Codeword(561) xor
                Codeword(638) xor Codeword(734) xor Codeword(874) xor Codeword(960) xor
                Codeword(1003) xor Codeword(1042) xor Codeword(1069) xor Codeword(1154) xor
                Codeword(1248) xor Codeword(1313) xor Codeword(1353) xor Codeword(1405) xor
                Codeword(1483) xor Codeword(1500) xor Codeword(1561) xor Codeword(1702) xor
                Codeword(1811) xor Codeword(1812) xor Codeword(1833) xor Codeword(1849) xor
                Codeword(1900) xor Codeword(1926) xor Codeword(2014) xor Codeword(2020);
 
     check68 <= Codeword(49) xor Codeword(112) xor Codeword(210) xor Codeword(256) xor
                Codeword(318) xor Codeword(381) xor Codeword(417) xor Codeword(485) xor
                Codeword(528) xor Codeword(601) xor Codeword(627) xor Codeword(694) xor
                Codeword(741) xor Codeword(791) xor Codeword(861) xor Codeword(897) xor
                Codeword(979) xor Codeword(1148) xor Codeword(1195) xor Codeword(1260) xor
                Codeword(1350) xor Codeword(1424) xor Codeword(1442) xor Codeword(1485) xor
                Codeword(1504) xor Codeword(1509) xor Codeword(1529) xor Codeword(1556) xor
                Codeword(1578) xor Codeword(1676) xor Codeword(1690) xor Codeword(1741);
 
     check69 <= Codeword(48) xor Codeword(101) xor Codeword(135) xor Codeword(215) xor
                Codeword(259) xor Codeword(283) xor Codeword(351) xor Codeword(498) xor
                Codeword(602) xor Codeword(674) xor Codeword(785) xor Codeword(836) xor
                Codeword(910) xor Codeword(951) xor Codeword(1051) xor Codeword(1152) xor
                Codeword(1272) xor Codeword(1282) xor Codeword(1364) xor Codeword(1517) xor
                Codeword(1540) xor Codeword(1563) xor Codeword(1607) xor Codeword(1759) xor
                Codeword(1773) xor Codeword(1779) xor Codeword(1839) xor Codeword(1948) xor
                Codeword(1951) xor Codeword(1982) xor Codeword(2015) xor Codeword(2021);
 
     check70 <= Codeword(47) xor Codeword(104) xor Codeword(136) xor Codeword(206) xor
                Codeword(246) xor Codeword(301) xor Codeword(389) xor Codeword(407) xor
                Codeword(450) xor Codeword(556) xor Codeword(572) xor Codeword(629) xor
                Codeword(713) xor Codeword(762) xor Codeword(822) xor Codeword(857) xor
                Codeword(921) xor Codeword(948) xor Codeword(1025) xor Codeword(1063) xor
                Codeword(1141) xor Codeword(1212) xor Codeword(1242) xor Codeword(1388) xor
                Codeword(1448) xor Codeword(1495) xor Codeword(1532) xor Codeword(1577) xor
                Codeword(1614) xor Codeword(1708) xor Codeword(1786) xor Codeword(1822);
 
     check71 <= Codeword(46) xor Codeword(95) xor Codeword(176) xor Codeword(276) xor
                Codeword(302) xor Codeword(353) xor Codeword(479) xor Codeword(538) xor
                Codeword(650) xor Codeword(739) xor Codeword(828) xor Codeword(883) xor
                Codeword(891) xor Codeword(964) xor Codeword(1034) xor Codeword(1121) xor
                Codeword(1198) xor Codeword(1233) xor Codeword(1284) xor Codeword(1431) xor
                Codeword(1452) xor Codeword(1481) xor Codeword(1541) xor Codeword(1651) xor
                Codeword(1707) xor Codeword(1813) xor Codeword(1847) xor Codeword(1937) xor
                Codeword(1952) xor Codeword(2018) xor Codeword(2030) xor Codeword(2039);
 
     check72 <= Codeword(45) xor Codeword(75) xor Codeword(162) xor Codeword(183) xor
                Codeword(243) xor Codeword(367) xor Codeword(435) xor Codeword(493) xor
                Codeword(552) xor Codeword(565) xor Codeword(657) xor Codeword(680) xor
                Codeword(775) xor Codeword(867) xor Codeword(935) xor Codeword(957) xor
                Codeword(1104) xor Codeword(1161) xor Codeword(1214) xor Codeword(1275) xor
                Codeword(1342) xor Codeword(1423) xor Codeword(1527) xor Codeword(1603) xor
                Codeword(1629) xor Codeword(1679) xor Codeword(1724) xor Codeword(1820) xor
                Codeword(1848) xor Codeword(1986) xor Codeword(2003) xor Codeword(2008);
 
     check73 <= Codeword(44) xor Codeword(56) xor Codeword(121) xor Codeword(219) xor
                Codeword(328) xor Codeword(363) xor Codeword(415) xor Codeword(507) xor
                Codeword(573) xor Codeword(708) xor Codeword(723) xor Codeword(795) xor
                Codeword(838) xor Codeword(923) xor Codeword(990) xor Codeword(1032) xor
                Codeword(1075) xor Codeword(1116) xor Codeword(1178) xor Codeword(1235) xor
                Codeword(1311) xor Codeword(1336) xor Codeword(1432) xor Codeword(1451) xor
                Codeword(1462) xor Codeword(1619) xor Codeword(1739) xor Codeword(1837) xor
                Codeword(1857) xor Codeword(1914) xor Codeword(1920) xor Codeword(1921);
 
     check74 <= Codeword(43) xor Codeword(70) xor Codeword(125) xor Codeword(221) xor
                Codeword(290) xor Codeword(384) xor Codeword(427) xor Codeword(501) xor
                Codeword(532) xor Codeword(658) xor Codeword(696) xor Codeword(764) xor
                Codeword(885) xor Codeword(938) xor Codeword(1023) xor Codeword(1073) xor
                Codeword(1127) xor Codeword(1187) xor Codeword(1254) xor Codeword(1318) xor
                Codeword(1339) xor Codeword(1387) xor Codeword(1397) xor Codeword(1446) xor
                Codeword(1583) xor Codeword(1634) xor Codeword(1658) xor Codeword(1758) xor
                Codeword(1791) xor Codeword(1796) xor Codeword(1836) xor Codeword(1880);
 
     check75 <= Codeword(42) xor Codeword(81) xor Codeword(170) xor Codeword(192) xor
                Codeword(278) xor Codeword(294) xor Codeword(347) xor Codeword(436) xor
                Codeword(468) xor Codeword(520) xor Codeword(615) xor Codeword(649) xor
                Codeword(682) xor Codeword(740) xor Codeword(807) xor Codeword(872) xor
                Codeword(903) xor Codeword(993) xor Codeword(1004) xor Codeword(1102) xor
                Codeword(1155) xor Codeword(1183) xor Codeword(1262) xor Codeword(1279) xor
                Codeword(1288) xor Codeword(1468) xor Codeword(1534) xor Codeword(1545) xor
                Codeword(1581) xor Codeword(1685) xor Codeword(1775) xor Codeword(1823);
 
     check76 <= Codeword(41) xor Codeword(106) xor Codeword(124) xor Codeword(174) xor
                Codeword(270) xor Codeword(332) xor Codeword(348) xor Codeword(408) xor
                Codeword(481) xor Codeword(509) xor Codeword(588) xor Codeword(619) xor
                Codeword(699) xor Codeword(761) xor Codeword(810) xor Codeword(835) xor
                Codeword(912) xor Codeword(997) xor Codeword(1041) xor Codeword(1086) xor
                Codeword(1143) xor Codeword(1188) xor Codeword(1257) xor Codeword(1286) xor
                Codeword(1365) xor Codeword(1460) xor Codeword(1475) xor Codeword(1547) xor
                Codeword(1609) xor Codeword(1653) xor Codeword(1694) xor Codeword(1742);
 
     check77 <= Codeword(119) xor Codeword(185) xor Codeword(257) xor Codeword(293) xor
                Codeword(383) xor Codeword(423) xor Codeword(477) xor Codeword(523) xor
                Codeword(568) xor Codeword(624) xor Codeword(717) xor Codeword(722) xor
                Codeword(731) xor Codeword(797) xor Codeword(865) xor Codeword(908) xor
                Codeword(987) xor Codeword(1055) xor Codeword(1088) xor Codeword(1177) xor
                Codeword(1263) xor Codeword(1316) xor Codeword(1349) xor Codeword(1409) xor
                Codeword(1435) xor Codeword(1624) xor Codeword(1659) xor Codeword(1810) xor
                Codeword(1845) xor Codeword(2013) xor Codeword(2017) xor Codeword(2031);
 
     check78 <= Codeword(40) xor Codeword(84) xor Codeword(159) xor Codeword(193) xor
                Codeword(274) xor Codeword(288) xor Codeword(374) xor Codeword(391) xor
                Codeword(395) xor Codeword(496) xor Codeword(544) xor Codeword(590) xor
                Codeword(662) xor Codeword(672) xor Codeword(772) xor Codeword(827) xor
                Codeword(863) xor Codeword(913) xor Codeword(965) xor Codeword(1009) xor
                Codeword(1076) xor Codeword(1146) xor Codeword(1200) xor Codeword(1253) xor
                Codeword(1300) xor Codeword(1361) xor Codeword(1392) xor Codeword(1437) xor
                Codeword(1593) xor Codeword(1616) xor Codeword(1680) xor Codeword(1743);
 
     check79 <= Codeword(39) xor Codeword(99) xor Codeword(167) xor Codeword(220) xor
                Codeword(325) xor Codeword(430) xor Codeword(463) xor Codeword(721) xor
                Codeword(742) xor Codeword(794) xor Codeword(902) xor Codeword(947) xor
                Codeword(1035) xor Codeword(1103) xor Codeword(1207) xor Codeword(1331) xor
                Codeword(1371) xor Codeword(1401) xor Codeword(1512) xor Codeword(1521) xor
                Codeword(1567) xor Codeword(1727) xor Codeword(1769) xor Codeword(1776) xor
                Codeword(1777) xor Codeword(1801) xor Codeword(1866) xor Codeword(1883) xor
                Codeword(1891) xor Codeword(1950) xor Codeword(2026) xor Codeword(2032);
 
     check80 <= Codeword(38) xor Codeword(62) xor Codeword(131) xor Codeword(182) xor
                Codeword(248) xor Codeword(337) xor Codeword(397) xor Codeword(549) xor
                Codeword(600) xor Codeword(632) xor Codeword(673) xor Codeword(733) xor
                Codeword(869) xor Codeword(926) xor Codeword(961) xor Codeword(1072) xor
                Codeword(1118) xor Codeword(1166) xor Codeword(1192) xor Codeword(1228) xor
                Codeword(1289) xor Codeword(1343) xor Codeword(1410) xor Codeword(1461) xor
                Codeword(1484) xor Codeword(1695) xor Codeword(1730) xor Codeword(1915) xor
                Codeword(1961) xor Codeword(1967) xor Codeword(2010) xor Codeword(2022);
 
     check81 <= Codeword(37) xor Codeword(72) xor Codeword(129) xor Codeword(262) xor
                Codeword(409) xor Codeword(495) xor Codeword(554) xor Codeword(563) xor
                Codeword(617) xor Codeword(804) xor Codeword(846) xor Codeword(972) xor
                Codeword(1012) xor Codeword(1095) xor Codeword(1114) xor Codeword(1168) xor
                Codeword(1267) xor Codeword(1317) xor Codeword(1496) xor Codeword(1546) xor
                Codeword(1560) xor Codeword(1580) xor Codeword(1647) xor Codeword(1655) xor
                Codeword(1867) xor Codeword(1874) xor Codeword(1878) xor Codeword(1949) xor
                Codeword(1956) xor Codeword(1957) xor Codeword(1971) xor Codeword(1973);
 
     check82 <= Codeword(36) xor Codeword(67) xor Codeword(165) xor Codeword(188) xor
                Codeword(254) xor Codeword(298) xor Codeword(336) xor Codeword(486) xor
                Codeword(543) xor Codeword(584) xor Codeword(626) xor Codeword(685) xor
                Codeword(738) xor Codeword(777) xor Codeword(829) xor Codeword(856) xor
                Codeword(916) xor Codeword(1000) xor Codeword(1027) xor Codeword(1082) xor
                Codeword(1119) xor Codeword(1216) xor Codeword(1269) xor Codeword(1374) xor
                Codeword(1396) xor Codeword(1490) xor Codeword(1568) xor Codeword(1601) xor
                Codeword(1670) xor Codeword(1763) xor Codeword(1788) xor Codeword(1824);
 
     check83 <= Codeword(35) xor Codeword(73) xor Codeword(144) xor Codeword(208) xor
                Codeword(232) xor Codeword(330) xor Codeword(425) xor Codeword(448) xor
                Codeword(511) xor Codeword(585) xor Codeword(633) xor Codeword(691) xor
                Codeword(821) xor Codeword(850) xor Codeword(918) xor Codeword(989) xor
                Codeword(1047) xor Codeword(1105) xor Codeword(1239) xor Codeword(1309) xor
                Codeword(1332) xor Codeword(1425) xor Codeword(1436) xor Codeword(1511) xor
                Codeword(1590) xor Codeword(1641) xor Codeword(1681) xor Codeword(1693) xor
                Codeword(1819) xor Codeword(1871) xor Codeword(1919) xor Codeword(1922);
 
     check84 <= Codeword(34) xor Codeword(61) xor Codeword(147) xor Codeword(222) xor
                Codeword(310) xor Codeword(371) xor Codeword(392) xor Codeword(453) xor
                Codeword(562) xor Codeword(663) xor Codeword(676) xor Codeword(766) xor
                Codeword(808) xor Codeword(854) xor Codeword(942) xor Codeword(975) xor
                Codeword(1057) xor Codeword(1097) xor Codeword(1132) xor Codeword(1211) xor
                Codeword(1404) xor Codeword(1455) xor Codeword(1463) xor Codeword(1474) xor
                Codeword(1625) xor Codeword(1678) xor Codeword(1761) xor Codeword(1804) xor
                Codeword(1863) xor Codeword(1870) xor Codeword(1897) xor Codeword(1907);
 
     check85 <= Codeword(33) xor Codeword(132) xor Codeword(218) xor Codeword(235) xor
                Codeword(313) xor Codeword(379) xor Codeword(505) xor Codeword(558) xor
                Codeword(608) xor Codeword(623) xor Codeword(677) xor Codeword(725) xor
                Codeword(843) xor Codeword(924) xor Codeword(1052) xor Codeword(1087) xor
                Codeword(1217) xor Codeword(1232) xor Codeword(1277) xor Codeword(1319) xor
                Codeword(1363) xor Codeword(1389) xor Codeword(1652) xor Codeword(1768) xor
                Codeword(1770) xor Codeword(1772) xor Codeword(1815) xor Codeword(1872) xor
                Codeword(1909) xor Codeword(2016) xor Codeword(2038) xor Codeword(2043);
 
     check86 <= Codeword(32) xor Codeword(166) xor Codeword(239) xor Codeword(343) xor
                Codeword(424) xor Codeword(452) xor Codeword(559) xor Codeword(571) xor
                Codeword(651) xor Codeword(703) xor Codeword(773) xor Codeword(877) xor
                Codeword(934) xor Codeword(953) xor Codeword(1058) xor Codeword(1101) xor
                Codeword(1112) xor Codeword(1122) xor Codeword(1310) xor Codeword(1358) xor
                Codeword(1620) xor Codeword(1756) xor Codeword(1762) xor Codeword(1802) xor
                Codeword(1916) xor Codeword(1944) xor Codeword(1946) xor Codeword(1954) xor
                Codeword(1983) xor Codeword(1993) xor Codeword(1996) xor Codeword(2001);
 
     check87 <= Codeword(31) xor Codeword(77) xor Codeword(128) xor Codeword(203) xor
                Codeword(229) xor Codeword(331) xor Codeword(341) xor Codeword(416) xor
                Codeword(503) xor Codeword(526) xor Codeword(576) xor Codeword(683) xor
                Codeword(799) xor Codeword(862) xor Codeword(963) xor Codeword(1046) xor
                Codeword(1124) xor Codeword(1206) xor Codeword(1268) xor Codeword(1426) xor
                Codeword(1459) xor Codeword(1544) xor Codeword(1554) xor Codeword(1731) xor
                Codeword(1765) xor Codeword(1832) xor Codeword(1842) xor Codeword(1853) xor
                Codeword(1869) xor Codeword(1917) xor Codeword(2000) xor Codeword(2005);
 
     check88 <= Codeword(30) xor Codeword(79) xor Codeword(156) xor Codeword(204) xor
                Codeword(263) xor Codeword(297) xor Codeword(377) xor Codeword(434) xor
                Codeword(484) xor Codeword(616) xor Codeword(695) xor Codeword(759) xor
                Codeword(813) xor Codeword(873) xor Codeword(917) xor Codeword(958) xor
                Codeword(1014) xor Codeword(1150) xor Codeword(1179) xor Codeword(1227) xor
                Codeword(1278) xor Codeword(1315) xor Codeword(1354) xor Codeword(1399) xor
                Codeword(1438) xor Codeword(1700) xor Codeword(1799) xor Codeword(1903) xor
                Codeword(1911) xor Codeword(1929) xor Codeword(2037) xor Codeword(2040);
 
     check89 <= Codeword(29) xor Codeword(102) xor Codeword(140) xor Codeword(184) xor
                Codeword(247) xor Codeword(355) xor Codeword(438) xor Codeword(491) xor
                Codeword(519) xor Codeword(575) xor Codeword(664) xor Codeword(704) xor
                Codeword(752) xor Codeword(884) xor Codeword(1130) xor Codeword(1167) xor
                Codeword(1213) xor Codeword(1293) xor Codeword(1377) xor Codeword(1421) xor
                Codeword(1585) xor Codeword(1643) xor Codeword(1686) xor Codeword(1725) xor
                Codeword(1861) xor Codeword(1892) xor Codeword(1894) xor Codeword(1918) xor
                Codeword(1935) xor Codeword(1972) xor Codeword(2025) xor Codeword(2033);
 
     check90 <= Codeword(28) xor Codeword(85) xor Codeword(168) xor Codeword(175) xor
                Codeword(258) xor Codeword(307) xor Codeword(358) xor Codeword(447) xor
                Codeword(459) xor Codeword(527) xor Codeword(661) xor Codeword(756) xor
                Codeword(783) xor Codeword(904) xor Codeword(952) xor Codeword(1084) xor
                Codeword(1142) xor Codeword(1181) xor Codeword(1291) xor Codeword(1330) xor
                Codeword(1383) xor Codeword(1559) xor Codeword(1630) xor Codeword(1703) xor
                Codeword(1834) xor Codeword(1841) xor Codeword(1846) xor Codeword(1881) xor
                Codeword(1882) xor Codeword(1888) xor Codeword(1923) xor Codeword(1925);
 
     check91 <= Codeword(27) xor Codeword(96) xor Codeword(158) xor Codeword(191) xor
                Codeword(269) xor Codeword(280) xor Codeword(344) xor Codeword(457) xor
                Codeword(606) xor Codeword(690) xor Codeword(746) xor Codeword(792) xor
                Codeword(845) xor Codeword(937) xor Codeword(978) xor Codeword(1007) xor
                Codeword(1059) xor Codeword(1151) xor Codeword(1193) xor Codeword(1256) xor
                Codeword(1367) xor Codeword(1384) xor Codeword(1398) xor Codeword(1591) xor
                Codeword(1645) xor Codeword(1733) xor Codeword(1792) xor Codeword(1905) xor
                Codeword(1979) xor Codeword(1999) xor Codeword(2028) xor Codeword(2034);
 
     check92 <= Codeword(26) xor Codeword(103) xor Codeword(145) xor Codeword(195) xor
                Codeword(242) xor Codeword(324) xor Codeword(378) xor Codeword(432) xor
                Codeword(489) xor Codeword(516) xor Codeword(613) xor Codeword(646) xor
                Codeword(718) xor Codeword(726) xor Codeword(786) xor Codeword(831) xor
                Codeword(887) xor Codeword(906) xor Codeword(984) xor Codeword(1030) xor
                Codeword(1070) xor Codeword(1123) xor Codeword(1191) xor Codeword(1270) xor
                Codeword(1298) xor Codeword(1369) xor Codeword(1385) xor Codeword(1478) xor
                Codeword(1613) xor Codeword(1687) xor Codeword(1697) xor Codeword(1744);
 
     check93 <= Codeword(25) xor Codeword(78) xor Codeword(164) xor Codeword(224) xor
                Codeword(231) xor Codeword(311) xor Codeword(340) xor Codeword(413) xor
                Codeword(471) xor Codeword(545) xor Codeword(581) xor Codeword(647) xor
                Codeword(698) xor Codeword(765) xor Codeword(790) xor Codeword(848) xor
                Codeword(919) xor Codeword(967) xor Codeword(1013) xor Codeword(1064) xor
                Codeword(1138) xor Codeword(1209) xor Codeword(1219) xor Codeword(1266) xor
                Codeword(1327) xor Codeword(1408) xor Codeword(1456) xor Codeword(1579) xor
                Codeword(1622) xor Codeword(1661) xor Codeword(1715) xor Codeword(1745);
 
     check94 <= Codeword(24) xor Codeword(92) xor Codeword(194) xor Codeword(329) xor
                Codeword(368) xor Codeword(421) xor Codeword(474) xor Codeword(522) xor
                Codeword(579) xor Codeword(719) xor Codeword(776) xor Codeword(780) xor
                Codeword(915) xor Codeword(969) xor Codeword(1024) xor Codeword(1068) xor
                Codeword(1164) xor Codeword(1175) xor Codeword(1230) xor Codeword(1375) xor
                Codeword(1412) xor Codeword(1467) xor Codeword(1482) xor Codeword(1617) xor
                Codeword(1656) xor Codeword(1805) xor Codeword(1887) xor Codeword(1895) xor
                Codeword(1901) xor Codeword(1933) xor Codeword(1936) xor Codeword(1943);
 
     check95 <= Codeword(23) xor Codeword(63) xor Codeword(134) xor Codeword(190) xor
                Codeword(234) xor Codeword(303) xor Codeword(352) xor Codeword(443) xor
                Codeword(460) xor Codeword(547) xor Codeword(611) xor Codeword(618) xor
                Codeword(678) xor Codeword(732) xor Codeword(814) xor Codeword(875) xor
                Codeword(932) xor Codeword(995) xor Codeword(1031) xor Codeword(1145) xor
                Codeword(1176) xor Codeword(1250) xor Codeword(1444) xor Codeword(1487) xor
                Codeword(1507) xor Codeword(1528) xor Codeword(1535) xor Codeword(1552) xor
                Codeword(1566) xor Codeword(1623) xor Codeword(1684) xor Codeword(1746);
 
     check96 <= Codeword(22) xor Codeword(98) xor Codeword(150) xor Codeword(172) xor
                Codeword(251) xor Codeword(380) xor Codeword(441) xor Codeword(490) xor
                Codeword(560) xor Codeword(592) xor Codeword(631) xor Codeword(675) xor
                Codeword(760) xor Codeword(798) xor Codeword(870) xor Codeword(899) xor
                Codeword(976) xor Codeword(1006) xor Codeword(1090) xor Codeword(1208) xor
                Codeword(1251) xor Codeword(1283) xor Codeword(1338) xor Codeword(1453) xor
                Codeword(1476) xor Codeword(1513) xor Codeword(1571) xor Codeword(1612) xor
                Codeword(1689) xor Codeword(1735) xor Codeword(1886) xor Codeword(1908);
 
     check97 <= Codeword(21) xor Codeword(65) xor Codeword(142) xor Codeword(180) xor
                Codeword(260) xor Codeword(316) xor Codeword(370) xor Codeword(419) xor
                Codeword(456) xor Codeword(557) xor Codeword(595) xor Codeword(636) xor
                Codeword(693) xor Codeword(748) xor Codeword(809) xor Codeword(876) xor
                Codeword(900) xor Codeword(988) xor Codeword(1020) xor Codeword(1077) xor
                Codeword(1125) xor Codeword(1199) xor Codeword(1229) xor Codeword(1324) xor
                Codeword(1368) xor Codeword(1406) xor Codeword(1447) xor Codeword(1575) xor
                Codeword(1596) xor Codeword(1633) xor Codeword(1665) xor Codeword(1747);
 
     check98 <= Codeword(20) xor Codeword(116) xor Codeword(199) xor Codeword(255) xor
                Codeword(308) xor Codeword(356) xor Codeword(400) xor Codeword(482) xor
                Codeword(518) xor Codeword(582) xor Codeword(668) xor Codeword(714) xor
                Codeword(735) xor Codeword(820) xor Codeword(866) xor Codeword(931) xor
                Codeword(996) xor Codeword(1048) xor Codeword(1215) xor Codeword(1382) xor
                Codeword(1450) xor Codeword(1520) xor Codeword(1551) xor Codeword(1570) xor
                Codeword(1584) xor Codeword(1638) xor Codeword(1699) xor Codeword(1781) xor
                Codeword(1818) xor Codeword(1968) xor Codeword(2036) xor Codeword(2041);
 
     check99 <= Codeword(19) xor Codeword(76) xor Codeword(126) xor Codeword(198) xor
                Codeword(261) xor Codeword(285) xor Codeword(376) xor Codeword(402) xor
                Codeword(467) xor Codeword(540) xor Codeword(612) xor Codeword(635) xor
                Codeword(715) xor Codeword(750) xor Codeword(793) xor Codeword(834) xor
                Codeword(925) xor Codeword(968) xor Codeword(1026) xor Codeword(1096) xor
                Codeword(1140) xor Codeword(1238) xor Codeword(1290) xor Codeword(1355) xor
                Codeword(1395) xor Codeword(1558) xor Codeword(1564) xor Codeword(1592) xor
                Codeword(1626) xor Codeword(1649) xor Codeword(1691) xor Codeword(1748);
 
     check100 <= Codeword(18) xor Codeword(94) xor Codeword(120) xor Codeword(178) xor
                Codeword(250) xor Codeword(295) xor Codeword(349) xor Codeword(444) xor
                Codeword(492) xor Codeword(541) xor Codeword(578) xor Codeword(692) xor
                Codeword(770) xor Codeword(782) xor Codeword(840) xor Codeword(941) xor
                Codeword(983) xor Codeword(1050) xor Codeword(1071) xor Codeword(1163) xor
                Codeword(1220) xor Codeword(1241) xor Codeword(1301) xor Codeword(1335) xor
                Codeword(1417) xor Codeword(1441) xor Codeword(1519) xor Codeword(1602) xor
                Codeword(1627) xor Codeword(1671) xor Codeword(1778) xor Codeword(1825);
 
     check101 <= Codeword(17) xor Codeword(58) xor Codeword(123) xor Codeword(211) xor
                Codeword(273) xor Codeword(289) xor Codeword(346) xor Codeword(420) xor
                Codeword(517) xor Codeword(603) xor Codeword(684) xor Codeword(724) xor
                Codeword(823) xor Codeword(830) xor Codeword(879) xor Codeword(889) xor
                Codeword(954) xor Codeword(1357) xor Codeword(1472) xor Codeword(1488) xor
                Codeword(1508) xor Codeword(1516) xor Codeword(1525) xor Codeword(1674) xor
                Codeword(1710) xor Codeword(1831) xor Codeword(1840) xor Codeword(1850) xor
                Codeword(1884) xor Codeword(1912) xor Codeword(1997) xor Codeword(2002);
 
     check102 <= Codeword(16) xor Codeword(59) xor Codeword(113) xor Codeword(214) xor
                Codeword(226) xor Codeword(361) xor Codeword(440) xor Codeword(472) xor
                Codeword(510) xor Codeword(589) xor Codeword(621) xor Codeword(702) xor
                Codeword(774) xor Codeword(881) xor Codeword(991) xor Codeword(1005) xor
                Codeword(1098) xor Codeword(1139) xor Codeword(1285) xor Codeword(1477) xor
                Codeword(1502) xor Codeword(1631) xor Codeword(1666) xor Codeword(1713) xor
                Codeword(1798) xor Codeword(1844) xor Codeword(1890) xor Codeword(1906) xor
                Codeword(1989) xor Codeword(2004) xor Codeword(2023) xor Codeword(2027);
 
     check103 <= Codeword(15) xor Codeword(93) xor Codeword(151) xor Codeword(200) xor
                Codeword(265) xor Codeword(284) xor Codeword(354) xor Codeword(410) xor
                Codeword(488) xor Codeword(525) xor Codeword(614) xor Codeword(642) xor
                Codeword(706) xor Codeword(802) xor Codeword(852) xor Codeword(888) xor
                Codeword(956) xor Codeword(1022) xor Codeword(1062) xor Codeword(1131) xor
                Codeword(1197) xor Codeword(1236) xor Codeword(1326) xor Codeword(1366) xor
                Codeword(1538) xor Codeword(1553) xor Codeword(1573) xor Codeword(1604) xor
                Codeword(1642) xor Codeword(1650) xor Codeword(1712) xor Codeword(1749);
 
     check104 <= Codeword(14) xor Codeword(86) xor Codeword(133) xor Codeword(179) xor
                Codeword(267) xor Codeword(317) xor Codeword(388) xor Codeword(396) xor
                Codeword(464) xor Codeword(530) xor Codeword(605) xor Codeword(640) xor
                Codeword(769) xor Codeword(811) xor Codeword(832) xor Codeword(939) xor
                Codeword(970) xor Codeword(1043) xor Codeword(1080) xor Codeword(1149) xor
                Codeword(1204) xor Codeword(1274) xor Codeword(1312) xor Codeword(1454) xor
                Codeword(1470) xor Codeword(1480) xor Codeword(1489) xor Codeword(1498) xor
                Codeword(1533) xor Codeword(1663) xor Codeword(1714) xor Codeword(1750);
 
     check105 <= Codeword(13) xor Codeword(146) xor Codeword(197) xor Codeword(237) xor
                Codeword(300) xor Codeword(338) xor Codeword(422) xor Codeword(462) xor
                Codeword(593) xor Codeword(705) xor Codeword(737) xor Codeword(806) xor
                Codeword(844) xor Codeword(922) xor Codeword(966) xor Codeword(1044) xor
                Codeword(1089) xor Codeword(1172) xor Codeword(1225) xor Codeword(1351) xor
                Codeword(1418) xor Codeword(1428) xor Codeword(1443) xor Codeword(1497) xor
                Codeword(1526) xor Codeword(1709) xor Codeword(1783) xor Codeword(1806) xor
                Codeword(1966) xor Codeword(2012) xor Codeword(2044) xor Codeword(2046);
 
     check106 <= Codeword(12) xor Codeword(157) xor Codeword(223) xor Codeword(272) xor
                Codeword(312) xor Codeword(333) xor Codeword(412) xor Codeword(529) xor
                Codeword(610) xor Codeword(700) xor Codeword(744) xor Codeword(812) xor
                Codeword(853) xor Codeword(929) xor Codeword(986) xor Codeword(1021) xor
                Codeword(1085) xor Codeword(1170) xor Codeword(1246) xor Codeword(1280) xor
                Codeword(1295) xor Codeword(1352) xor Codeword(1394) xor Codeword(1514) xor
                Codeword(1594) xor Codeword(1637) xor Codeword(1803) xor Codeword(1807) xor
                Codeword(1885) xor Codeword(1938) xor Codeword(1953) xor Codeword(1963);
 
     check107 <= Codeword(110) xor Codeword(127) xor Codeword(207) xor Codeword(230) xor
                Codeword(323) xor Codeword(335) xor Codeword(469) xor Codeword(586) xor
                Codeword(656) xor Codeword(681) xor Codeword(728) xor Codeword(801) xor
                Codeword(880) xor Codeword(895) xor Codeword(949) xor Codeword(1153) xor
                Codeword(1202) xor Codeword(1244) xor Codeword(1302) xor Codeword(1333) xor
                Codeword(1415) xor Codeword(1445) xor Codeword(1729) xor Codeword(1793) xor
                Codeword(1797) xor Codeword(1817) xor Codeword(1835) xor Codeword(1889) xor
                Codeword(1977) xor Codeword(1981) xor Codeword(2045) xor Codeword(2047);
 
     check108 <= Codeword(11) xor Codeword(105) xor Codeword(115) xor Codeword(181) xor
                Codeword(238) xor Codeword(296) xor Codeword(385) xor Codeword(418) xor
                Codeword(500) xor Codeword(508) xor Codeword(583) xor Codeword(643) xor
                Codeword(689) xor Codeword(730) xor Codeword(826) xor Codeword(839) xor
                Codeword(893) xor Codeword(950) xor Codeword(1029) xor Codeword(1108) xor
                Codeword(1147) xor Codeword(1184) xor Codeword(1299) xor Codeword(1376) xor
                Codeword(1471) xor Codeword(1523) xor Codeword(1548) xor Codeword(1595) xor
                Codeword(1644) xor Codeword(1683) xor Codeword(1717) xor Codeword(1751);
 
     check109 <= Codeword(10) xor Codeword(100) xor Codeword(160) xor Codeword(171) xor
                Codeword(266) xor Codeword(362) xor Codeword(454) xor Codeword(598) xor
                Codeword(711) xor Codeword(754) xor Codeword(778) xor Codeword(927) xor
                Codeword(985) xor Codeword(1129) xor Codeword(1169) xor Codeword(1186) xor
                Codeword(1258) xor Codeword(1303) xor Codeword(1337) xor Codeword(1588) xor
                Codeword(1615) xor Codeword(1672) xor Codeword(1732) xor Codeword(1734) xor
                Codeword(1767) xor Codeword(1858) xor Codeword(1893) xor Codeword(1927) xor
                Codeword(1939) xor Codeword(2007) xor Codeword(2029) xor Codeword(2042);
 
     check110 <= Codeword(9) xor Codeword(83) xor Codeword(118) xor Codeword(212) xor
                Codeword(225) xor Codeword(326) xor Codeword(345) xor Codeword(446) xor
                Codeword(504) xor Codeword(536) xor Codeword(591) xor Codeword(639) xor
                Codeword(710) xor Codeword(736) xor Codeword(816) xor Codeword(847) xor
                Codeword(909) xor Codeword(977) xor Codeword(1107) xor Codeword(1136) xor
                Codeword(1165) xor Codeword(1173) xor Codeword(1261) xor Codeword(1294) xor
                Codeword(1341) xor Codeword(1439) xor Codeword(1458) xor Codeword(1494) xor
                Codeword(1505) xor Codeword(1628) xor Codeword(1704) xor Codeword(1752);
 
     check111 <= Codeword(8) xor Codeword(90) xor Codeword(138) xor Codeword(177) xor
                Codeword(252) xor Codeword(287) xor Codeword(357) xor Codeword(405) xor
                Codeword(451) xor Codeword(534) xor Codeword(567) xor Codeword(665) xor
                Codeword(687) xor Codeword(747) xor Codeword(818) xor Codeword(868) xor
                Codeword(911) xor Codeword(994) xor Codeword(1033) xor Codeword(1092) xor
                Codeword(1159) xor Codeword(1203) xor Codeword(1218) xor Codeword(1247) xor
                Codeword(1314) xor Codeword(1390) xor Codeword(1465) xor Codeword(1536) xor
                Codeword(1550) xor Codeword(1668) xor Codeword(1782) xor Codeword(1826);
 
     check112 <= Codeword(7) xor Codeword(54) xor Codeword(148) xor Codeword(205) xor
                Codeword(233) xor Codeword(305) xor Codeword(369) xor Codeword(398) xor
                Codeword(497) xor Codeword(513) xor Codeword(577) xor Codeword(652) xor
                Codeword(669) xor Codeword(755) xor Codeword(788) xor Codeword(882) xor
                Codeword(896) xor Codeword(999) xor Codeword(1028) xor Codeword(1060) xor
                Codeword(1094) xor Codeword(1157) xor Codeword(1321) xor Codeword(1340) xor
                Codeword(1473) xor Codeword(1518) xor Codeword(1524) xor Codeword(1598) xor
                Codeword(1640) xor Codeword(1667) xor Codeword(1698) xor Codeword(1753);
 
     check113 <= Codeword(6) xor Codeword(108) xor Codeword(143) xor Codeword(202) xor
                Codeword(253) xor Codeword(314) xor Codeword(339) xor Codeword(429) xor
                Codeword(550) xor Codeword(570) xor Codeword(622) xor Codeword(671) xor
                Codeword(729) xor Codeword(824) xor Codeword(878) xor Codeword(928) xor
                Codeword(1011) xor Codeword(1066) xor Codeword(1134) xor Codeword(1194) xor
                Codeword(1243) xor Codeword(1305) xor Codeword(1329) xor Codeword(1393) xor
                Codeword(1440) xor Codeword(1503) xor Codeword(1610) xor Codeword(1677) xor
                Codeword(1728) xor Codeword(1737) xor Codeword(1794) xor Codeword(1827);
 
     check114 <= Codeword(5) xor Codeword(88) xor Codeword(149) xor Codeword(216) xor
                Codeword(268) xor Codeword(309) xor Codeword(387) xor Codeword(439) xor
                Codeword(461) xor Codeword(553) xor Codeword(574) xor Codeword(667) xor
                Codeword(712) xor Codeword(743) xor Codeword(781) xor Codeword(842) xor
                Codeword(892) xor Codeword(998) xor Codeword(1018) xor Codeword(1099) xor
                Codeword(1180) xor Codeword(1271) xor Codeword(1307) xor Codeword(1373) xor
                Codeword(1422) xor Codeword(1429) xor Codeword(1486) xor Codeword(1555) xor
                Codeword(1611) xor Codeword(1736) xor Codeword(1809) xor Codeword(1828);
 
     check115 <= Codeword(4) xor Codeword(68) xor Codeword(137) xor Codeword(209) xor
                Codeword(264) xor Codeword(315) xor Codeword(372) xor Codeword(433) xor
                Codeword(473) xor Codeword(537) xor Codeword(564) xor Codeword(654) xor
                Codeword(688) xor Codeword(771) xor Codeword(789) xor Codeword(864) xor
                Codeword(920) xor Codeword(992) xor Codeword(1039) xor Codeword(1111) xor
                Codeword(1117) xor Codeword(1205) xor Codeword(1222) xor Codeword(1255) xor
                Codeword(1380) xor Codeword(1420) xor Codeword(1469) xor Codeword(1530) xor
                Codeword(1605) xor Codeword(1639) xor Codeword(1654) xor Codeword(1754);
 
     check116 <= Codeword(71) xor Codeword(163) xor Codeword(187) xor Codeword(228) xor
                Codeword(304) xor Codeword(390) xor Codeword(437) xor Codeword(483) xor
                Codeword(514) xor Codeword(599) xor Codeword(620) xor Codeword(709) xor
                Codeword(749) xor Codeword(817) xor Codeword(905) xor Codeword(974) xor
                Codeword(1037) xor Codeword(1067) xor Codeword(1160) xor Codeword(1196) xor
                Codeword(1224) xor Codeword(1226) xor Codeword(1347) xor Codeword(1386) xor
                Codeword(1542) xor Codeword(1632) xor Codeword(1662) xor Codeword(1785) xor
                Codeword(1947) xor Codeword(1998) xor Codeword(2024) xor Codeword(2035);
 
     check117 <= Codeword(3) xor Codeword(55) xor Codeword(111) xor Codeword(196) xor
                Codeword(426) xor Codeword(455) xor Codeword(533) xor Codeword(648) xor
                Codeword(679) xor Codeword(841) xor Codeword(930) xor Codeword(981) xor
                Codeword(1016) xor Codeword(1093) xor Codeword(1135) xor Codeword(1185) xor
                Codeword(1273) xor Codeword(1325) xor Codeword(1345) xor Codeword(1449) xor
                Codeword(1537) xor Codeword(1576) xor Codeword(1657) xor Codeword(1701) xor
                Codeword(1808) xor Codeword(1864) xor Codeword(1877) xor Codeword(1913) xor
                Codeword(1931) xor Codeword(1934) xor Codeword(1965) xor Codeword(1974);
 
     check118 <= Codeword(2) xor Codeword(89) xor Codeword(152) xor Codeword(249) xor
                Codeword(282) xor Codeword(359) xor Codeword(406) xor Codeword(499) xor
                Codeword(506) xor Codeword(594) xor Codeword(645) xor Codeword(803) xor
                Codeword(833) xor Codeword(945) xor Codeword(1053) xor Codeword(1106) xor
                Codeword(1156) xor Codeword(1201) xor Codeword(1259) xor Codeword(1281) xor
                Codeword(1378) xor Codeword(1403) xor Codeword(1433) xor Codeword(1492) xor
                Codeword(1531) xor Codeword(1599) xor Codeword(1660) xor Codeword(1711) xor
                Codeword(1873) xor Codeword(1924) xor Codeword(1984) xor Codeword(1985);
 
     check119 <= Codeword(1) xor Codeword(107) xor Codeword(154) xor Codeword(227) xor
                Codeword(319) xor Codeword(445) xor Codeword(546) xor Codeword(604) xor
                Codeword(659) xor Codeword(727) xor Codeword(784) xor Codeword(851) xor
                Codeword(1002) xor Codeword(1056) xor Codeword(1081) xor Codeword(1126) xor
                Codeword(1306) xor Codeword(1359) xor Codeword(1413) xor Codeword(1427) xor
                Codeword(1464) xor Codeword(1522) xor Codeword(1648) xor Codeword(1688) xor
                Codeword(1800) xor Codeword(1879) xor Codeword(1941) xor Codeword(1942) xor
                Codeword(1945) xor Codeword(1955) xor Codeword(1969) xor Codeword(1975);
 
     check120 <= Codeword(0) xor Codeword(80) xor Codeword(321) xor Codeword(360) xor
                Codeword(401) xor Codeword(502) xor Codeword(515) xor Codeword(653) xor
                Codeword(745) xor Codeword(805) xor Codeword(855) xor Codeword(980) xor
                Codeword(1040) xor Codeword(1061) xor Codeword(1252) xor Codeword(1320) xor
                Codeword(1362) xor Codeword(1407) xor Codeword(1491) xor Codeword(1562) xor
                Codeword(1589) xor Codeword(1716) xor Codeword(1726) xor Codeword(1780) xor
                Codeword(1790) xor Codeword(1852) xor Codeword(1862) xor Codeword(1899) xor
                Codeword(1904) xor Codeword(1958) xor Codeword(2006) xor Codeword(2009);
 
     check121 <= Codeword(64) xor Codeword(161) xor Codeword(217) xor Codeword(236) xor
                Codeword(291) xor Codeword(350) xor Codeword(411) xor Codeword(466) xor
                Codeword(566) xor Codeword(628) xor Codeword(670) xor Codeword(767) xor
                Codeword(819) xor Codeword(901) xor Codeword(959) xor Codeword(1017) xor
                Codeword(1083) xor Codeword(1137) xor Codeword(1189) xor Codeword(1223) xor
                Codeword(1249) xor Codeword(1296) xor Codeword(1348) xor Codeword(1411) xor
                Codeword(1479) xor Codeword(1501) xor Codeword(1572) xor Codeword(1646) xor
                Codeword(1696) xor Codeword(1723) xor Codeword(1766) xor Codeword(1829);
 
     check122 <= Codeword(91) xor Codeword(114) xor Codeword(201) xor Codeword(241) xor
                Codeword(327) xor Codeword(375) xor Codeword(475) xor Codeword(551) xor
                Codeword(607) xor Codeword(637) xor Codeword(686) xor Codeword(768) xor
                Codeword(815) xor Codeword(898) xor Codeword(962) xor Codeword(1036) xor
                Codeword(1128) xor Codeword(1182) xor Codeword(1264) xor Codeword(1328) xor
                Codeword(1379) xor Codeword(1400) xor Codeword(1565) xor Codeword(1673) xor
                Codeword(1760) xor Codeword(1771) xor Codeword(1774) xor Codeword(1789) xor
                Codeword(1865) xor Codeword(1928) xor Codeword(1990) xor Codeword(1991);
 
     check123 <= Codeword(82) xor Codeword(122) xor Codeword(213) xor Codeword(279) xor
                Codeword(382) xor Codeword(428) xor Codeword(470) xor Codeword(512) xor
                Codeword(569) xor Codeword(630) xor Codeword(716) xor Codeword(849) xor
                Codeword(914) xor Codeword(946) xor Codeword(1008) xor Codeword(1091) xor
                Codeword(1110) xor Codeword(1115) xor Codeword(1297) xor Codeword(1344) xor
                Codeword(1543) xor Codeword(1569) xor Codeword(1600) xor Codeword(1636) xor
                Codeword(1682) xor Codeword(1722) xor Codeword(1814) xor Codeword(1838) xor
                Codeword(1868) xor Codeword(1876) xor Codeword(1987) xor Codeword(1988);
 
     check124 <= Codeword(69) xor Codeword(153) xor Codeword(240) xor Codeword(292) xor
                Codeword(364) xor Codeword(414) xor Codeword(476) xor Codeword(542) xor
                Codeword(634) xor Codeword(886) xor Codeword(907) xor Codeword(1049) xor
                Codeword(1109) xor Codeword(1133) xor Codeword(1234) xor Codeword(1308) xor
                Codeword(1370) xor Codeword(1419) xor Codeword(1457) xor Codeword(1597) xor
                Codeword(1608) xor Codeword(1721) xor Codeword(1795) xor Codeword(1821) xor
                Codeword(1843) xor Codeword(1856) xor Codeword(1898) xor Codeword(1910) xor
                Codeword(1932) xor Codeword(1962) xor Codeword(1970) xor Codeword(1976);
 
     check125 <= Codeword(87) xor Codeword(169) xor Codeword(320) xor Codeword(366) xor
                Codeword(431) xor Codeword(465) xor Codeword(539) xor Codeword(596) xor
                Codeword(625) xor Codeword(753) xor Codeword(800) xor Codeword(837) xor
                Codeword(936) xor Codeword(1001) xor Codeword(1019) xor Codeword(1078) xor
                Codeword(1113) xor Codeword(1304) xor Codeword(1356) xor Codeword(1434) xor
                Codeword(1493) xor Codeword(1510) xor Codeword(1539) xor Codeword(1692) xor
                Codeword(1719) xor Codeword(1738) xor Codeword(1784) xor Codeword(1816) xor
                Codeword(1859) xor Codeword(1896) xor Codeword(1959) xor Codeword(1964);
 
     check126 <= Codeword(60) xor Codeword(139) xor Codeword(186) xor Codeword(271) xor
                Codeword(281) xor Codeword(334) xor Codeword(394) xor Codeword(487) xor
                Codeword(555) xor Codeword(660) xor Codeword(720) xor Codeword(758) xor
                Codeword(779) xor Codeword(860) xor Codeword(890) xor Codeword(971) xor
                Codeword(1010) xor Codeword(1079) xor Codeword(1162) xor Codeword(1237) xor
                Codeword(1276) xor Codeword(1323) xor Codeword(1334) xor Codeword(1381) xor
                Codeword(1515) xor Codeword(1549) xor Codeword(1586) xor Codeword(1635) xor
                Codeword(1720) xor Codeword(1757) xor Codeword(1764) xor Codeword(1830);
 
     check127 <= Codeword(52) xor Codeword(57) xor Codeword(117) xor Codeword(173) xor
                Codeword(277) xor Codeword(306) xor Codeword(373) xor Codeword(403) xor
                Codeword(494) xor Codeword(548) xor Codeword(597) xor Codeword(644) xor
                Codeword(697) xor Codeword(825) xor Codeword(858) xor Codeword(940) xor
                Codeword(955) xor Codeword(1054) xor Codeword(1120) xor Codeword(1210) xor
                Codeword(1221) xor Codeword(1240) xor Codeword(1292) xor Codeword(1372) xor
                Codeword(1414) xor Codeword(1430) xor Codeword(1499) xor Codeword(1506) xor
                Codeword(1587) xor Codeword(1618) xor Codeword(1706) xor Codeword(1755);
 
     check128 <= Codeword(53) xor Codeword(108) xor Codeword(129) xor Codeword(198) xor
                Codeword(244) xor Codeword(298) xor Codeword(341) xor Codeword(391) xor
                Codeword(441) xor Codeword(457) xor Codeword(534) xor Codeword(579) xor
                Codeword(640) xor Codeword(710) xor Codeword(762) xor Codeword(795) xor
                Codeword(858) xor Codeword(893) xor Codeword(1002) xor Codeword(1037) xor
                Codeword(1073) xor Codeword(1157) xor Codeword(1170) xor Codeword(1244) xor
                Codeword(1286) xor Codeword(1345) xor Codeword(1493) xor Codeword(1573) xor
                Codeword(1581) xor Codeword(1707) xor Codeword(1781) xor Codeword(1831);
 
     check129 <= Codeword(51) xor Codeword(56) xor Codeword(116) xor Codeword(172) xor
                Codeword(276) xor Codeword(305) xor Codeword(372) xor Codeword(402) xor
                Codeword(493) xor Codeword(547) xor Codeword(596) xor Codeword(643) xor
                Codeword(696) xor Codeword(824) xor Codeword(857) xor Codeword(939) xor
                Codeword(954) xor Codeword(1053) xor Codeword(1107) xor Codeword(1119) xor
                Codeword(1209) xor Codeword(1220) xor Codeword(1291) xor Codeword(1371) xor
                Codeword(1413) xor Codeword(1429) xor Codeword(1499) xor Codeword(1586) xor
                Codeword(1617) xor Codeword(1655) xor Codeword(1705) xor Codeword(1756);
 
     check130 <= Codeword(50) xor Codeword(73) xor Codeword(140) xor Codeword(188) xor
                Codeword(245) xor Codeword(285) xor Codeword(385) xor Codeword(398) xor
                Codeword(477) xor Codeword(520) xor Codeword(586) xor Codeword(654) xor
                Codeword(706) xor Codeword(756) xor Codeword(786) xor Codeword(835) xor
                Codeword(981) xor Codeword(1014) xor Codeword(1099) xor Codeword(1189) xor
                Codeword(1230) xor Codeword(1292) xor Codeword(1359) xor Codeword(1401) xor
                Codeword(1439) xor Codeword(1465) xor Codeword(1513) xor Codeword(1556) xor
                Codeword(1620) xor Codeword(1718) xor Codeword(1773) xor Codeword(1832);
 
     check131 <= Codeword(65) xor Codeword(154) xor Codeword(206) xor Codeword(243) xor
                Codeword(307) xor Codeword(334) xor Codeword(403) xor Codeword(479) xor
                Codeword(530) xor Codeword(608) xor Codeword(665) xor Codeword(700) xor
                Codeword(750) xor Codeword(791) xor Codeword(870) xor Codeword(887) xor
                Codeword(932) xor Codeword(972) xor Codeword(1044) xor Codeword(1064) xor
                Codeword(1143) xor Codeword(1173) xor Codeword(1264) xor Codeword(1321) xor
                Codeword(1377) xor Codeword(1551) xor Codeword(1572) xor Codeword(1605) xor
                Codeword(1608) xor Codeword(1674) xor Codeword(1792) xor Codeword(1833);
 
     check132 <= Codeword(49) xor Codeword(151) xor Codeword(214) xor Codeword(274) xor
                Codeword(321) xor Codeword(364) xor Codeword(448) xor Codeword(615) xor
                Codeword(637) xor Codeword(704) xor Codeword(733) xor Codeword(873) xor
                Codeword(914) xor Codeword(959) xor Codeword(1041) xor Codeword(1185) xor
                Codeword(1247) xor Codeword(1352) xor Codeword(1404) xor Codeword(1482) xor
                Codeword(1500) xor Codeword(1560) xor Codeword(1635) xor Codeword(1778) xor
                Codeword(1809) xor Codeword(1940) xor Codeword(1947) xor Codeword(1982) xor
                Codeword(2017) xor Codeword(2042) xor Codeword(2044) xor Codeword(2047);
 
     check133 <= Codeword(48) xor Codeword(209) xor Codeword(255) xor Codeword(317) xor
                Codeword(380) xor Codeword(416) xor Codeword(527) xor Codeword(600) xor
                Codeword(626) xor Codeword(693) xor Codeword(740) xor Codeword(790) xor
                Codeword(860) xor Codeword(896) xor Codeword(978) xor Codeword(1058) xor
                Codeword(1147) xor Codeword(1194) xor Codeword(1259) xor Codeword(1349) xor
                Codeword(1423) xor Codeword(1441) xor Codeword(1509) xor Codeword(1528) xor
                Codeword(1555) xor Codeword(1577) xor Codeword(1675) xor Codeword(1878) xor
                Codeword(1929) xor Codeword(1938) xor Codeword(1945) xor Codeword(1952);
 
     check134 <= Codeword(47) xor Codeword(100) xor Codeword(134) xor Codeword(258) xor
                Codeword(423) xor Codeword(497) xor Codeword(518) xor Codeword(763) xor
                Codeword(950) xor Codeword(1050) xor Codeword(1068) xor Codeword(1151) xor
                Codeword(1271) xor Codeword(1281) xor Codeword(1284) xor Codeword(1607) xor
                Codeword(1628) xor Codeword(1668) xor Codeword(1694) xor Codeword(1750) xor
                Codeword(1787) xor Codeword(1850) xor Codeword(1856) xor Codeword(1869) xor
                Codeword(1880) xor Codeword(1941) xor Codeword(1964) xor Codeword(1965) xor
                Codeword(2001) xor Codeword(2008) xor Codeword(2014) xor Codeword(2023);
 
     check135 <= Codeword(46) xor Codeword(103) xor Codeword(135) xor Codeword(205) xor
                Codeword(388) xor Codeword(449) xor Codeword(555) xor Codeword(571) xor
                Codeword(712) xor Codeword(761) xor Codeword(821) xor Codeword(920) xor
                Codeword(947) xor Codeword(1062) xor Codeword(1140) xor Codeword(1211) xor
                Codeword(1357) xor Codeword(1387) xor Codeword(1447) xor Codeword(1487) xor
                Codeword(1532) xor Codeword(1537) xor Codeword(1686) xor Codeword(1816) xor
                Codeword(1817) xor Codeword(1824) xor Codeword(1846) xor Codeword(1851) xor
                Codeword(1886) xor Codeword(1994) xor Codeword(2005) xor Codeword(2010);
 
     check136 <= Codeword(45) xor Codeword(94) xor Codeword(111) xor Codeword(175) xor
                Codeword(275) xor Codeword(301) xor Codeword(352) xor Codeword(408) xor
                Codeword(478) xor Codeword(537) xor Codeword(607) xor Codeword(649) xor
                Codeword(670) xor Codeword(738) xor Codeword(827) xor Codeword(882) xor
                Codeword(890) xor Codeword(1097) xor Codeword(1120) xor Codeword(1197) xor
                Codeword(1232) xor Codeword(1283) xor Codeword(1451) xor Codeword(1480) xor
                Codeword(1540) xor Codeword(1636) xor Codeword(1777) xor Codeword(1845) xor
                Codeword(1894) xor Codeword(1939) xor Codeword(1949) xor Codeword(1953);
 
     check137 <= Codeword(44) xor Codeword(74) xor Codeword(161) xor Codeword(182) xor
                Codeword(242) xor Codeword(282) xor Codeword(366) xor Codeword(434) xor
                Codeword(492) xor Codeword(551) xor Codeword(564) xor Codeword(656) xor
                Codeword(679) xor Codeword(774) xor Codeword(796) xor Codeword(934) xor
                Codeword(956) xor Codeword(1028) xor Codeword(1103) xor Codeword(1160) xor
                Codeword(1213) xor Codeword(1274) xor Codeword(1341) xor Codeword(1422) xor
                Codeword(1427) xor Codeword(1526) xor Codeword(1678) xor Codeword(1693) xor
                Codeword(1724) xor Codeword(1731) xor Codeword(1893) xor Codeword(1909);
 
     check138 <= Codeword(43) xor Codeword(55) xor Codeword(120) xor Codeword(218) xor
                Codeword(268) xor Codeword(327) xor Codeword(362) xor Codeword(414) xor
                Codeword(466) xor Codeword(506) xor Codeword(572) xor Codeword(653) xor
                Codeword(707) xor Codeword(776) xor Codeword(794) xor Codeword(837) xor
                Codeword(922) xor Codeword(989) xor Codeword(1031) xor Codeword(1074) xor
                Codeword(1115) xor Codeword(1177) xor Codeword(1310) xor Codeword(1431) xor
                Codeword(1450) xor Codeword(1461) xor Codeword(1618) xor Codeword(1680) xor
                Codeword(1712) xor Codeword(1744) xor Codeword(1794) xor Codeword(1834);
 
     check139 <= Codeword(42) xor Codeword(69) xor Codeword(124) xor Codeword(220) xor
                Codeword(252) xor Codeword(289) xor Codeword(383) xor Codeword(426) xor
                Codeword(500) xor Codeword(531) xor Codeword(601) xor Codeword(657) xor
                Codeword(695) xor Codeword(884) xor Codeword(937) xor Codeword(999) xor
                Codeword(1022) xor Codeword(1072) xor Codeword(1126) xor Codeword(1186) xor
                Codeword(1253) xor Codeword(1317) xor Codeword(1338) xor Codeword(1386) xor
                Codeword(1396) xor Codeword(1445) xor Codeword(1582) xor Codeword(1633) xor
                Codeword(1746) xor Codeword(1779) xor Codeword(1815) xor Codeword(1881);
 
     check140 <= Codeword(41) xor Codeword(80) xor Codeword(170) xor Codeword(191) xor
                Codeword(277) xor Codeword(293) xor Codeword(346) xor Codeword(435) xor
                Codeword(467) xor Codeword(519) xor Codeword(614) xor Codeword(648) xor
                Codeword(681) xor Codeword(739) xor Codeword(806) xor Codeword(871) xor
                Codeword(902) xor Codeword(992) xor Codeword(1101) xor Codeword(1154) xor
                Codeword(1182) xor Codeword(1261) xor Codeword(1278) xor Codeword(1287) xor
                Codeword(1467) xor Codeword(1504) xor Codeword(1533) xor Codeword(1544) xor
                Codeword(1580) xor Codeword(1611) xor Codeword(1708) xor Codeword(1757);
 
     check141 <= Codeword(123) xor Codeword(173) xor Codeword(269) xor Codeword(332) xor
                Codeword(347) xor Codeword(407) xor Codeword(480) xor Codeword(508) xor
                Codeword(618) xor Codeword(698) xor Codeword(760) xor Codeword(809) xor
                Codeword(834) xor Codeword(911) xor Codeword(996) xor Codeword(1040) xor
                Codeword(1085) xor Codeword(1142) xor Codeword(1187) xor Codeword(1332) xor
                Codeword(1364) xor Codeword(1459) xor Codeword(1474) xor Codeword(1546) xor
                Codeword(1741) xor Codeword(1788) xor Codeword(1810) xor Codeword(1814) xor
                Codeword(1848) xor Codeword(1872) xor Codeword(1879) xor Codeword(1910);
 
     check142 <= Codeword(40) xor Codeword(96) xor Codeword(118) xor Codeword(256) xor
                Codeword(382) xor Codeword(422) xor Codeword(522) xor Codeword(567) xor
                Codeword(623) xor Codeword(907) xor Codeword(986) xor Codeword(1054) xor
                Codeword(1129) xor Codeword(1262) xor Codeword(1315) xor Codeword(1348) xor
                Codeword(1408) xor Codeword(1623) xor Codeword(1658) xor Codeword(1747) xor
                Codeword(1797) xor Codeword(1818) xor Codeword(1827) xor Codeword(1873) xor
                Codeword(1899) xor Codeword(1902) xor Codeword(1918) xor Codeword(1955) xor
                Codeword(1973) xor Codeword(1989) xor Codeword(1998) xor Codeword(2003);
 
     check143 <= Codeword(39) xor Codeword(83) xor Codeword(158) xor Codeword(192) xor
                Codeword(273) xor Codeword(287) xor Codeword(373) xor Codeword(394) xor
                Codeword(495) xor Codeword(543) xor Codeword(589) xor Codeword(661) xor
                Codeword(671) xor Codeword(771) xor Codeword(862) xor Codeword(912) xor
                Codeword(964) xor Codeword(1008) xor Codeword(1075) xor Codeword(1145) xor
                Codeword(1199) xor Codeword(1252) xor Codeword(1299) xor Codeword(1360) xor
                Codeword(1391) xor Codeword(1436) xor Codeword(1455) xor Codeword(1592) xor
                Codeword(1615) xor Codeword(1679) xor Codeword(1688) xor Codeword(1758);
 
     check144 <= Codeword(38) xor Codeword(98) xor Codeword(166) xor Codeword(219) xor
                Codeword(249) xor Codeword(324) xor Codeword(333) xor Codeword(429) xor
                Codeword(462) xor Codeword(553) xor Codeword(602) xor Codeword(663) xor
                Codeword(720) xor Codeword(741) xor Codeword(793) xor Codeword(876) xor
                Codeword(901) xor Codeword(946) xor Codeword(1034) xor Codeword(1102) xor
                Codeword(1206) xor Codeword(1301) xor Codeword(1330) xor Codeword(1370) xor
                Codeword(1400) xor Codeword(1511) xor Codeword(1520) xor Codeword(1566) xor
                Codeword(1583) xor Codeword(1643) xor Codeword(1785) xor Codeword(1835);
 
     check145 <= Codeword(37) xor Codeword(61) xor Codeword(130) xor Codeword(181) xor
                Codeword(247) xor Codeword(331) xor Codeword(336) xor Codeword(396) xor
                Codeword(463) xor Codeword(548) xor Codeword(599) xor Codeword(631) xor
                Codeword(672) xor Codeword(732) xor Codeword(819) xor Codeword(868) xor
                Codeword(925) xor Codeword(960) xor Codeword(1024) xor Codeword(1071) xor
                Codeword(1117) xor Codeword(1165) xor Codeword(1191) xor Codeword(1227) xor
                Codeword(1288) xor Codeword(1342) xor Codeword(1409) xor Codeword(1442) xor
                Codeword(1460) xor Codeword(1492) xor Codeword(1669) xor Codeword(1759);
 
     check146 <= Codeword(36) xor Codeword(71) xor Codeword(128) xor Codeword(261) xor
                Codeword(299) xor Codeword(494) xor Codeword(562) xor Codeword(716) xor
                Codeword(775) xor Codeword(803) xor Codeword(845) xor Codeword(971) xor
                Codeword(1011) xor Codeword(1266) xor Codeword(1316) xor Codeword(1457) xor
                Codeword(1496) xor Codeword(1535) xor Codeword(1545) xor Codeword(1646) xor
                Codeword(1654) xor Codeword(1689) xor Codeword(1854) xor Codeword(1890) xor
                Codeword(1946) xor Codeword(1948) xor Codeword(1972) xor Codeword(1980) xor
                Codeword(1991) xor Codeword(1997) xor Codeword(2032) xor Codeword(2039);
 
     check147 <= Codeword(35) xor Codeword(66) xor Codeword(164) xor Codeword(187) xor
                Codeword(253) xor Codeword(297) xor Codeword(335) xor Codeword(406) xor
                Codeword(485) xor Codeword(542) xor Codeword(583) xor Codeword(625) xor
                Codeword(684) xor Codeword(722) xor Codeword(737) xor Codeword(828) xor
                Codeword(855) xor Codeword(915) xor Codeword(1026) xor Codeword(1081) xor
                Codeword(1118) xor Codeword(1215) xor Codeword(1268) xor Codeword(1285) xor
                Codeword(1373) xor Codeword(1489) xor Codeword(1567) xor Codeword(1600) xor
                Codeword(1739) xor Codeword(1752) xor Codeword(1807) xor Codeword(1836);
 
     check148 <= Codeword(34) xor Codeword(72) xor Codeword(143) xor Codeword(207) xor
                Codeword(231) xor Codeword(329) xor Codeword(390) xor Codeword(424) xor
                Codeword(504) xor Codeword(510) xor Codeword(584) xor Codeword(632) xor
                Codeword(690) xor Codeword(768) xor Codeword(820) xor Codeword(849) xor
                Codeword(917) xor Codeword(988) xor Codeword(1046) xor Codeword(1104) xor
                Codeword(1198) xor Codeword(1238) xor Codeword(1308) xor Codeword(1331) xor
                Codeword(1335) xor Codeword(1424) xor Codeword(1435) xor Codeword(1510) xor
                Codeword(1589) xor Codeword(1640) xor Codeword(1803) xor Codeword(1837);
 
     check149 <= Codeword(33) xor Codeword(60) xor Codeword(146) xor Codeword(221) xor
                Codeword(241) xor Codeword(309) xor Codeword(370) xor Codeword(446) xor
                Codeword(452) xor Codeword(516) xor Codeword(561) xor Codeword(662) xor
                Codeword(675) xor Codeword(765) xor Codeword(807) xor Codeword(853) xor
                Codeword(941) xor Codeword(974) xor Codeword(1056) xor Codeword(1096) xor
                Codeword(1131) xor Codeword(1210) xor Codeword(1275) xor Codeword(1296) xor
                Codeword(1354) xor Codeword(1403) xor Codeword(1454) xor Codeword(1462) xor
                Codeword(1473) xor Codeword(1624) xor Codeword(1726) xor Codeword(1838);
 
     check150 <= Codeword(32) xor Codeword(86) xor Codeword(131) xor Codeword(217) xor
                Codeword(312) xor Codeword(378) xor Codeword(392) xor Codeword(505) xor
                Codeword(557) xor Codeword(622) xor Codeword(826) xor Codeword(842) xor
                Codeword(923) xor Codeword(991) xor Codeword(1051) xor Codeword(1086) xor
                Codeword(1138) xor Codeword(1216) xor Codeword(1231) xor Codeword(1276) xor
                Codeword(1318) xor Codeword(1362) xor Codeword(1388) xor Codeword(1602) xor
                Codeword(1749) xor Codeword(1805) xor Codeword(1847) xor Codeword(1858) xor
                Codeword(1859) xor Codeword(1911) xor Codeword(1925) xor Codeword(1930);
 
     check151 <= Codeword(31) xor Codeword(92) xor Codeword(165) xor Codeword(184) xor
                Codeword(238) xor Codeword(342) xor Codeword(451) xor Codeword(570) xor
                Codeword(650) xor Codeword(702) xor Codeword(800) xor Codeword(933) xor
                Codeword(952) xor Codeword(1057) xor Codeword(1110) xor Codeword(1192) xor
                Codeword(1239) xor Codeword(1547) xor Codeword(1562) xor Codeword(1619) xor
                Codeword(1667) xor Codeword(1714) xor Codeword(1822) xor Codeword(1864) xor
                Codeword(1867) xor Codeword(1912) xor Codeword(1950) xor Codeword(2021) xor
                Codeword(2029) xor Codeword(2031) xor Codeword(2034) xor Codeword(2041);
 
     check152 <= Codeword(30) xor Codeword(76) xor Codeword(127) xor Codeword(202) xor
                Codeword(228) xor Codeword(330) xor Codeword(340) xor Codeword(415) xor
                Codeword(502) xor Codeword(525) xor Codeword(575) xor Codeword(628) xor
                Codeword(682) xor Codeword(748) xor Codeword(798) xor Codeword(861) xor
                Codeword(942) xor Codeword(962) xor Codeword(1045) xor Codeword(1079) xor
                Codeword(1123) xor Codeword(1205) xor Codeword(1267) xor Codeword(1300) xor
                Codeword(1363) xor Codeword(1390) xor Codeword(1458) xor Codeword(1543) xor
                Codeword(1711) xor Codeword(1742) xor Codeword(1802) xor Codeword(1839);
 
     check153 <= Codeword(29) xor Codeword(78) xor Codeword(155) xor Codeword(203) xor
                Codeword(262) xor Codeword(296) xor Codeword(376) xor Codeword(433) xor
                Codeword(509) xor Codeword(616) xor Codeword(652) xor Codeword(694) xor
                Codeword(758) xor Codeword(812) xor Codeword(872) xor Codeword(916) xor
                Codeword(957) xor Codeword(1077) xor Codeword(1149) xor Codeword(1178) xor
                Codeword(1226) xor Codeword(1314) xor Codeword(1353) xor Codeword(1398) xor
                Codeword(1437) xor Codeword(1484) xor Codeword(1553) xor Codeword(1587) xor
                Codeword(1651) xor Codeword(1699) xor Codeword(1729) xor Codeword(1840);
 
     check154 <= Codeword(28) xor Codeword(139) xor Codeword(183) xor Codeword(246) xor
                Codeword(322) xor Codeword(490) xor Codeword(574) xor Codeword(703) xor
                Codeword(751) xor Codeword(805) xor Codeword(883) xor Codeword(930) xor
                Codeword(963) xor Codeword(1020) xor Codeword(1166) xor Codeword(1254) xor
                Codeword(1376) xor Codeword(1420) xor Codeword(1434) xor Codeword(1584) xor
                Codeword(1642) xor Codeword(1685) xor Codeword(1706) xor Codeword(1855) xor
                Codeword(1868) xor Codeword(1891) xor Codeword(1942) xor Codeword(1999) xor
                Codeword(2013) xor Codeword(2015) xor Codeword(2045) xor Codeword(2046);
 
     check155 <= Codeword(27) xor Codeword(84) xor Codeword(167) xor Codeword(174) xor
                Codeword(257) xor Codeword(306) xor Codeword(357) xor Codeword(447) xor
                Codeword(458) xor Codeword(526) xor Codeword(569) xor Codeword(660) xor
                Codeword(676) xor Codeword(755) xor Codeword(782) xor Codeword(856) xor
                Codeword(903) xor Codeword(951) xor Codeword(1005) xor Codeword(1083) xor
                Codeword(1141) xor Codeword(1180) xor Codeword(1234) xor Codeword(1290) xor
                Codeword(1329) xor Codeword(1382) xor Codeword(1421) xor Codeword(1456) xor
                Codeword(1595) xor Codeword(1657) xor Codeword(1702) xor Codeword(1760);
 
     check156 <= Codeword(26) xor Codeword(95) xor Codeword(157) xor Codeword(343) xor
                Codeword(437) xor Codeword(456) xor Codeword(558) xor Codeword(605) xor
                Codeword(745) xor Codeword(844) xor Codeword(936) xor Codeword(977) xor
                Codeword(1003) xor Codeword(1006) xor Codeword(1150) xor Codeword(1255) xor
                Codeword(1303) xor Codeword(1366) xor Codeword(1397) xor Codeword(1508) xor
                Codeword(1644) xor Codeword(1661) xor Codeword(1728) xor Codeword(1789) xor
                Codeword(1913) xor Codeword(1921) xor Codeword(1936) xor Codeword(1971) xor
                Codeword(1975) xor Codeword(1984) xor Codeword(2019) xor Codeword(2022);
 
     check157 <= Codeword(25) xor Codeword(102) xor Codeword(144) xor Codeword(194) xor
                Codeword(323) xor Codeword(377) xor Codeword(431) xor Codeword(488) xor
                Codeword(515) xor Codeword(612) xor Codeword(645) xor Codeword(717) xor
                Codeword(725) xor Codeword(785) xor Codeword(830) xor Codeword(886) xor
                Codeword(905) xor Codeword(983) xor Codeword(1029) xor Codeword(1069) xor
                Codeword(1122) xor Codeword(1190) xor Codeword(1269) xor Codeword(1297) xor
                Codeword(1368) xor Codeword(1384) xor Codeword(1392) xor Codeword(1477) xor
                Codeword(1612) xor Codeword(1687) xor Codeword(1696) xor Codeword(1761);
 
     check158 <= Codeword(24) xor Codeword(77) xor Codeword(163) xor Codeword(224) xor
                Codeword(230) xor Codeword(310) xor Codeword(339) xor Codeword(412) xor
                Codeword(470) xor Codeword(544) xor Codeword(580) xor Codeword(646) xor
                Codeword(697) xor Codeword(764) xor Codeword(789) xor Codeword(847) xor
                Codeword(918) xor Codeword(966) xor Codeword(1012) xor Codeword(1063) xor
                Codeword(1137) xor Codeword(1208) xor Codeword(1218) xor Codeword(1265) xor
                Codeword(1326) xor Codeword(1337) xor Codeword(1407) xor Codeword(1475) xor
                Codeword(1578) xor Codeword(1621) xor Codeword(1660) xor Codeword(1762);
 
     check159 <= Codeword(23) xor Codeword(91) xor Codeword(136) xor Codeword(271) xor
                Codeword(367) xor Codeword(420) xor Codeword(473) xor Codeword(521) xor
                Codeword(578) xor Codeword(624) xor Codeword(866) xor Codeword(968) xor
                Codeword(1023) xor Codeword(1067) xor Codeword(1113) xor Codeword(1229) xor
                Codeword(1374) xor Codeword(1481) xor Codeword(1512) xor Codeword(1616) xor
                Codeword(1735) xor Codeword(1755) xor Codeword(1775) xor Codeword(1900) xor
                Codeword(1951) xor Codeword(1956) xor Codeword(1958) xor Codeword(1967) xor
                Codeword(1969) xor Codeword(1974) xor Codeword(1985) xor Codeword(1987);
 
     check160 <= Codeword(22) xor Codeword(62) xor Codeword(133) xor Codeword(189) xor
                Codeword(233) xor Codeword(302) xor Codeword(351) xor Codeword(442) xor
                Codeword(459) xor Codeword(546) xor Codeword(610) xor Codeword(617) xor
                Codeword(677) xor Codeword(731) xor Codeword(813) xor Codeword(874) xor
                Codeword(931) xor Codeword(994) xor Codeword(1030) xor Codeword(1109) xor
                Codeword(1144) xor Codeword(1175) xor Codeword(1249) xor Codeword(1443) xor
                Codeword(1527) xor Codeword(1534) xor Codeword(1552) xor Codeword(1565) xor
                Codeword(1576) xor Codeword(1622) xor Codeword(1683) xor Codeword(1763);
 
     check161 <= Codeword(21) xor Codeword(97) xor Codeword(149) xor Codeword(171) xor
                Codeword(250) xor Codeword(300) xor Codeword(379) xor Codeword(440) xor
                Codeword(489) xor Codeword(559) xor Codeword(630) xor Codeword(674) xor
                Codeword(759) xor Codeword(797) xor Codeword(869) xor Codeword(898) xor
                Codeword(975) xor Codeword(1207) xor Codeword(1250) xor Codeword(1411) xor
                Codeword(1452) xor Codeword(1531) xor Codeword(1570) xor Codeword(1650) xor
                Codeword(1743) xor Codeword(1745) xor Codeword(1784) xor Codeword(1790) xor
                Codeword(1823) xor Codeword(1830) xor Codeword(1861) xor Codeword(1882);
 
     check162 <= Codeword(20) xor Codeword(64) xor Codeword(141) xor Codeword(179) xor
                Codeword(259) xor Codeword(315) xor Codeword(369) xor Codeword(418) xor
                Codeword(455) xor Codeword(556) xor Codeword(594) xor Codeword(635) xor
                Codeword(692) xor Codeword(747) xor Codeword(808) xor Codeword(875) xor
                Codeword(899) xor Codeword(987) xor Codeword(1019) xor Codeword(1076) xor
                Codeword(1124) xor Codeword(1228) xor Codeword(1323) xor Codeword(1367) xor
                Codeword(1405) xor Codeword(1446) xor Codeword(1575) xor Codeword(1632) xor
                Codeword(1664) xor Codeword(1725) xor Codeword(1919) xor Codeword(1923);
 
     check163 <= Codeword(19) xor Codeword(79) xor Codeword(115) xor Codeword(254) xor
                Codeword(355) xor Codeword(399) xor Codeword(481) xor Codeword(517) xor
                Codeword(581) xor Codeword(668) xor Codeword(734) xor Codeword(865) xor
                Codeword(995) xor Codeword(1047) xor Codeword(1087) xor Codeword(1121) xor
                Codeword(1381) xor Codeword(1550) xor Codeword(1569) xor Codeword(1637) xor
                Codeword(1663) xor Codeword(1698) xor Codeword(1801) xor Codeword(1874) xor
                Codeword(1896) xor Codeword(1907) xor Codeword(1915) xor Codeword(1960) xor
                Codeword(1976) xor Codeword(1979) xor Codeword(2006) xor Codeword(2011);
 
     check164 <= Codeword(18) xor Codeword(75) xor Codeword(125) xor Codeword(197) xor
                Codeword(260) xor Codeword(375) xor Codeword(401) xor Codeword(539) xor
                Codeword(611) xor Codeword(634) xor Codeword(714) xor Codeword(749) xor
                Codeword(792) xor Codeword(833) xor Codeword(924) xor Codeword(967) xor
                Codeword(1025) xor Codeword(1095) xor Codeword(1139) xor Codeword(1237) xor
                Codeword(1289) xor Codeword(1394) xor Codeword(1494) xor Codeword(1516) xor
                Codeword(1557) xor Codeword(1563) xor Codeword(1690) xor Codeword(1732) xor
                Codeword(1826) xor Codeword(1897) xor Codeword(1914) xor Codeword(1916);
 
     check165 <= Codeword(17) xor Codeword(93) xor Codeword(119) xor Codeword(177) xor
                Codeword(294) xor Codeword(348) xor Codeword(443) xor Codeword(491) xor
                Codeword(540) xor Codeword(629) xor Codeword(691) xor Codeword(769) xor
                Codeword(781) xor Codeword(839) xor Codeword(940) xor Codeword(982) xor
                Codeword(1049) xor Codeword(1070) xor Codeword(1162) xor Codeword(1219) xor
                Codeword(1416) xor Codeword(1440) xor Codeword(1519) xor Codeword(1601) xor
                Codeword(1701) xor Codeword(1780) xor Codeword(1806) xor Codeword(1811) xor
                Codeword(1906) xor Codeword(1917) xor Codeword(2018) xor Codeword(2026);
 
     check166 <= Codeword(16) xor Codeword(57) xor Codeword(122) xor Codeword(210) xor
                Codeword(288) xor Codeword(345) xor Codeword(419) xor Codeword(483) xor
                Codeword(667) xor Codeword(683) xor Codeword(723) xor Codeword(777) xor
                Codeword(822) xor Codeword(878) xor Codeword(888) xor Codeword(953) xor
                Codeword(1007) xor Codeword(1111) xor Codeword(1163) xor Codeword(1309) xor
                Codeword(1356) xor Codeword(1415) xor Codeword(1471) xor Codeword(1515) xor
                Codeword(1525) xor Codeword(1579) xor Codeword(1673) xor Codeword(1709) xor
                Codeword(1808) xor Codeword(1862) xor Codeword(1863) xor Codeword(1883);
 
     check167 <= Codeword(15) xor Codeword(58) xor Codeword(112) xor Codeword(213) xor
                Codeword(225) xor Codeword(292) xor Codeword(360) xor Codeword(471) xor
                Codeword(588) xor Codeword(701) xor Codeword(773) xor Codeword(784) xor
                Codeword(880) xor Codeword(990) xor Codeword(1004) xor Codeword(1167) xor
                Codeword(1214) xor Codeword(1240) xor Codeword(1369) xor Codeword(1393) xor
                Codeword(1502) xor Codeword(1574) xor Codeword(1630) xor Codeword(1665) xor
                Codeword(1791) xor Codeword(1895) xor Codeword(1927) xor Codeword(1990) xor
                Codeword(2030) xor Codeword(2035) xor Codeword(2037) xor Codeword(2043);
 
     check168 <= Codeword(14) xor Codeword(150) xor Codeword(199) xor Codeword(264) xor
                Codeword(283) xor Codeword(353) xor Codeword(409) xor Codeword(487) xor
                Codeword(524) xor Codeword(613) xor Codeword(641) xor Codeword(705) xor
                Codeword(724) xor Codeword(801) xor Codeword(851) xor Codeword(943) xor
                Codeword(955) xor Codeword(1021) xor Codeword(1061) xor Codeword(1130) xor
                Codeword(1196) xor Codeword(1235) xor Codeword(1277) xor Codeword(1325) xor
                Codeword(1365) xor Codeword(1603) xor Codeword(1641) xor Codeword(1649) xor
                Codeword(1734) xor Codeword(1786) xor Codeword(1996) xor Codeword(2000);
 
     check169 <= Codeword(13) xor Codeword(85) xor Codeword(132) xor Codeword(178) xor
                Codeword(266) xor Codeword(316) xor Codeword(387) xor Codeword(395) xor
                Codeword(529) xor Codeword(604) xor Codeword(639) xor Codeword(810) xor
                Codeword(831) xor Codeword(938) xor Codeword(969) xor Codeword(1042) xor
                Codeword(1148) xor Codeword(1203) xor Codeword(1273) xor Codeword(1311) xor
                Codeword(1453) xor Codeword(1469) xor Codeword(1479) xor Codeword(1488) xor
                Codeword(1498) xor Codeword(1539) xor Codeword(1713) xor Codeword(1751) xor
                Codeword(1819) xor Codeword(1961) xor Codeword(1962) xor Codeword(1977);
 
     check170 <= Codeword(12) xor Codeword(101) xor Codeword(145) xor Codeword(236) xor
                Codeword(337) xor Codeword(421) xor Codeword(461) xor Codeword(592) xor
                Codeword(620) xor Codeword(843) xor Codeword(965) xor Codeword(1043) xor
                Codeword(1088) xor Codeword(1153) xor Codeword(1171) xor Codeword(1328) xor
                Codeword(1350) xor Codeword(1417) xor Codeword(1497) xor Codeword(1524) xor
                Codeword(1588) xor Codeword(1626) xor Codeword(1681) xor Codeword(1800) xor
                Codeword(1804) xor Codeword(1898) xor Codeword(1924) xor Codeword(1959) xor
                Codeword(1986) xor Codeword(1993) xor Codeword(2020) xor Codeword(2025);
 
     check171 <= Codeword(105) xor Codeword(156) xor Codeword(222) xor Codeword(311) xor
                Codeword(411) xor Codeword(476) xor Codeword(528) xor Codeword(609) xor
                Codeword(699) xor Codeword(743) xor Codeword(811) xor Codeword(852) xor
                Codeword(928) xor Codeword(985) xor Codeword(1084) xor Codeword(1245) xor
                Codeword(1279) xor Codeword(1294) xor Codeword(1351) xor Codeword(1430) xor
                Codeword(1514) xor Codeword(1518) xor Codeword(1593) xor Codeword(1692) xor
                Codeword(1730) xor Codeword(1798) xor Codeword(1857) xor Codeword(1889) xor
                Codeword(1892) xor Codeword(1922) xor Codeword(1933) xor Codeword(1937);
 
     check172 <= Codeword(11) xor Codeword(110) xor Codeword(126) xor Codeword(229) xor
                Codeword(400) xor Codeword(468) xor Codeword(523) xor Codeword(585) xor
                Codeword(655) xor Codeword(727) xor Codeword(879) xor Codeword(894) xor
                Codeword(948) xor Codeword(1013) xor Codeword(1089) xor Codeword(1152) xor
                Codeword(1201) xor Codeword(1243) xor Codeword(1383) xor Codeword(1414) xor
                Codeword(1591) xor Codeword(1613) xor Codeword(1754) xor Codeword(1795) xor
                Codeword(1866) xor Codeword(1875) xor Codeword(1908) xor Codeword(1957) xor
                Codeword(1983) xor Codeword(2009) xor Codeword(2027) xor Codeword(2033);
 
     check173 <= Codeword(10) xor Codeword(104) xor Codeword(114) xor Codeword(180) xor
                Codeword(237) xor Codeword(295) xor Codeword(384) xor Codeword(417) xor
                Codeword(499) xor Codeword(642) xor Codeword(688) xor Codeword(729) xor
                Codeword(825) xor Codeword(838) xor Codeword(892) xor Codeword(949) xor
                Codeword(1060) xor Codeword(1146) xor Codeword(1183) xor Codeword(1298) xor
                Codeword(1375) xor Codeword(1470) xor Codeword(1522) xor Codeword(1594) xor
                Codeword(1682) xor Codeword(1716) xor Codeword(1727) xor Codeword(1820) xor
                Codeword(1829) xor Codeword(1853) xor Codeword(1934) xor Codeword(1944);
 
     check174 <= Codeword(9) xor Codeword(99) xor Codeword(159) xor Codeword(265) xor
                Codeword(361) xor Codeword(453) xor Codeword(514) xor Codeword(597) xor
                Codeword(753) xor Codeword(984) xor Codeword(1033) xor Codeword(1100) xor
                Codeword(1128) xor Codeword(1168) xor Codeword(1257) xor Codeword(1302) xor
                Codeword(1336) xor Codeword(1425) xor Codeword(1614) xor Codeword(1671) xor
                Codeword(1736) xor Codeword(1770) xor Codeword(1799) xor Codeword(1849) xor
                Codeword(1877) xor Codeword(1887) xor Codeword(1904) xor Codeword(1966) xor
                Codeword(1970) xor Codeword(1988) xor Codeword(1992) xor Codeword(1995);
 
     check175 <= Codeword(8) xor Codeword(82) xor Codeword(117) xor Codeword(211) xor
                Codeword(278) xor Codeword(325) xor Codeword(344) xor Codeword(445) xor
                Codeword(503) xor Codeword(535) xor Codeword(590) xor Codeword(638) xor
                Codeword(709) xor Codeword(735) xor Codeword(815) xor Codeword(846) xor
                Codeword(908) xor Codeword(976) xor Codeword(1106) xor Codeword(1135) xor
                Codeword(1164) xor Codeword(1172) xor Codeword(1260) xor Codeword(1293) xor
                Codeword(1340) xor Codeword(1395) xor Codeword(1438) xor Codeword(1495) xor
                Codeword(1505) xor Codeword(1606) xor Codeword(1627) xor Codeword(1764);
 
     check176 <= Codeword(7) xor Codeword(89) xor Codeword(137) xor Codeword(176) xor
                Codeword(251) xor Codeword(286) xor Codeword(356) xor Codeword(404) xor
                Codeword(450) xor Codeword(533) xor Codeword(566) xor Codeword(664) xor
                Codeword(686) xor Codeword(746) xor Codeword(817) xor Codeword(867) xor
                Codeword(910) xor Codeword(993) xor Codeword(1032) xor Codeword(1091) xor
                Codeword(1158) xor Codeword(1169) xor Codeword(1202) xor Codeword(1246) xor
                Codeword(1313) xor Codeword(1389) xor Codeword(1464) xor Codeword(1536) xor
                Codeword(1549) xor Codeword(1625) xor Codeword(1691) xor Codeword(1765);
 
     check177 <= Codeword(6) xor Codeword(109) xor Codeword(147) xor Codeword(204) xor
                Codeword(232) xor Codeword(304) xor Codeword(368) xor Codeword(397) xor
                Codeword(496) xor Codeword(512) xor Codeword(576) xor Codeword(651) xor
                Codeword(721) xor Codeword(754) xor Codeword(787) xor Codeword(881) xor
                Codeword(895) xor Codeword(998) xor Codeword(1027) xor Codeword(1059) xor
                Codeword(1093) xor Codeword(1156) xor Codeword(1320) xor Codeword(1339) xor
                Codeword(1472) xor Codeword(1517) xor Codeword(1523) xor Codeword(1538) xor
                Codeword(1597) xor Codeword(1639) xor Codeword(1697) xor Codeword(1766);
 
     check178 <= Codeword(5) xor Codeword(107) xor Codeword(142) xor Codeword(201) xor
                Codeword(313) xor Codeword(338) xor Codeword(428) xor Codeword(549) xor
                Codeword(621) xor Codeword(728) xor Codeword(823) xor Codeword(877) xor
                Codeword(927) xor Codeword(1010) xor Codeword(1065) xor Codeword(1133) xor
                Codeword(1193) xor Codeword(1242) xor Codeword(1282) xor Codeword(1304) xor
                Codeword(1503) xor Codeword(1599) xor Codeword(1609) xor Codeword(1676) xor
                Codeword(1704) xor Codeword(1796) xor Codeword(1813) xor Codeword(1871) xor
                Codeword(1888) xor Codeword(1920) xor Codeword(1963) xor Codeword(1978);
 
     check179 <= Codeword(4) xor Codeword(87) xor Codeword(148) xor Codeword(215) xor
                Codeword(267) xor Codeword(308) xor Codeword(386) xor Codeword(438) xor
                Codeword(460) xor Codeword(552) xor Codeword(573) xor Codeword(666) xor
                Codeword(711) xor Codeword(742) xor Codeword(780) xor Codeword(841) xor
                Codeword(891) xor Codeword(997) xor Codeword(1017) xor Codeword(1098) xor
                Codeword(1114) xor Codeword(1179) xor Codeword(1270) xor Codeword(1306) xor
                Codeword(1372) xor Codeword(1428) xor Codeword(1483) xor Codeword(1610) xor
                Codeword(1670) xor Codeword(1717) xor Codeword(1771) xor Codeword(1841);
 
     check180 <= Codeword(67) xor Codeword(208) xor Codeword(263) xor Codeword(314) xor
                Codeword(371) xor Codeword(432) xor Codeword(472) xor Codeword(536) xor
                Codeword(563) xor Codeword(687) xor Codeword(770) xor Codeword(788) xor
                Codeword(863) xor Codeword(919) xor Codeword(1038) xor Codeword(1116) xor
                Codeword(1204) xor Codeword(1221) xor Codeword(1379) xor Codeword(1419) xor
                Codeword(1468) xor Codeword(1507) xor Codeword(1529) xor Codeword(1604) xor
                Codeword(1638) xor Codeword(1695) xor Codeword(1738) xor Codeword(1885) xor
                Codeword(1901) xor Codeword(1935) xor Codeword(2016) xor Codeword(2024);
 
     check181 <= Codeword(3) xor Codeword(70) xor Codeword(162) xor Codeword(186) xor
                Codeword(227) xor Codeword(303) xor Codeword(389) xor Codeword(436) xor
                Codeword(482) xor Codeword(513) xor Codeword(598) xor Codeword(619) xor
                Codeword(708) xor Codeword(816) xor Codeword(864) xor Codeword(904) xor
                Codeword(973) xor Codeword(1036) xor Codeword(1066) xor Codeword(1159) xor
                Codeword(1195) xor Codeword(1223) xor Codeword(1225) xor Codeword(1312) xor
                Codeword(1346) xor Codeword(1385) xor Codeword(1476) xor Codeword(1541) xor
                Codeword(1631) xor Codeword(1710) xor Codeword(1733) xor Codeword(1842);
 
     check182 <= Codeword(2) xor Codeword(54) xor Codeword(169) xor Codeword(195) xor
                Codeword(248) xor Codeword(328) xor Codeword(350) xor Codeword(425) xor
                Codeword(454) xor Codeword(532) xor Codeword(582) xor Codeword(647) xor
                Codeword(678) xor Codeword(772) xor Codeword(829) xor Codeword(840) xor
                Codeword(929) xor Codeword(1015) xor Codeword(1092) xor Codeword(1134) xor
                Codeword(1184) xor Codeword(1272) xor Codeword(1324) xor Codeword(1334) xor
                Codeword(1344) xor Codeword(1448) xor Codeword(1486) xor Codeword(1647) xor
                Codeword(1656) xor Codeword(1700) xor Codeword(1772) xor Codeword(1843);
 
     check183 <= Codeword(1) xor Codeword(88) xor Codeword(190) xor Codeword(281) xor
                Codeword(358) xor Codeword(405) xor Codeword(498) xor Codeword(560) xor
                Codeword(593) xor Codeword(644) xor Codeword(718) xor Codeword(730) xor
                Codeword(802) xor Codeword(832) xor Codeword(921) xor Codeword(944) xor
                Codeword(1052) xor Codeword(1105) xor Codeword(1155) xor Codeword(1200) xor
                Codeword(1258) xor Codeword(1280) xor Codeword(1402) xor Codeword(1432) xor
                Codeword(1491) xor Codeword(1530) xor Codeword(1598) xor Codeword(1659) xor
                Codeword(1776) xor Codeword(1860) xor Codeword(1926) xor Codeword(1931);
 
     check184 <= Codeword(0) xor Codeword(106) xor Codeword(153) xor Codeword(193) xor
                Codeword(226) xor Codeword(318) xor Codeword(354) xor Codeword(444) xor
                Codeword(484) xor Codeword(545) xor Codeword(603) xor Codeword(658) xor
                Codeword(689) xor Codeword(726) xor Codeword(783) xor Codeword(850) xor
                Codeword(909) xor Codeword(1001) xor Codeword(1055) xor Codeword(1080) xor
                Codeword(1125) xor Codeword(1176) xor Codeword(1305) xor Codeword(1358) xor
                Codeword(1412) xor Codeword(1426) xor Codeword(1463) xor Codeword(1521) xor
                Codeword(1558) xor Codeword(1648) xor Codeword(1652) xor Codeword(1767);
 
     check185 <= Codeword(121) xor Codeword(272) xor Codeword(320) xor Codeword(359) xor
                Codeword(501) xor Codeword(577) xor Codeword(680) xor Codeword(804) xor
                Codeword(926) xor Codeword(979) xor Codeword(1039) xor Codeword(1174) xor
                Codeword(1251) xor Codeword(1319) xor Codeword(1361) xor Codeword(1406) xor
                Codeword(1449) xor Codeword(1490) xor Codeword(1561) xor Codeword(1677) xor
                Codeword(1715) xor Codeword(1723) xor Codeword(1865) xor Codeword(1876) xor
                Codeword(1903) xor Codeword(1943) xor Codeword(1954) xor Codeword(1981) xor
                Codeword(2007) xor Codeword(2012) xor Codeword(2028) xor Codeword(2036);
 
     check186 <= Codeword(63) xor Codeword(160) xor Codeword(216) xor Codeword(235) xor
                Codeword(290) xor Codeword(349) xor Codeword(410) xor Codeword(465) xor
                Codeword(507) xor Codeword(565) xor Codeword(627) xor Codeword(669) xor
                Codeword(766) xor Codeword(818) xor Codeword(900) xor Codeword(958) xor
                Codeword(1016) xor Codeword(1082) xor Codeword(1136) xor Codeword(1188) xor
                Codeword(1222) xor Codeword(1248) xor Codeword(1295) xor Codeword(1347) xor
                Codeword(1410) xor Codeword(1478) xor Codeword(1501) xor Codeword(1571) xor
                Codeword(1645) xor Codeword(1666) xor Codeword(1928) xor Codeword(1932);
 
     check187 <= Codeword(90) xor Codeword(113) xor Codeword(200) xor Codeword(240) xor
                Codeword(326) xor Codeword(374) xor Codeword(439) xor Codeword(474) xor
                Codeword(550) xor Codeword(606) xor Codeword(636) xor Codeword(685) xor
                Codeword(767) xor Codeword(814) xor Codeword(854) xor Codeword(897) xor
                Codeword(961) xor Codeword(1035) xor Codeword(1094) xor Codeword(1127) xor
                Codeword(1181) xor Codeword(1263) xor Codeword(1327) xor Codeword(1378) xor
                Codeword(1399) xor Codeword(1554) xor Codeword(1564) xor Codeword(1590) xor
                Codeword(1629) xor Codeword(1672) xor Codeword(1722) xor Codeword(1768);
 
     check188 <= Codeword(81) xor Codeword(212) xor Codeword(279) xor Codeword(284) xor
                Codeword(381) xor Codeword(427) xor Codeword(469) xor Codeword(511) xor
                Codeword(568) xor Codeword(715) xor Codeword(744) xor Codeword(779) xor
                Codeword(848) xor Codeword(913) xor Codeword(945) xor Codeword(1090) xor
                Codeword(1108) xor Codeword(1212) xor Codeword(1256) xor Codeword(1343) xor
                Codeword(1542) xor Codeword(1568) xor Codeword(1721) xor Codeword(1737) xor
                Codeword(1774) xor Codeword(1783) xor Codeword(1812) xor Codeword(1825) xor
                Codeword(1828) xor Codeword(1852) xor Codeword(1870) xor Codeword(1884);
 
     check189 <= Codeword(68) xor Codeword(152) xor Codeword(223) xor Codeword(239) xor
                Codeword(291) xor Codeword(363) xor Codeword(413) xor Codeword(475) xor
                Codeword(541) xor Codeword(587) xor Codeword(633) xor Codeword(713) xor
                Codeword(736) xor Codeword(799) xor Codeword(885) xor Codeword(906) xor
                Codeword(980) xor Codeword(1048) xor Codeword(1132) xor Codeword(1233) xor
                Codeword(1307) xor Codeword(1418) xor Codeword(1444) xor Codeword(1506) xor
                Codeword(1559) xor Codeword(1596) xor Codeword(1662) xor Codeword(1719) xor
                Codeword(1740) xor Codeword(1748) xor Codeword(1793) xor Codeword(1844);
 
     check190 <= Codeword(168) xor Codeword(196) xor Codeword(234) xor Codeword(319) xor
                Codeword(365) xor Codeword(430) xor Codeword(464) xor Codeword(538) xor
                Codeword(595) xor Codeword(673) xor Codeword(752) xor Codeword(836) xor
                Codeword(935) xor Codeword(1000) xor Codeword(1018) xor Codeword(1112) xor
                Codeword(1241) xor Codeword(1355) xor Codeword(1433) xor Codeword(1466) xor
                Codeword(1485) xor Codeword(1653) xor Codeword(1720) xor Codeword(1753) xor
                Codeword(1782) xor Codeword(1821) xor Codeword(1905) xor Codeword(1968) xor
                Codeword(2002) xor Codeword(2004) xor Codeword(2038) xor Codeword(2040);
 
     check191 <= Codeword(52) xor Codeword(59) xor Codeword(138) xor Codeword(185) xor
                Codeword(270) xor Codeword(280) xor Codeword(393) xor Codeword(486) xor
                Codeword(554) xor Codeword(591) xor Codeword(659) xor Codeword(719) xor
                Codeword(757) xor Codeword(778) xor Codeword(859) xor Codeword(889) xor
                Codeword(970) xor Codeword(1009) xor Codeword(1078) xor Codeword(1161) xor
                Codeword(1217) xor Codeword(1224) xor Codeword(1236) xor Codeword(1322) xor
                Codeword(1333) xor Codeword(1380) xor Codeword(1548) xor Codeword(1585) xor
                Codeword(1634) xor Codeword(1684) xor Codeword(1703) xor Codeword(1769);
 
     check192 <= Codeword(53) xor Codeword(107) xor Codeword(128) xor Codeword(197) xor
                Codeword(243) xor Codeword(297) xor Codeword(340) xor Codeword(440) xor
                Codeword(456) xor Codeword(533) xor Codeword(578) xor Codeword(639) xor
                Codeword(709) xor Codeword(761) xor Codeword(794) xor Codeword(857) xor
                Codeword(892) xor Codeword(1001) xor Codeword(1036) xor Codeword(1072) xor
                Codeword(1156) xor Codeword(1243) xor Codeword(1344) xor Codeword(1415) xor
                Codeword(1455) xor Codeword(1485) xor Codeword(1518) xor Codeword(1580) xor
                Codeword(1663) xor Codeword(1734) xor Codeword(1788) xor Codeword(1845);
 
     check193 <= Codeword(51) xor Codeword(58) xor Codeword(137) xor Codeword(269) xor
                Codeword(333) xor Codeword(485) xor Codeword(590) xor Codeword(658) xor
                Codeword(756) xor Codeword(858) xor Codeword(888) xor Codeword(969) xor
                Codeword(1008) xor Codeword(1160) xor Codeword(1216) xor Codeword(1223) xor
                Codeword(1235) xor Codeword(1321) xor Codeword(1379) xor Codeword(1584) xor
                Codeword(1633) xor Codeword(1683) xor Codeword(1702) xor Codeword(1877) xor
                Codeword(1899) xor Codeword(1944) xor Codeword(1985) xor Codeword(2022) xor
                Codeword(2027) xor Codeword(2032) xor Codeword(2040) xor Codeword(2042);
 
     check194 <= Codeword(50) xor Codeword(55) xor Codeword(115) xor Codeword(171) xor
                Codeword(275) xor Codeword(304) xor Codeword(371) xor Codeword(401) xor
                Codeword(492) xor Codeword(546) xor Codeword(595) xor Codeword(642) xor
                Codeword(695) xor Codeword(823) xor Codeword(938) xor Codeword(953) xor
                Codeword(1052) xor Codeword(1106) xor Codeword(1118) xor Codeword(1208) xor
                Codeword(1219) xor Codeword(1239) xor Codeword(1290) xor Codeword(1370) xor
                Codeword(1412) xor Codeword(1428) xor Codeword(1499) xor Codeword(1585) xor
                Codeword(1616) xor Codeword(1654) xor Codeword(1792) xor Codeword(1846);
 
     check195 <= Codeword(72) xor Codeword(139) xor Codeword(187) xor Codeword(244) xor
                Codeword(384) xor Codeword(397) xor Codeword(519) xor Codeword(585) xor
                Codeword(705) xor Codeword(755) xor Codeword(785) xor Codeword(834) xor
                Codeword(942) xor Codeword(1098) xor Codeword(1188) xor Codeword(1229) xor
                Codeword(1291) xor Codeword(1358) xor Codeword(1400) xor Codeword(1438) xor
                Codeword(1464) xor Codeword(1555) xor Codeword(1619) xor Codeword(1668) xor
                Codeword(1718) xor Codeword(1729) xor Codeword(1732) xor Codeword(1790) xor
                Codeword(1827) xor Codeword(1833) xor Codeword(1843) xor Codeword(1885);
 
     check196 <= Codeword(49) xor Codeword(64) xor Codeword(153) xor Codeword(205) xor
                Codeword(242) xor Codeword(306) xor Codeword(402) xor Codeword(478) xor
                Codeword(529) xor Codeword(664) xor Codeword(699) xor Codeword(749) xor
                Codeword(790) xor Codeword(830) xor Codeword(869) xor Codeword(931) xor
                Codeword(971) xor Codeword(1043) xor Codeword(1063) xor Codeword(1142) xor
                Codeword(1172) xor Codeword(1263) xor Codeword(1320) xor Codeword(1376) xor
                Codeword(1550) xor Codeword(1571) xor Codeword(1604) xor Codeword(1673) xor
                Codeword(1728) xor Codeword(1740) xor Codeword(1769) xor Codeword(1847);
 
     check197 <= Codeword(48) xor Codeword(96) xor Codeword(150) xor Codeword(213) xor
                Codeword(273) xor Codeword(320) xor Codeword(363) xor Codeword(504) xor
                Codeword(523) xor Codeword(614) xor Codeword(636) xor Codeword(703) xor
                Codeword(732) xor Codeword(872) xor Codeword(887) xor Codeword(913) xor
                Codeword(958) xor Codeword(1040) xor Codeword(1068) xor Codeword(1153) xor
                Codeword(1184) xor Codeword(1246) xor Codeword(1312) xor Codeword(1351) xor
                Codeword(1403) xor Codeword(1457) xor Codeword(1481) xor Codeword(1500) xor
                Codeword(1634) xor Codeword(1670) xor Codeword(1701) xor Codeword(1770);
 
     check198 <= Codeword(47) xor Codeword(105) xor Codeword(111) xor Codeword(208) xor
                Codeword(254) xor Codeword(316) xor Codeword(379) xor Codeword(415) xor
                Codeword(484) xor Codeword(526) xor Codeword(599) xor Codeword(625) xor
                Codeword(692) xor Codeword(739) xor Codeword(789) xor Codeword(859) xor
                Codeword(895) xor Codeword(977) xor Codeword(1057) xor Codeword(1146) xor
                Codeword(1193) xor Codeword(1258) xor Codeword(1348) xor Codeword(1422) xor
                Codeword(1440) xor Codeword(1484) xor Codeword(1487) xor Codeword(1509) xor
                Codeword(1527) xor Codeword(1674) xor Codeword(1689) xor Codeword(1771);
 
     check199 <= Codeword(46) xor Codeword(99) xor Codeword(133) xor Codeword(214) xor
                Codeword(257) xor Codeword(282) xor Codeword(350) xor Codeword(422) xor
                Codeword(496) xor Codeword(517) xor Codeword(601) xor Codeword(667) xor
                Codeword(673) xor Codeword(762) xor Codeword(784) xor Codeword(835) xor
                Codeword(909) xor Codeword(949) xor Codeword(1049) xor Codeword(1067) xor
                Codeword(1150) xor Codeword(1270) xor Codeword(1280) xor Codeword(1283) xor
                Codeword(1363) xor Codeword(1539) xor Codeword(1562) xor Codeword(1607) xor
                Codeword(1627) xor Codeword(1748) xor Codeword(1765) xor Codeword(1848);
 
     check200 <= Codeword(45) xor Codeword(102) xor Codeword(134) xor Codeword(204) xor
                Codeword(245) xor Codeword(300) xor Codeword(387) xor Codeword(406) xor
                Codeword(448) xor Codeword(554) xor Codeword(570) xor Codeword(628) xor
                Codeword(711) xor Codeword(760) xor Codeword(820) xor Codeword(856) xor
                Codeword(919) xor Codeword(946) xor Codeword(1024) xor Codeword(1061) xor
                Codeword(1139) xor Codeword(1210) xor Codeword(1241) xor Codeword(1356) xor
                Codeword(1386) xor Codeword(1446) xor Codeword(1532) xor Codeword(1576) xor
                Codeword(1613) xor Codeword(1685) xor Codeword(1707) xor Codeword(1772);
 
     check201 <= Codeword(44) xor Codeword(93) xor Codeword(169) xor Codeword(174) xor
                Codeword(274) xor Codeword(351) xor Codeword(407) xor Codeword(477) xor
                Codeword(536) xor Codeword(606) xor Codeword(648) xor Codeword(669) xor
                Codeword(737) xor Codeword(881) xor Codeword(889) xor Codeword(963) xor
                Codeword(1033) xor Codeword(1096) xor Codeword(1119) xor Codeword(1196) xor
                Codeword(1231) xor Codeword(1430) xor Codeword(1450) xor Codeword(1479) xor
                Codeword(1531) xor Codeword(1535) xor Codeword(1747) xor Codeword(1750) xor
                Codeword(1758) xor Codeword(1812) xor Codeword(1835) xor Codeword(1886);
 
     check202 <= Codeword(43) xor Codeword(73) xor Codeword(160) xor Codeword(181) xor
                Codeword(281) xor Codeword(365) xor Codeword(433) xor Codeword(491) xor
                Codeword(550) xor Codeword(563) xor Codeword(655) xor Codeword(678) xor
                Codeword(773) xor Codeword(795) xor Codeword(933) xor Codeword(955) xor
                Codeword(1027) xor Codeword(1102) xor Codeword(1159) xor Codeword(1273) xor
                Codeword(1328) xor Codeword(1340) xor Codeword(1426) xor Codeword(1602) xor
                Codeword(1724) xor Codeword(1726) xor Codeword(1761) xor Codeword(1803) xor
                Codeword(1839) xor Codeword(1841) xor Codeword(1868) xor Codeword(1887);
 
     check203 <= Codeword(42) xor Codeword(54) xor Codeword(119) xor Codeword(217) xor
                Codeword(267) xor Codeword(326) xor Codeword(361) xor Codeword(413) xor
                Codeword(465) xor Codeword(560) xor Codeword(571) xor Codeword(706) xor
                Codeword(793) xor Codeword(836) xor Codeword(988) xor Codeword(1030) xor
                Codeword(1073) xor Codeword(1234) xor Codeword(1392) xor Codeword(1460) xor
                Codeword(1617) xor Codeword(1679) xor Codeword(1828) xor Codeword(1871) xor
                Codeword(1903) xor Codeword(1912) xor Codeword(1924) xor Codeword(1953) xor
                Codeword(1955) xor Codeword(1956) xor Codeword(2000) xor Codeword(2006);
 
     check204 <= Codeword(41) xor Codeword(68) xor Codeword(123) xor Codeword(219) xor
                Codeword(251) xor Codeword(288) xor Codeword(382) xor Codeword(425) xor
                Codeword(499) xor Codeword(530) xor Codeword(600) xor Codeword(656) xor
                Codeword(694) xor Codeword(763) xor Codeword(826) xor Codeword(883) xor
                Codeword(936) xor Codeword(998) xor Codeword(1021) xor Codeword(1071) xor
                Codeword(1125) xor Codeword(1252) xor Codeword(1316) xor Codeword(1385) xor
                Codeword(1581) xor Codeword(1632) xor Codeword(1657) xor Codeword(1745) xor
                Codeword(1752) xor Codeword(1763) xor Codeword(1795) xor Codeword(1849);
 
     check205 <= Codeword(170) xor Codeword(276) xor Codeword(345) xor Codeword(434) xor
                Codeword(613) xor Codeword(647) xor Codeword(738) xor Codeword(870) xor
                Codeword(901) xor Codeword(1058) xor Codeword(1181) xor Codeword(1260) xor
                Codeword(1286) xor Codeword(1543) xor Codeword(1553) xor Codeword(1610) xor
                Codeword(1684) xor Codeword(1810) xor Codeword(1914) xor Codeword(1967) xor
                Codeword(1977) xor Codeword(1984) xor Codeword(1989) xor Codeword(1994) xor
                Codeword(1997) xor Codeword(2009) xor Codeword(2015) xor Codeword(2016) xor
                Codeword(2025) xor Codeword(2029) xor Codeword(2036) xor Codeword(2044);
 
     check206 <= Codeword(40) xor Codeword(122) xor Codeword(172) xor Codeword(332) xor
                Codeword(346) xor Codeword(479) xor Codeword(587) xor Codeword(617) xor
                Codeword(697) xor Codeword(759) xor Codeword(808) xor Codeword(833) xor
                Codeword(910) xor Codeword(995) xor Codeword(1039) xor Codeword(1084) xor
                Codeword(1141) xor Codeword(1186) xor Codeword(1256) xor Codeword(1285) xor
                Codeword(1331) xor Codeword(1458) xor Codeword(1473) xor Codeword(1545) xor
                Codeword(1652) xor Codeword(1693) xor Codeword(1824) xor Codeword(1829) xor
                Codeword(1869) xor Codeword(1921) xor Codeword(1930) xor Codeword(1938);
 
     check207 <= Codeword(39) xor Codeword(95) xor Codeword(117) xor Codeword(255) xor
                Codeword(292) xor Codeword(381) xor Codeword(391) xor Codeword(421) xor
                Codeword(521) xor Codeword(566) xor Codeword(622) xor Codeword(716) xor
                Codeword(730) xor Codeword(796) xor Codeword(864) xor Codeword(906) xor
                Codeword(985) xor Codeword(1053) xor Codeword(1087) xor Codeword(1128) xor
                Codeword(1176) xor Codeword(1261) xor Codeword(1314) xor Codeword(1347) xor
                Codeword(1407) xor Codeword(1434) xor Codeword(1591) xor Codeword(1622) xor
                Codeword(1725) xor Codeword(1881) xor Codeword(1954) xor Codeword(1963);
 
     check208 <= Codeword(38) xor Codeword(82) xor Codeword(157) xor Codeword(191) xor
                Codeword(286) xor Codeword(372) xor Codeword(393) xor Codeword(494) xor
                Codeword(542) xor Codeword(588) xor Codeword(660) xor Codeword(770) xor
                Codeword(861) xor Codeword(911) xor Codeword(1074) xor Codeword(1144) xor
                Codeword(1251) xor Codeword(1298) xor Codeword(1359) xor Codeword(1435) xor
                Codeword(1454) xor Codeword(1551) xor Codeword(1614) xor Codeword(1678) xor
                Codeword(1767) xor Codeword(1813) xor Codeword(1815) xor Codeword(1862) xor
                Codeword(1884) xor Codeword(1894) xor Codeword(1916) xor Codeword(1919);
 
     check209 <= Codeword(37) xor Codeword(97) xor Codeword(165) xor Codeword(218) xor
                Codeword(323) xor Codeword(428) xor Codeword(461) xor Codeword(552) xor
                Codeword(662) xor Codeword(719) xor Codeword(740) xor Codeword(792) xor
                Codeword(875) xor Codeword(900) xor Codeword(945) xor Codeword(1101) xor
                Codeword(1205) xor Codeword(1329) xor Codeword(1399) xor Codeword(1510) xor
                Codeword(1565) xor Codeword(1582) xor Codeword(1642) xor Codeword(1710) xor
                Codeword(1844) xor Codeword(1880) xor Codeword(1907) xor Codeword(1908) xor
                Codeword(1917) xor Codeword(1922) xor Codeword(1931) xor Codeword(1939);
 
     check210 <= Codeword(36) xor Codeword(60) xor Codeword(129) xor Codeword(180) xor
                Codeword(246) xor Codeword(330) xor Codeword(335) xor Codeword(395) xor
                Codeword(462) xor Codeword(547) xor Codeword(598) xor Codeword(630) xor
                Codeword(671) xor Codeword(731) xor Codeword(818) xor Codeword(867) xor
                Codeword(924) xor Codeword(959) xor Codeword(1023) xor Codeword(1070) xor
                Codeword(1116) xor Codeword(1164) xor Codeword(1190) xor Codeword(1226) xor
                Codeword(1287) xor Codeword(1341) xor Codeword(1408) xor Codeword(1441) xor
                Codeword(1459) xor Codeword(1491) xor Codeword(1694) xor Codeword(1773);
 
     check211 <= Codeword(35) xor Codeword(70) xor Codeword(127) xor Codeword(206) xor
                Codeword(260) xor Codeword(298) xor Codeword(408) xor Codeword(493) xor
                Codeword(553) xor Codeword(561) xor Codeword(715) xor Codeword(774) xor
                Codeword(802) xor Codeword(844) xor Codeword(930) xor Codeword(970) xor
                Codeword(1010) xor Codeword(1094) xor Codeword(1167) xor Codeword(1192) xor
                Codeword(1265) xor Codeword(1315) xor Codeword(1496) xor Codeword(1513) xor
                Codeword(1534) xor Codeword(1544) xor Codeword(1559) xor Codeword(1579) xor
                Codeword(1645) xor Codeword(1738) xor Codeword(1743) xor Codeword(1850);
 
     check212 <= Codeword(34) xor Codeword(65) xor Codeword(163) xor Codeword(186) xor
                Codeword(296) xor Codeword(405) xor Codeword(541) xor Codeword(683) xor
                Codeword(827) xor Codeword(999) xor Codeword(1025) xor Codeword(1080) xor
                Codeword(1117) xor Codeword(1267) xor Codeword(1372) xor Codeword(1395) xor
                Codeword(1488) xor Codeword(1566) xor Codeword(1712) xor Codeword(1730) xor
                Codeword(1737) xor Codeword(1796) xor Codeword(1865) xor Codeword(1875) xor
                Codeword(1895) xor Codeword(1896) xor Codeword(1898) xor Codeword(1900) xor
                Codeword(1902) xor Codeword(1905) xor Codeword(1934) xor Codeword(1945);
 
     check213 <= Codeword(33) xor Codeword(71) xor Codeword(142) xor Codeword(230) xor
                Codeword(389) xor Codeword(503) xor Codeword(583) xor Codeword(631) xor
                Codeword(767) xor Codeword(848) xor Codeword(916) xor Codeword(987) xor
                Codeword(1045) xor Codeword(1103) xor Codeword(1197) xor Codeword(1237) xor
                Codeword(1307) xor Codeword(1330) xor Codeword(1423) xor Codeword(1639) xor
                Codeword(1680) xor Codeword(1692) xor Codeword(1915) xor Codeword(1918) xor
                Codeword(1957) xor Codeword(1974) xor Codeword(1975) xor Codeword(2002) xor
                Codeword(2012) xor Codeword(2018) xor Codeword(2021) xor Codeword(2037);
 
     check214 <= Codeword(32) xor Codeword(59) xor Codeword(145) xor Codeword(220) xor
                Codeword(240) xor Codeword(308) xor Codeword(369) xor Codeword(445) xor
                Codeword(451) xor Codeword(515) xor Codeword(615) xor Codeword(661) xor
                Codeword(674) xor Codeword(764) xor Codeword(806) xor Codeword(852) xor
                Codeword(940) xor Codeword(973) xor Codeword(1055) xor Codeword(1095) xor
                Codeword(1130) xor Codeword(1209) xor Codeword(1274) xor Codeword(1295) xor
                Codeword(1353) xor Codeword(1402) xor Codeword(1453) xor Codeword(1461) xor
                Codeword(1472) xor Codeword(1623) xor Codeword(1677) xor Codeword(1774);
 
     check215 <= Codeword(31) xor Codeword(85) xor Codeword(130) xor Codeword(216) xor
                Codeword(234) xor Codeword(311) xor Codeword(377) xor Codeword(446) xor
                Codeword(505) xor Codeword(556) xor Codeword(607) xor Codeword(621) xor
                Codeword(676) xor Codeword(724) xor Codeword(825) xor Codeword(841) xor
                Codeword(922) xor Codeword(990) xor Codeword(1050) xor Codeword(1085) xor
                Codeword(1137) xor Codeword(1215) xor Codeword(1224) xor Codeword(1230) xor
                Codeword(1317) xor Codeword(1361) xor Codeword(1387) xor Codeword(1425) xor
                Codeword(1601) xor Codeword(1608) xor Codeword(1651) xor Codeword(1775);
 
     check216 <= Codeword(30) xor Codeword(91) xor Codeword(164) xor Codeword(183) xor
                Codeword(237) xor Codeword(299) xor Codeword(341) xor Codeword(423) xor
                Codeword(450) xor Codeword(558) xor Codeword(649) xor Codeword(701) xor
                Codeword(772) xor Codeword(876) xor Codeword(932) xor Codeword(951) xor
                Codeword(1056) xor Codeword(1100) xor Codeword(1108) xor Codeword(1121) xor
                Codeword(1191) xor Codeword(1238) xor Codeword(1309) xor Codeword(1357) xor
                Codeword(1546) xor Codeword(1561) xor Codeword(1618) xor Codeword(1713) xor
                Codeword(1766) xor Codeword(1797) xor Codeword(1821) xor Codeword(1888);
 
     check217 <= Codeword(29) xor Codeword(75) xor Codeword(126) xor Codeword(201) xor
                Codeword(227) xor Codeword(329) xor Codeword(339) xor Codeword(414) xor
                Codeword(501) xor Codeword(524) xor Codeword(574) xor Codeword(627) xor
                Codeword(681) xor Codeword(747) xor Codeword(797) xor Codeword(860) xor
                Codeword(941) xor Codeword(961) xor Codeword(1044) xor Codeword(1078) xor
                Codeword(1122) xor Codeword(1204) xor Codeword(1266) xor Codeword(1299) xor
                Codeword(1332) xor Codeword(1362) xor Codeword(1389) xor Codeword(1542) xor
                Codeword(1606) xor Codeword(1628) xor Codeword(1667) xor Codeword(1776);
 
     check218 <= Codeword(28) xor Codeword(77) xor Codeword(154) xor Codeword(202) xor
                Codeword(261) xor Codeword(295) xor Codeword(375) xor Codeword(432) xor
                Codeword(483) xor Codeword(508) xor Codeword(616) xor Codeword(651) xor
                Codeword(693) xor Codeword(757) xor Codeword(811) xor Codeword(871) xor
                Codeword(915) xor Codeword(956) xor Codeword(1013) xor Codeword(1076) xor
                Codeword(1148) xor Codeword(1177) xor Codeword(1225) xor Codeword(1277) xor
                Codeword(1313) xor Codeword(1352) xor Codeword(1397) xor Codeword(1436) xor
                Codeword(1492) xor Codeword(1586) xor Codeword(1698) xor Codeword(1777);
 
     check219 <= Codeword(27) xor Codeword(101) xor Codeword(138) xor Codeword(182) xor
                Codeword(321) xor Codeword(354) xor Codeword(437) xor Codeword(489) xor
                Codeword(518) xor Codeword(573) xor Codeword(663) xor Codeword(702) xor
                Codeword(750) xor Codeword(804) xor Codeword(882) xor Codeword(929) xor
                Codeword(962) xor Codeword(1019) xor Codeword(1089) xor Codeword(1129) xor
                Codeword(1165) xor Codeword(1212) xor Codeword(1253) xor Codeword(1292) xor
                Codeword(1375) xor Codeword(1419) xor Codeword(1433) xor Codeword(1641) xor
                Codeword(1705) xor Codeword(1757) xor Codeword(1801) xor Codeword(1851);
 
     check220 <= Codeword(26) xor Codeword(83) xor Codeword(166) xor Codeword(173) xor
                Codeword(256) xor Codeword(305) xor Codeword(356) xor Codeword(447) xor
                Codeword(457) xor Codeword(525) xor Codeword(568) xor Codeword(659) xor
                Codeword(675) xor Codeword(754) xor Codeword(781) xor Codeword(855) xor
                Codeword(902) xor Codeword(950) xor Codeword(1004) xor Codeword(1082) xor
                Codeword(1140) xor Codeword(1179) xor Codeword(1233) xor Codeword(1282) xor
                Codeword(1289) xor Codeword(1381) xor Codeword(1420) xor Codeword(1475) xor
                Codeword(1594) xor Codeword(1629) xor Codeword(1656) xor Codeword(1778);
 
     check221 <= Codeword(25) xor Codeword(94) xor Codeword(156) xor Codeword(190) xor
                Codeword(268) xor Codeword(331) xor Codeword(342) xor Codeword(436) xor
                Codeword(455) xor Codeword(557) xor Codeword(604) xor Codeword(624) xor
                Codeword(689) xor Codeword(791) xor Codeword(843) xor Codeword(935) xor
                Codeword(976) xor Codeword(1111) xor Codeword(1149) xor Codeword(1302) xor
                Codeword(1334) xor Codeword(1365) xor Codeword(1396) xor Codeword(1590) xor
                Codeword(1660) xor Codeword(1704) xor Codeword(1727) xor Codeword(1876) xor
                Codeword(1882) xor Codeword(1935) xor Codeword(1940) xor Codeword(1946);
 
     check222 <= Codeword(24) xor Codeword(143) xor Codeword(241) xor Codeword(376) xor
                Codeword(430) xor Codeword(487) xor Codeword(611) xor Codeword(644) xor
                Codeword(777) xor Codeword(885) xor Codeword(904) xor Codeword(982) xor
                Codeword(1189) xor Codeword(1268) xor Codeword(1367) xor Codeword(1391) xor
                Codeword(1687) xor Codeword(1749) xor Codeword(1820) xor Codeword(1823) xor
                Codeword(1870) xor Codeword(1913) xor Codeword(1932) xor Codeword(1969) xor
                Codeword(1973) xor Codeword(1982) xor Codeword(2007) xor Codeword(2023) xor
                Codeword(2033) xor Codeword(2035) xor Codeword(2041) xor Codeword(2046);
 
     check223 <= Codeword(23) xor Codeword(76) xor Codeword(162) xor Codeword(224) xor
                Codeword(229) xor Codeword(309) xor Codeword(338) xor Codeword(411) xor
                Codeword(469) xor Codeword(543) xor Codeword(579) xor Codeword(645) xor
                Codeword(696) xor Codeword(788) xor Codeword(846) xor Codeword(917) xor
                Codeword(965) xor Codeword(1011) xor Codeword(1062) xor Codeword(1136) xor
                Codeword(1169) xor Codeword(1207) xor Codeword(1264) xor Codeword(1325) xor
                Codeword(1336) xor Codeword(1406) xor Codeword(1474) xor Codeword(1577) xor
                Codeword(1620) xor Codeword(1659) xor Codeword(1714) xor Codeword(1779);
 
     check224 <= Codeword(22) xor Codeword(90) xor Codeword(135) xor Codeword(193) xor
                Codeword(270) xor Codeword(328) xor Codeword(366) xor Codeword(419) xor
                Codeword(472) xor Codeword(520) xor Codeword(623) xor Codeword(718) xor
                Codeword(775) xor Codeword(779) xor Codeword(865) xor Codeword(914) xor
                Codeword(967) xor Codeword(1022) xor Codeword(1066) xor Codeword(1112) xor
                Codeword(1174) xor Codeword(1228) xor Codeword(1284) xor Codeword(1373) xor
                Codeword(1411) xor Codeword(1442) xor Codeword(1480) xor Codeword(1511) xor
                Codeword(1615) xor Codeword(1655) xor Codeword(1708) xor Codeword(1780);
 
     check225 <= Codeword(21) xor Codeword(61) xor Codeword(132) xor Codeword(188) xor
                Codeword(232) xor Codeword(301) xor Codeword(441) xor Codeword(458) xor
                Codeword(545) xor Codeword(609) xor Codeword(812) xor Codeword(873) xor
                Codeword(993) xor Codeword(1029) xor Codeword(1143) xor Codeword(1248) xor
                Codeword(1486) xor Codeword(1506) xor Codeword(1526) xor Codeword(1533) xor
                Codeword(1552) xor Codeword(1564) xor Codeword(1621) xor Codeword(1682) xor
                Codeword(1739) xor Codeword(1800) xor Codeword(1873) xor Codeword(1874) xor
                Codeword(1925) xor Codeword(1948) xor Codeword(1958) xor Codeword(1965);
 
     check226 <= Codeword(20) xor Codeword(148) xor Codeword(378) xor Codeword(488) xor
                Codeword(591) xor Codeword(758) xor Codeword(868) xor Codeword(897) xor
                Codeword(974) xor Codeword(1005) xor Codeword(1206) xor Codeword(1249) xor
                Codeword(1337) xor Codeword(1410) xor Codeword(1451) xor Codeword(1466) xor
                Codeword(1530) xor Codeword(1569) xor Codeword(1611) xor Codeword(1649) xor
                Codeword(1688) xor Codeword(1825) xor Codeword(1943) xor Codeword(1964) xor
                Codeword(1970) xor Codeword(1990) xor Codeword(1993) xor Codeword(2003) xor
                Codeword(2017) xor Codeword(2026) xor Codeword(2034) xor Codeword(2045);
 
     check227 <= Codeword(19) xor Codeword(63) xor Codeword(140) xor Codeword(178) xor
                Codeword(258) xor Codeword(314) xor Codeword(368) xor Codeword(417) xor
                Codeword(454) xor Codeword(555) xor Codeword(593) xor Codeword(634) xor
                Codeword(691) xor Codeword(746) xor Codeword(807) xor Codeword(874) xor
                Codeword(898) xor Codeword(986) xor Codeword(1018) xor Codeword(1075) xor
                Codeword(1123) xor Codeword(1198) xor Codeword(1227) xor Codeword(1322) xor
                Codeword(1366) xor Codeword(1404) xor Codeword(1445) xor Codeword(1575) xor
                Codeword(1595) xor Codeword(1631) xor Codeword(1706) xor Codeword(1781);
 
     check228 <= Codeword(18) xor Codeword(78) xor Codeword(114) xor Codeword(198) xor
                Codeword(253) xor Codeword(307) xor Codeword(398) xor Codeword(480) xor
                Codeword(580) xor Codeword(668) xor Codeword(713) xor Codeword(733) xor
                Codeword(819) xor Codeword(994) xor Codeword(1046) xor Codeword(1086) xor
                Codeword(1120) xor Codeword(1275) xor Codeword(1303) xor Codeword(1380) xor
                Codeword(1449) xor Codeword(1549) xor Codeword(1568) xor Codeword(1583) xor
                Codeword(1697) xor Codeword(1863) xor Codeword(1937) xor Codeword(1942) xor
                Codeword(1962) xor Codeword(1972) xor Codeword(1998) xor Codeword(2004);
 
     check229 <= Codeword(17) xor Codeword(74) xor Codeword(124) xor Codeword(259) xor
                Codeword(374) xor Codeword(466) xor Codeword(538) xor Codeword(610) xor
                Codeword(633) xor Codeword(832) xor Codeword(923) xor Codeword(966) xor
                Codeword(1236) xor Codeword(1288) xor Codeword(1354) xor Codeword(1495) xor
                Codeword(1515) xor Codeword(1556) xor Codeword(1625) xor Codeword(1798) xor
                Codeword(1842) xor Codeword(1878) xor Codeword(1959) xor Codeword(1976) xor
                Codeword(1981) xor Codeword(1988) xor Codeword(1991) xor Codeword(2001) xor
                Codeword(2010) xor Codeword(2019) xor Codeword(2031) xor Codeword(2043);
 
     check230 <= Codeword(16) xor Codeword(118) xor Codeword(176) xor Codeword(249) xor
                Codeword(293) xor Codeword(347) xor Codeword(442) xor Codeword(490) xor
                Codeword(539) xor Codeword(577) xor Codeword(690) xor Codeword(780) xor
                Codeword(838) xor Codeword(939) xor Codeword(981) xor Codeword(1048) xor
                Codeword(1069) xor Codeword(1161) xor Codeword(1218) xor Codeword(1240) xor
                Codeword(1300) xor Codeword(1519) xor Codeword(1600) xor Codeword(1626) xor
                Codeword(1700) xor Codeword(1809) xor Codeword(1819) xor Codeword(1831) xor
                Codeword(1949) xor Codeword(1978) xor Codeword(1996) xor Codeword(2005);
 
     check231 <= Codeword(15) xor Codeword(56) xor Codeword(209) xor Codeword(272) xor
                Codeword(287) xor Codeword(344) xor Codeword(418) xor Codeword(482) xor
                Codeword(516) xor Codeword(602) xor Codeword(666) xor Codeword(682) xor
                Codeword(722) xor Codeword(776) xor Codeword(821) xor Codeword(877) xor
                Codeword(943) xor Codeword(952) xor Codeword(1006) xor Codeword(1162) xor
                Codeword(1217) xor Codeword(1308) xor Codeword(1355) xor Codeword(1414) xor
                Codeword(1470) xor Codeword(1507) xor Codeword(1525) xor Codeword(1578) xor
                Codeword(1647) xor Codeword(1672) xor Codeword(1804) xor Codeword(1852);
 
     check232 <= Codeword(14) xor Codeword(57) xor Codeword(212) xor Codeword(278) xor
                Codeword(291) xor Codeword(359) xor Codeword(439) xor Codeword(470) xor
                Codeword(509) xor Codeword(700) xor Codeword(783) xor Codeword(879) xor
                Codeword(989) xor Codeword(1097) xor Codeword(1138) xor Codeword(1166) xor
                Codeword(1213) xor Codeword(1368) xor Codeword(1476) xor Codeword(1502) xor
                Codeword(1504) xor Codeword(1573) xor Codeword(1664) xor Codeword(1746) xor
                Codeword(1756) xor Codeword(1760) xor Codeword(1864) xor Codeword(1910) xor
                Codeword(1920) xor Codeword(1951) xor Codeword(1952) xor Codeword(1966);
 
     check233 <= Codeword(13) xor Codeword(92) xor Codeword(149) xor Codeword(263) xor
                Codeword(352) xor Codeword(486) xor Codeword(612) xor Codeword(640) xor
                Codeword(723) xor Codeword(850) xor Codeword(954) xor Codeword(1195) xor
                Codeword(1276) xor Codeword(1324) xor Codeword(1364) xor Codeword(1494) xor
                Codeword(1537) xor Codeword(1640) xor Codeword(1711) xor Codeword(1832) xor
                Codeword(1834) xor Codeword(1892) xor Codeword(1909) xor Codeword(1960) xor
                Codeword(1983) xor Codeword(1995) xor Codeword(2008) xor Codeword(2013) xor
                Codeword(2020) xor Codeword(2028) xor Codeword(2039) xor Codeword(2047);
 
     check234 <= Codeword(12) xor Codeword(84) xor Codeword(131) xor Codeword(177) xor
                Codeword(265) xor Codeword(315) xor Codeword(386) xor Codeword(394) xor
                Codeword(463) xor Codeword(528) xor Codeword(603) xor Codeword(638) xor
                Codeword(768) xor Codeword(809) xor Codeword(886) xor Codeword(937) xor
                Codeword(968) xor Codeword(1041) xor Codeword(1147) xor Codeword(1202) xor
                Codeword(1272) xor Codeword(1310) xor Codeword(1383) xor Codeword(1452) xor
                Codeword(1468) xor Codeword(1478) xor Codeword(1498) xor Codeword(1662) xor
                Codeword(1753) xor Codeword(1791) xor Codeword(1808) xor Codeword(1853);
 
     check235 <= Codeword(100) xor Codeword(144) xor Codeword(196) xor Codeword(235) xor
                Codeword(336) xor Codeword(420) xor Codeword(460) xor Codeword(619) xor
                Codeword(704) xor Codeword(736) xor Codeword(805) xor Codeword(842) xor
                Codeword(921) xor Codeword(964) xor Codeword(1042) xor Codeword(1152) xor
                Codeword(1170) xor Codeword(1327) xor Codeword(1349) xor Codeword(1416) xor
                Codeword(1427) xor Codeword(1497) xor Codeword(1523) xor Codeword(1558) xor
                Codeword(1799) xor Codeword(1818) xor Codeword(1826) xor Codeword(1830) xor
                Codeword(1837) xor Codeword(1838) xor Codeword(1867) xor Codeword(1889);
 
     check236 <= Codeword(11) xor Codeword(104) xor Codeword(155) xor Codeword(221) xor
                Codeword(271) xor Codeword(310) xor Codeword(390) xor Codeword(410) xor
                Codeword(475) xor Codeword(527) xor Codeword(608) xor Codeword(653) xor
                Codeword(698) xor Codeword(742) xor Codeword(810) xor Codeword(851) xor
                Codeword(927) xor Codeword(984) xor Codeword(1020) xor Codeword(1083) xor
                Codeword(1244) xor Codeword(1278) xor Codeword(1293) xor Codeword(1350) xor
                Codeword(1393) xor Codeword(1429) xor Codeword(1514) xor Codeword(1517) xor
                Codeword(1592) xor Codeword(1636) xor Codeword(1669) xor Codeword(1782);
 
     check237 <= Codeword(10) xor Codeword(110) xor Codeword(125) xor Codeword(228) xor
                Codeword(322) xor Codeword(334) xor Codeword(399) xor Codeword(467) xor
                Codeword(522) xor Codeword(584) xor Codeword(654) xor Codeword(680) xor
                Codeword(726) xor Codeword(800) xor Codeword(878) xor Codeword(893) xor
                Codeword(947) xor Codeword(1012) xor Codeword(1088) xor Codeword(1151) xor
                Codeword(1200) xor Codeword(1242) xor Codeword(1301) xor Codeword(1382) xor
                Codeword(1413) xor Codeword(1444) xor Codeword(1574) xor Codeword(1612) xor
                Codeword(1650) xor Codeword(1695) xor Codeword(1789) xor Codeword(1854);
 
     check238 <= Codeword(9) xor Codeword(103) xor Codeword(113) xor Codeword(179) xor
                Codeword(236) xor Codeword(294) xor Codeword(383) xor Codeword(416) xor
                Codeword(498) xor Codeword(507) xor Codeword(582) xor Codeword(641) xor
                Codeword(687) xor Codeword(728) xor Codeword(824) xor Codeword(837) xor
                Codeword(891) xor Codeword(948) xor Codeword(1028) xor Codeword(1059) xor
                Codeword(1079) xor Codeword(1145) xor Codeword(1182) xor Codeword(1297) xor
                Codeword(1374) xor Codeword(1469) xor Codeword(1521) xor Codeword(1547) xor
                Codeword(1593) xor Codeword(1643) xor Codeword(1715) xor Codeword(1783);
 
     check239 <= Codeword(8) xor Codeword(98) xor Codeword(158) xor Codeword(223) xor
                Codeword(264) xor Codeword(284) xor Codeword(360) xor Codeword(392) xor
                Codeword(452) xor Codeword(513) xor Codeword(596) xor Codeword(620) xor
                Codeword(710) xor Codeword(752) xor Codeword(829) xor Codeword(866) xor
                Codeword(926) xor Codeword(983) xor Codeword(1032) xor Codeword(1099) xor
                Codeword(1127) xor Codeword(1185) xor Codeword(1424) xor Codeword(1572) xor
                Codeword(1587) xor Codeword(1717) xor Codeword(1794) xor Codeword(1811) xor
                Codeword(1814) xor Codeword(1817) xor Codeword(1866) xor Codeword(1890);
 
     check240 <= Codeword(7) xor Codeword(81) xor Codeword(116) xor Codeword(210) xor
                Codeword(277) xor Codeword(324) xor Codeword(343) xor Codeword(444) xor
                Codeword(502) xor Codeword(534) xor Codeword(589) xor Codeword(637) xor
                Codeword(708) xor Codeword(734) xor Codeword(814) xor Codeword(845) xor
                Codeword(907) xor Codeword(975) xor Codeword(1105) xor Codeword(1113) xor
                Codeword(1134) xor Codeword(1171) xor Codeword(1259) xor Codeword(1339) xor
                Codeword(1394) xor Codeword(1437) xor Codeword(1505) xor Codeword(1605) xor
                Codeword(1686) xor Codeword(1703) xor Codeword(1806) xor Codeword(1855);
 
     check241 <= Codeword(6) xor Codeword(88) xor Codeword(175) xor Codeword(250) xor
                Codeword(285) xor Codeword(355) xor Codeword(403) xor Codeword(449) xor
                Codeword(532) xor Codeword(565) xor Codeword(685) xor Codeword(745) xor
                Codeword(816) xor Codeword(992) xor Codeword(1031) xor Codeword(1090) xor
                Codeword(1157) xor Codeword(1168) xor Codeword(1201) xor Codeword(1245) xor
                Codeword(1388) xor Codeword(1463) xor Codeword(1536) xor Codeword(1548) xor
                Codeword(1624) xor Codeword(1690) xor Codeword(1802) xor Codeword(1891) xor
                Codeword(1893) xor Codeword(1901) xor Codeword(1941) xor Codeword(1947);
 
     check242 <= Codeword(5) xor Codeword(108) xor Codeword(146) xor Codeword(203) xor
                Codeword(231) xor Codeword(303) xor Codeword(367) xor Codeword(396) xor
                Codeword(495) xor Codeword(511) xor Codeword(575) xor Codeword(650) xor
                Codeword(720) xor Codeword(753) xor Codeword(786) xor Codeword(880) xor
                Codeword(894) xor Codeword(997) xor Codeword(1003) xor Codeword(1026) xor
                Codeword(1092) xor Codeword(1155) xor Codeword(1319) xor Codeword(1338) xor
                Codeword(1471) xor Codeword(1522) xor Codeword(1596) xor Codeword(1638) xor
                Codeword(1666) xor Codeword(1696) xor Codeword(1786) xor Codeword(1856);
 
     check243 <= Codeword(4) xor Codeword(106) xor Codeword(141) xor Codeword(200) xor
                Codeword(252) xor Codeword(312) xor Codeword(337) xor Codeword(427) xor
                Codeword(476) xor Codeword(548) xor Codeword(569) xor Codeword(670) xor
                Codeword(727) xor Codeword(822) xor Codeword(1009) xor Codeword(1064) xor
                Codeword(1132) xor Codeword(1281) xor Codeword(1335) xor Codeword(1439) xor
                Codeword(1503) xor Codeword(1598) xor Codeword(1675) xor Codeword(1744) xor
                Codeword(1764) xor Codeword(1816) xor Codeword(1872) xor Codeword(1904) xor
                Codeword(1927) xor Codeword(1950) xor Codeword(1968) xor Codeword(1971);
 
     check244 <= Codeword(147) xor Codeword(266) xor Codeword(385) xor Codeword(459) xor
                Codeword(551) xor Codeword(572) xor Codeword(665) xor Codeword(741) xor
                Codeword(840) xor Codeword(890) xor Codeword(996) xor Codeword(1016) xor
                Codeword(1178) xor Codeword(1269) xor Codeword(1305) xor Codeword(1371) xor
                Codeword(1421) xor Codeword(1482) xor Codeword(1554) xor Codeword(1609) xor
                Codeword(1716) xor Codeword(1807) xor Codeword(1980) xor Codeword(1986) xor
                Codeword(1987) xor Codeword(1992) xor Codeword(1999) xor Codeword(2011) xor
                Codeword(2014) xor Codeword(2024) xor Codeword(2030) xor Codeword(2038);
 
     check245 <= Codeword(3) xor Codeword(66) xor Codeword(136) xor Codeword(207) xor
                Codeword(262) xor Codeword(313) xor Codeword(370) xor Codeword(431) xor
                Codeword(471) xor Codeword(535) xor Codeword(562) xor Codeword(686) xor
                Codeword(769) xor Codeword(787) xor Codeword(862) xor Codeword(918) xor
                Codeword(991) xor Codeword(1037) xor Codeword(1109) xor Codeword(1115) xor
                Codeword(1203) xor Codeword(1220) xor Codeword(1254) xor Codeword(1378) xor
                Codeword(1418) xor Codeword(1467) xor Codeword(1528) xor Codeword(1603) xor
                Codeword(1637) xor Codeword(1653) xor Codeword(1759) xor Codeword(1857);
 
     check246 <= Codeword(2) xor Codeword(69) xor Codeword(161) xor Codeword(185) xor
                Codeword(226) xor Codeword(302) xor Codeword(388) xor Codeword(435) xor
                Codeword(481) xor Codeword(512) xor Codeword(597) xor Codeword(618) xor
                Codeword(707) xor Codeword(748) xor Codeword(815) xor Codeword(863) xor
                Codeword(903) xor Codeword(972) xor Codeword(1035) xor Codeword(1065) xor
                Codeword(1158) xor Codeword(1194) xor Codeword(1222) xor Codeword(1311) xor
                Codeword(1345) xor Codeword(1384) xor Codeword(1524) xor Codeword(1540) xor
                Codeword(1630) xor Codeword(1661) xor Codeword(1709) xor Codeword(1784);
 
     check247 <= Codeword(1) xor Codeword(109) xor Codeword(168) xor Codeword(194) xor
                Codeword(247) xor Codeword(327) xor Codeword(349) xor Codeword(424) xor
                Codeword(453) xor Codeword(531) xor Codeword(581) xor Codeword(646) xor
                Codeword(677) xor Codeword(771) xor Codeword(828) xor Codeword(839) xor
                Codeword(928) xor Codeword(980) xor Codeword(1014) xor Codeword(1091) xor
                Codeword(1133) xor Codeword(1183) xor Codeword(1271) xor Codeword(1323) xor
                Codeword(1333) xor Codeword(1343) xor Codeword(1447) xor Codeword(1483) xor
                Codeword(1646) xor Codeword(1699) xor Codeword(1755) xor Codeword(1858);
 
     check248 <= Codeword(0) xor Codeword(87) xor Codeword(151) xor Codeword(189) xor
                Codeword(248) xor Codeword(280) xor Codeword(357) xor Codeword(404) xor
                Codeword(497) xor Codeword(559) xor Codeword(592) xor Codeword(643) xor
                Codeword(717) xor Codeword(729) xor Codeword(801) xor Codeword(831) xor
                Codeword(920) xor Codeword(1002) xor Codeword(1051) xor Codeword(1104) xor
                Codeword(1154) xor Codeword(1199) xor Codeword(1257) xor Codeword(1279) xor
                Codeword(1377) xor Codeword(1401) xor Codeword(1431) xor Codeword(1490) xor
                Codeword(1529) xor Codeword(1597) xor Codeword(1658) xor Codeword(1785);
 
     check249 <= Codeword(152) xor Codeword(192) xor Codeword(225) xor Codeword(317) xor
                Codeword(353) xor Codeword(443) xor Codeword(544) xor Codeword(657) xor
                Codeword(688) xor Codeword(725) xor Codeword(782) xor Codeword(849) xor
                Codeword(908) xor Codeword(1000) xor Codeword(1054) xor Codeword(1124) xor
                Codeword(1175) xor Codeword(1304) xor Codeword(1390) xor Codeword(1462) xor
                Codeword(1520) xor Codeword(1557) xor Codeword(1648) xor Codeword(1723) xor
                Codeword(1735) xor Codeword(1736) xor Codeword(1741) xor Codeword(1751) xor
                Codeword(1822) xor Codeword(1840) xor Codeword(1883) xor Codeword(1911);
 
     check250 <= Codeword(79) xor Codeword(120) xor Codeword(184) xor Codeword(319) xor
                Codeword(358) xor Codeword(400) xor Codeword(500) xor Codeword(514) xor
                Codeword(576) xor Codeword(652) xor Codeword(679) xor Codeword(744) xor
                Codeword(803) xor Codeword(854) xor Codeword(925) xor Codeword(978) xor
                Codeword(1038) xor Codeword(1173) xor Codeword(1250) xor Codeword(1318) xor
                Codeword(1360) xor Codeword(1405) xor Codeword(1448) xor Codeword(1489) xor
                Codeword(1508) xor Codeword(1512) xor Codeword(1560) xor Codeword(1588) xor
                Codeword(1676) xor Codeword(1762) xor Codeword(1928) xor Codeword(1933);
 
     check251 <= Codeword(62) xor Codeword(159) xor Codeword(215) xor Codeword(289) xor
                Codeword(348) xor Codeword(409) xor Codeword(464) xor Codeword(506) xor
                Codeword(564) xor Codeword(626) xor Codeword(721) xor Codeword(765) xor
                Codeword(817) xor Codeword(899) xor Codeword(957) xor Codeword(1015) xor
                Codeword(1081) xor Codeword(1135) xor Codeword(1187) xor Codeword(1221) xor
                Codeword(1247) xor Codeword(1294) xor Codeword(1346) xor Codeword(1409) xor
                Codeword(1477) xor Codeword(1501) xor Codeword(1570) xor Codeword(1644) xor
                Codeword(1665) xor Codeword(1722) xor Codeword(1793) xor Codeword(1859);
 
     check252 <= Codeword(89) xor Codeword(112) xor Codeword(199) xor Codeword(239) xor
                Codeword(325) xor Codeword(373) xor Codeword(438) xor Codeword(473) xor
                Codeword(549) xor Codeword(605) xor Codeword(635) xor Codeword(684) xor
                Codeword(766) xor Codeword(813) xor Codeword(853) xor Codeword(896) xor
                Codeword(960) xor Codeword(1034) xor Codeword(1093) xor Codeword(1126) xor
                Codeword(1180) xor Codeword(1262) xor Codeword(1326) xor Codeword(1398) xor
                Codeword(1563) xor Codeword(1589) xor Codeword(1671) xor Codeword(1721) xor
                Codeword(1731) xor Codeword(1742) xor Codeword(1805) xor Codeword(1860);
 
     check253 <= Codeword(80) xor Codeword(121) xor Codeword(211) xor Codeword(279) xor
                Codeword(283) xor Codeword(380) xor Codeword(426) xor Codeword(468) xor
                Codeword(510) xor Codeword(567) xor Codeword(629) xor Codeword(714) xor
                Codeword(743) xor Codeword(778) xor Codeword(847) xor Codeword(912) xor
                Codeword(944) xor Codeword(1007) xor Codeword(1060) xor Codeword(1114) xor
                Codeword(1211) xor Codeword(1255) xor Codeword(1296) xor Codeword(1342) xor
                Codeword(1541) xor Codeword(1567) xor Codeword(1599) xor Codeword(1635) xor
                Codeword(1681) xor Codeword(1719) xor Codeword(1768) xor Codeword(1861);
 
     check254 <= Codeword(67) xor Codeword(222) xor Codeword(238) xor Codeword(290) xor
                Codeword(362) xor Codeword(412) xor Codeword(474) xor Codeword(540) xor
                Codeword(586) xor Codeword(632) xor Codeword(712) xor Codeword(735) xor
                Codeword(798) xor Codeword(884) xor Codeword(905) xor Codeword(979) xor
                Codeword(1047) xor Codeword(1107) xor Codeword(1131) xor Codeword(1232) xor
                Codeword(1306) xor Codeword(1369) xor Codeword(1417) xor Codeword(1443) xor
                Codeword(1456) xor Codeword(1493) xor Codeword(1516) xor Codeword(1720) xor
                Codeword(1733) xor Codeword(1754) xor Codeword(1923) xor Codeword(1926);
 
     check255 <= Codeword(52) xor Codeword(86) xor Codeword(167) xor Codeword(195) xor
                Codeword(233) xor Codeword(318) xor Codeword(364) xor Codeword(429) xor
                Codeword(537) xor Codeword(594) xor Codeword(672) xor Codeword(751) xor
                Codeword(799) xor Codeword(934) xor Codeword(1017) xor Codeword(1077) xor
                Codeword(1110) xor Codeword(1163) xor Codeword(1214) xor Codeword(1432) xor
                Codeword(1465) xor Codeword(1538) xor Codeword(1691) xor Codeword(1787) xor
                Codeword(1836) xor Codeword(1879) xor Codeword(1897) xor Codeword(1906) xor
                Codeword(1929) xor Codeword(1936) xor Codeword(1961) xor Codeword(1979);
 
     check256 <= Codeword(53) xor Codeword(106) xor Codeword(127) xor Codeword(242) xor
                Codeword(296) xor Codeword(339) xor Codeword(455) xor Codeword(532) xor
                Codeword(638) xor Codeword(708) xor Codeword(760) xor Codeword(793) xor
                Codeword(891) xor Codeword(1000) xor Codeword(1035) xor Codeword(1071) xor
                Codeword(1155) xor Codeword(1242) xor Codeword(1285) xor Codeword(1343) xor
                Codeword(1414) xor Codeword(1454) xor Codeword(1517) xor Codeword(1747) xor
                Codeword(1780) xor Codeword(1846) xor Codeword(1929) xor Codeword(1959) xor
                Codeword(1962) xor Codeword(1990) xor Codeword(1995) xor Codeword(1997);
 
     check257 <= Codeword(51) xor Codeword(85) xor Codeword(166) xor Codeword(194) xor
                Codeword(232) xor Codeword(317) xor Codeword(363) xor Codeword(428) xor
                Codeword(463) xor Codeword(536) xor Codeword(593) xor Codeword(624) xor
                Codeword(671) xor Codeword(750) xor Codeword(798) xor Codeword(835) xor
                Codeword(933) xor Codeword(999) xor Codeword(1016) xor Codeword(1076) xor
                Codeword(1108) xor Codeword(1162) xor Codeword(1213) xor Codeword(1240) xor
                Codeword(1303) xor Codeword(1354) xor Codeword(1431) xor Codeword(1464) xor
                Codeword(1484) xor Codeword(1652) xor Codeword(1690) xor Codeword(1786);
 
     check258 <= Codeword(50) xor Codeword(57) xor Codeword(331) xor Codeword(553) xor
                Codeword(589) xor Codeword(657) xor Codeword(718) xor Codeword(755) xor
                Codeword(829) xor Codeword(857) xor Codeword(943) xor Codeword(968) xor
                Codeword(1077) xor Codeword(1159) xor Codeword(1215) xor Codeword(1222) xor
                Codeword(1320) xor Codeword(1378) xor Codeword(1547) xor Codeword(1574) xor
                Codeword(1632) xor Codeword(1682) xor Codeword(1770) xor Codeword(1778) xor
                Codeword(1801) xor Codeword(1834) xor Codeword(1884) xor Codeword(1901) xor
                Codeword(1921) xor Codeword(1922) xor Codeword(1945) xor Codeword(1954);
 
     check259 <= Codeword(54) xor Codeword(114) xor Codeword(274) xor Codeword(303) xor
                Codeword(370) xor Codeword(491) xor Codeword(545) xor Codeword(594) xor
                Codeword(641) xor Codeword(694) xor Codeword(822) xor Codeword(856) xor
                Codeword(937) xor Codeword(952) xor Codeword(1051) xor Codeword(1105) xor
                Codeword(1117) xor Codeword(1207) xor Codeword(1218) xor Codeword(1238) xor
                Codeword(1289) xor Codeword(1499) xor Codeword(1584) xor Codeword(1615) xor
                Codeword(1728) xor Codeword(1735) xor Codeword(1738) xor Codeword(1833) xor
                Codeword(1844) xor Codeword(1970) xor Codeword(1981) xor Codeword(1986);
 
     check260 <= Codeword(49) xor Codeword(71) xor Codeword(138) xor Codeword(186) xor
                Codeword(243) xor Codeword(383) xor Codeword(396) xor Codeword(584) xor
                Codeword(754) xor Codeword(833) xor Codeword(941) xor Codeword(980) xor
                Codeword(1013) xor Codeword(1187) xor Codeword(1228) xor Codeword(1290) xor
                Codeword(1399) xor Codeword(1437) xor Codeword(1463) xor Codeword(1618) xor
                Codeword(1718) xor Codeword(1765) xor Codeword(1771) xor Codeword(1822) xor
                Codeword(1857) xor Codeword(1943) xor Codeword(1963) xor Codeword(1988) xor
                Codeword(2015) xor Codeword(2020) xor Codeword(2023) xor Codeword(2030);
 
     check261 <= Codeword(48) xor Codeword(63) xor Codeword(152) xor Codeword(204) xor
                Codeword(305) xor Codeword(333) xor Codeword(401) xor Codeword(477) xor
                Codeword(528) xor Codeword(607) xor Codeword(698) xor Codeword(777) xor
                Codeword(789) xor Codeword(868) xor Codeword(970) xor Codeword(1042) xor
                Codeword(1062) xor Codeword(1141) xor Codeword(1171) xor Codeword(1262) xor
                Codeword(1319) xor Codeword(1375) xor Codeword(1493) xor Codeword(1549) xor
                Codeword(1570) xor Codeword(1603) xor Codeword(1672) xor Codeword(1704) xor
                Codeword(1761) xor Codeword(1842) xor Codeword(1874) xor Codeword(1891);
 
     check262 <= Codeword(47) xor Codeword(95) xor Codeword(149) xor Codeword(212) xor
                Codeword(319) xor Codeword(362) xor Codeword(392) xor Codeword(503) xor
                Codeword(522) xor Codeword(613) xor Codeword(635) xor Codeword(702) xor
                Codeword(731) xor Codeword(830) xor Codeword(871) xor Codeword(912) xor
                Codeword(957) xor Codeword(1039) xor Codeword(1067) xor Codeword(1152) xor
                Codeword(1183) xor Codeword(1245) xor Codeword(1311) xor Codeword(1350) xor
                Codeword(1402) xor Codeword(1480) xor Codeword(1500) xor Codeword(1559) xor
                Codeword(1633) xor Codeword(1700) xor Codeword(1807) xor Codeword(1862);
 
     check263 <= Codeword(46) xor Codeword(104) xor Codeword(169) xor Codeword(207) xor
                Codeword(253) xor Codeword(315) xor Codeword(378) xor Codeword(414) xor
                Codeword(525) xor Codeword(598) xor Codeword(691) xor Codeword(738) xor
                Codeword(788) xor Codeword(858) xor Codeword(894) xor Codeword(976) xor
                Codeword(1056) xor Codeword(1145) xor Codeword(1257) xor Codeword(1347) xor
                Codeword(1492) xor Codeword(1509) xor Codeword(1526) xor Codeword(1554) xor
                Codeword(1576) xor Codeword(1673) xor Codeword(1743) xor Codeword(1840) xor
                Codeword(1841) xor Codeword(1905) xor Codeword(1971) xor Codeword(1978);
 
     check264 <= Codeword(45) xor Codeword(98) xor Codeword(132) xor Codeword(213) xor
                Codeword(256) xor Codeword(281) xor Codeword(349) xor Codeword(421) xor
                Codeword(495) xor Codeword(600) xor Codeword(666) xor Codeword(672) xor
                Codeword(761) xor Codeword(783) xor Codeword(834) xor Codeword(908) xor
                Codeword(948) xor Codeword(1048) xor Codeword(1066) xor Codeword(1149) xor
                Codeword(1269) xor Codeword(1279) xor Codeword(1362) xor Codeword(1516) xor
                Codeword(1531) xor Codeword(1561) xor Codeword(1607) xor Codeword(1693) xor
                Codeword(1753) xor Codeword(1802) xor Codeword(1806) xor Codeword(1863);
 
     check265 <= Codeword(44) xor Codeword(133) xor Codeword(203) xor Codeword(244) xor
                Codeword(386) xor Codeword(405) xor Codeword(504) xor Codeword(627) xor
                Codeword(759) xor Codeword(855) xor Codeword(918) xor Codeword(945) xor
                Codeword(1023) xor Codeword(1209) xor Codeword(1355) xor Codeword(1385) xor
                Codeword(1445) xor Codeword(1486) xor Codeword(1532) xor Codeword(1612) xor
                Codeword(1757) xor Codeword(1845) xor Codeword(1858) xor Codeword(1888) xor
                Codeword(1906) xor Codeword(1915) xor Codeword(1992) xor Codeword(1993) xor
                Codeword(2028) xor Codeword(2032) xor Codeword(2043) xor Codeword(2046);
 
     check266 <= Codeword(43) xor Codeword(168) xor Codeword(173) xor Codeword(273) xor
                Codeword(300) xor Codeword(535) xor Codeword(605) xor Codeword(647) xor
                Codeword(721) xor Codeword(880) xor Codeword(888) xor Codeword(962) xor
                Codeword(1032) xor Codeword(1095) xor Codeword(1118) xor Codeword(1195) xor
                Codeword(1230) xor Codeword(1429) xor Codeword(1478) xor Codeword(1530) xor
                Codeword(1534) xor Codeword(1539) xor Codeword(1635) xor Codeword(1725) xor
                Codeword(1815) xor Codeword(1824) xor Codeword(1827) xor Codeword(1898) xor
                Codeword(1908) xor Codeword(1965) xor Codeword(1996) xor Codeword(2006);
 
     check267 <= Codeword(42) xor Codeword(72) xor Codeword(159) xor Codeword(180) xor
                Codeword(241) xor Codeword(280) xor Codeword(364) xor Codeword(432) xor
                Codeword(490) xor Codeword(549) xor Codeword(562) xor Codeword(654) xor
                Codeword(677) xor Codeword(794) xor Codeword(866) xor Codeword(932) xor
                Codeword(954) xor Codeword(1026) xor Codeword(1101) xor Codeword(1158) xor
                Codeword(1212) xor Codeword(1272) xor Codeword(1327) xor Codeword(1339) xor
                Codeword(1390) xor Codeword(1421) xor Codeword(1601) xor Codeword(1628) xor
                Codeword(1677) xor Codeword(1692) xor Codeword(1724) xor Codeword(1864);
 
     check268 <= Codeword(41) xor Codeword(109) xor Codeword(118) xor Codeword(216) xor
                Codeword(266) xor Codeword(325) xor Codeword(360) xor Codeword(412) xor
                Codeword(464) xor Codeword(559) xor Codeword(570) xor Codeword(652) xor
                Codeword(705) xor Codeword(775) xor Codeword(792) xor Codeword(921) xor
                Codeword(987) xor Codeword(1029) xor Codeword(1072) xor Codeword(1114) xor
                Codeword(1176) xor Codeword(1233) xor Codeword(1309) xor Codeword(1335) xor
                Codeword(1391) xor Codeword(1430) xor Codeword(1449) xor Codeword(1459) xor
                Codeword(1616) xor Codeword(1678) xor Codeword(1711) xor Codeword(1787);
 
     check269 <= Codeword(67) xor Codeword(122) xor Codeword(218) xor Codeword(250) xor
                Codeword(287) xor Codeword(381) xor Codeword(424) xor Codeword(498) xor
                Codeword(529) xor Codeword(599) xor Codeword(655) xor Codeword(693) xor
                Codeword(762) xor Codeword(825) xor Codeword(882) xor Codeword(935) xor
                Codeword(997) xor Codeword(1070) xor Codeword(1124) xor Codeword(1185) xor
                Codeword(1251) xor Codeword(1315) xor Codeword(1337) xor Codeword(1384) xor
                Codeword(1395) xor Codeword(1444) xor Codeword(1580) xor Codeword(1631) xor
                Codeword(1656) xor Codeword(1739) xor Codeword(1810) xor Codeword(1892);
 
     check270 <= Codeword(40) xor Codeword(79) xor Codeword(170) xor Codeword(190) xor
                Codeword(275) xor Codeword(292) xor Codeword(344) xor Codeword(433) xor
                Codeword(466) xor Codeword(518) xor Codeword(612) xor Codeword(646) xor
                Codeword(680) xor Codeword(737) xor Codeword(805) xor Codeword(869) xor
                Codeword(900) xor Codeword(991) xor Codeword(1057) xor Codeword(1100) xor
                Codeword(1153) xor Codeword(1180) xor Codeword(1259) xor Codeword(1277) xor
                Codeword(1383) xor Codeword(1442) xor Codeword(1542) xor Codeword(1579) xor
                Codeword(1609) xor Codeword(1683) xor Codeword(1707) xor Codeword(1788);
 
     check271 <= Codeword(39) xor Codeword(105) xor Codeword(171) xor Codeword(268) xor
                Codeword(332) xor Codeword(345) xor Codeword(406) xor Codeword(478) xor
                Codeword(507) xor Codeword(586) xor Codeword(696) xor Codeword(758) xor
                Codeword(807) xor Codeword(832) xor Codeword(994) xor Codeword(1038) xor
                Codeword(1083) xor Codeword(1140) xor Codeword(1255) xor Codeword(1330) xor
                Codeword(1363) xor Codeword(1472) xor Codeword(1544) xor Codeword(1606) xor
                Codeword(1608) xor Codeword(1803) xor Codeword(1849) xor Codeword(1852) xor
                Codeword(1895) xor Codeword(1911) xor Codeword(1941) xor Codeword(1948);
 
     check272 <= Codeword(38) xor Codeword(94) xor Codeword(116) xor Codeword(184) xor
                Codeword(254) xor Codeword(291) xor Codeword(380) xor Codeword(420) xor
                Codeword(476) xor Codeword(520) xor Codeword(565) xor Codeword(621) xor
                Codeword(715) xor Codeword(729) xor Codeword(795) xor Codeword(863) xor
                Codeword(905) xor Codeword(984) xor Codeword(1052) xor Codeword(1086) xor
                Codeword(1127) xor Codeword(1175) xor Codeword(1260) xor Codeword(1313) xor
                Codeword(1346) xor Codeword(1406) xor Codeword(1433) xor Codeword(1455) xor
                Codeword(1621) xor Codeword(1657) xor Codeword(1706) xor Codeword(1789);
 
     check273 <= Codeword(37) xor Codeword(81) xor Codeword(156) xor Codeword(272) xor
                Codeword(285) xor Codeword(371) xor Codeword(493) xor Codeword(541) xor
                Codeword(659) xor Codeword(670) xor Codeword(769) xor Codeword(826) xor
                Codeword(860) xor Codeword(910) xor Codeword(963) xor Codeword(1007) xor
                Codeword(1073) xor Codeword(1143) xor Codeword(1198) xor Codeword(1250) xor
                Codeword(1297) xor Codeword(1358) xor Codeword(1453) xor Codeword(1550) xor
                Codeword(1726) xor Codeword(1736) xor Codeword(1817) xor Codeword(1910) xor
                Codeword(1918) xor Codeword(1984) xor Codeword(2031) xor Codeword(2042);
 
     check274 <= Codeword(36) xor Codeword(164) xor Codeword(217) xor Codeword(248) xor
                Codeword(390) xor Codeword(427) xor Codeword(460) xor Codeword(551) xor
                Codeword(601) xor Codeword(661) xor Codeword(739) xor Codeword(874) xor
                Codeword(899) xor Codeword(944) xor Codeword(1033) xor Codeword(1204) xor
                Codeword(1275) xor Codeword(1282) xor Codeword(1300) xor Codeword(1369) xor
                Codeword(1398) xor Codeword(1564) xor Codeword(1581) xor Codeword(1641) xor
                Codeword(1650) xor Codeword(1709) xor Codeword(1985) xor Codeword(2002) xor
                Codeword(2017) xor Codeword(2019) xor Codeword(2029) xor Codeword(2033);
 
     check275 <= Codeword(35) xor Codeword(59) xor Codeword(128) xor Codeword(179) xor
                Codeword(329) xor Codeword(394) xor Codeword(461) xor Codeword(546) xor
                Codeword(597) xor Codeword(817) xor Codeword(923) xor Codeword(958) xor
                Codeword(1022) xor Codeword(1069) xor Codeword(1113) xor Codeword(1115) xor
                Codeword(1189) xor Codeword(1225) xor Codeword(1286) xor Codeword(1340) xor
                Codeword(1407) xor Codeword(1440) xor Codeword(1458) xor Codeword(1490) xor
                Codeword(1668) xor Codeword(1813) xor Codeword(1825) xor Codeword(1848) xor
                Codeword(1851) xor Codeword(1873) xor Codeword(1875) xor Codeword(1893);
 
     check276 <= Codeword(34) xor Codeword(69) xor Codeword(126) xor Codeword(205) xor
                Codeword(259) xor Codeword(297) xor Codeword(407) xor Codeword(492) xor
                Codeword(552) xor Codeword(615) xor Codeword(667) xor Codeword(714) xor
                Codeword(773) xor Codeword(801) xor Codeword(843) xor Codeword(929) xor
                Codeword(969) xor Codeword(1009) xor Codeword(1093) xor Codeword(1166) xor
                Codeword(1191) xor Codeword(1264) xor Codeword(1314) xor Codeword(1456) xor
                Codeword(1496) xor Codeword(1533) xor Codeword(1543) xor Codeword(1578) xor
                Codeword(1644) xor Codeword(1653) xor Codeword(1688) xor Codeword(1790);
 
     check277 <= Codeword(33) xor Codeword(64) xor Codeword(162) xor Codeword(185) xor
                Codeword(252) xor Codeword(295) xor Codeword(334) xor Codeword(391) xor
                Codeword(404) xor Codeword(484) xor Codeword(540) xor Codeword(582) xor
                Codeword(682) xor Codeword(736) xor Codeword(854) xor Codeword(914) xor
                Codeword(998) xor Codeword(1116) xor Codeword(1266) xor Codeword(1371) xor
                Codeword(1394) xor Codeword(1565) xor Codeword(1599) xor Codeword(1669) xor
                Codeword(1751) xor Codeword(1758) xor Codeword(1808) xor Codeword(1936) xor
                Codeword(1951) xor Codeword(2000) xor Codeword(2004) xor Codeword(2010);
 
     check278 <= Codeword(32) xor Codeword(70) xor Codeword(141) xor Codeword(229) xor
                Codeword(328) xor Codeword(388) xor Codeword(423) xor Codeword(502) xor
                Codeword(509) xor Codeword(630) xor Codeword(689) xor Codeword(766) xor
                Codeword(819) xor Codeword(847) xor Codeword(915) xor Codeword(986) xor
                Codeword(1044) xor Codeword(1102) xor Codeword(1163) xor Codeword(1196) xor
                Codeword(1236) xor Codeword(1306) xor Codeword(1329) xor Codeword(1422) xor
                Codeword(1434) xor Codeword(1588) xor Codeword(1638) xor Codeword(1679) xor
                Codeword(1782) xor Codeword(1854) xor Codeword(1934) xor Codeword(1949);
 
     check279 <= Codeword(31) xor Codeword(58) xor Codeword(144) xor Codeword(219) xor
                Codeword(239) xor Codeword(368) xor Codeword(444) xor Codeword(450) xor
                Codeword(614) xor Codeword(660) xor Codeword(851) xor Codeword(939) xor
                Codeword(972) xor Codeword(1054) xor Codeword(1208) xor Codeword(1273) xor
                Codeword(1294) xor Codeword(1352) xor Codeword(1401) xor Codeword(1452) xor
                Codeword(1460) xor Codeword(1471) xor Codeword(1622) xor Codeword(1676) xor
                Codeword(1768) xor Codeword(1779) xor Codeword(1964) xor Codeword(1991) xor
                Codeword(2007) xor Codeword(2011) xor Codeword(2013) xor Codeword(2025);
 
     check280 <= Codeword(30) xor Codeword(84) xor Codeword(129) xor Codeword(215) xor
                Codeword(233) xor Codeword(310) xor Codeword(376) xor Codeword(445) xor
                Codeword(505) xor Codeword(555) xor Codeword(606) xor Codeword(675) xor
                Codeword(723) xor Codeword(824) xor Codeword(840) xor Codeword(989) xor
                Codeword(1049) xor Codeword(1084) xor Codeword(1136) xor Codeword(1223) xor
                Codeword(1229) xor Codeword(1316) xor Codeword(1360) xor Codeword(1386) xor
                Codeword(1424) xor Codeword(1600) xor Codeword(1708) xor Codeword(1740) xor
                Codeword(1777) xor Codeword(1896) xor Codeword(1924) xor Codeword(1927);
 
     check281 <= Codeword(29) xor Codeword(90) xor Codeword(163) xor Codeword(182) xor
                Codeword(236) xor Codeword(298) xor Codeword(340) xor Codeword(422) xor
                Codeword(449) xor Codeword(557) xor Codeword(569) xor Codeword(648) xor
                Codeword(700) xor Codeword(771) xor Codeword(799) xor Codeword(875) xor
                Codeword(931) xor Codeword(950) xor Codeword(1055) xor Codeword(1060) xor
                Codeword(1099) xor Codeword(1120) xor Codeword(1190) xor Codeword(1237) xor
                Codeword(1308) xor Codeword(1356) xor Codeword(1545) xor Codeword(1560) xor
                Codeword(1591) xor Codeword(1617) xor Codeword(1666) xor Codeword(1791);
 
     check282 <= Codeword(28) xor Codeword(74) xor Codeword(125) xor Codeword(200) xor
                Codeword(226) xor Codeword(338) xor Codeword(413) xor Codeword(500) xor
                Codeword(573) xor Codeword(626) xor Codeword(746) xor Codeword(859) xor
                Codeword(940) xor Codeword(960) xor Codeword(1043) xor Codeword(1203) xor
                Codeword(1265) xor Codeword(1298) xor Codeword(1331) xor Codeword(1361) xor
                Codeword(1388) xor Codeword(1541) xor Codeword(1605) xor Codeword(1627) xor
                Codeword(1766) xor Codeword(1785) xor Codeword(1974) xor Codeword(2003) xor
                Codeword(2009) xor Codeword(2040) xor Codeword(2041) xor Codeword(2047);
 
     check283 <= Codeword(27) xor Codeword(76) xor Codeword(153) xor Codeword(201) xor
                Codeword(260) xor Codeword(294) xor Codeword(374) xor Codeword(431) xor
                Codeword(482) xor Codeword(616) xor Codeword(650) xor Codeword(692) xor
                Codeword(756) xor Codeword(810) xor Codeword(870) xor Codeword(955) xor
                Codeword(1012) xor Codeword(1075) xor Codeword(1147) xor Codeword(1276) xor
                Codeword(1351) xor Codeword(1396) xor Codeword(1435) xor Codeword(1491) xor
                Codeword(1524) xor Codeword(1585) xor Codeword(1697) xor Codeword(1829) xor
                Codeword(1835) xor Codeword(1900) xor Codeword(1947) xor Codeword(1955);
 
     check284 <= Codeword(26) xor Codeword(100) xor Codeword(137) xor Codeword(181) xor
                Codeword(245) xor Codeword(320) xor Codeword(353) xor Codeword(436) xor
                Codeword(488) xor Codeword(517) xor Codeword(572) xor Codeword(662) xor
                Codeword(701) xor Codeword(749) xor Codeword(803) xor Codeword(881) xor
                Codeword(928) xor Codeword(961) xor Codeword(1018) xor Codeword(1088) xor
                Codeword(1128) xor Codeword(1164) xor Codeword(1211) xor Codeword(1252) xor
                Codeword(1291) xor Codeword(1374) xor Codeword(1418) xor Codeword(1432) xor
                Codeword(1583) xor Codeword(1640) xor Codeword(1684) xor Codeword(1792);
 
     check285 <= Codeword(25) xor Codeword(82) xor Codeword(165) xor Codeword(172) xor
                Codeword(255) xor Codeword(304) xor Codeword(355) xor Codeword(447) xor
                Codeword(456) xor Codeword(524) xor Codeword(567) xor Codeword(658) xor
                Codeword(674) xor Codeword(753) xor Codeword(780) xor Codeword(901) xor
                Codeword(949) xor Codeword(1081) xor Codeword(1139) xor Codeword(1178) xor
                Codeword(1232) xor Codeword(1281) xor Codeword(1288) xor Codeword(1380) xor
                Codeword(1419) xor Codeword(1474) xor Codeword(1504) xor Codeword(1593) xor
                Codeword(1701) xor Codeword(1731) xor Codeword(1755) xor Codeword(1865);
 
     check286 <= Codeword(24) xor Codeword(93) xor Codeword(155) xor Codeword(189) xor
                Codeword(267) xor Codeword(330) xor Codeword(341) xor Codeword(435) xor
                Codeword(454) xor Codeword(556) xor Codeword(603) xor Codeword(623) xor
                Codeword(688) xor Codeword(744) xor Codeword(790) xor Codeword(842) xor
                Codeword(887) xor Codeword(934) xor Codeword(975) xor Codeword(1005) xor
                Codeword(1148) xor Codeword(1192) xor Codeword(1254) xor Codeword(1333) xor
                Codeword(1364) xor Codeword(1507) xor Codeword(1589) xor Codeword(1643) xor
                Codeword(1659) xor Codeword(1752) xor Codeword(1764) xor Codeword(1866);
 
     check287 <= Codeword(23) xor Codeword(101) xor Codeword(142) xor Codeword(193) xor
                Codeword(240) xor Codeword(322) xor Codeword(375) xor Codeword(429) xor
                Codeword(486) xor Codeword(514) xor Codeword(610) xor Codeword(643) xor
                Codeword(716) xor Codeword(722) xor Codeword(724) xor Codeword(784) xor
                Codeword(884) xor Codeword(903) xor Codeword(981) xor Codeword(1028) xor
                Codeword(1068) xor Codeword(1121) xor Codeword(1188) xor Codeword(1267) xor
                Codeword(1296) xor Codeword(1334) xor Codeword(1366) xor Codeword(1476) xor
                Codeword(1551) xor Codeword(1611) xor Codeword(1687) xor Codeword(1793);
 
     check288 <= Codeword(22) xor Codeword(75) xor Codeword(161) xor Codeword(224) xor
                Codeword(228) xor Codeword(308) xor Codeword(337) xor Codeword(410) xor
                Codeword(468) xor Codeword(542) xor Codeword(578) xor Codeword(644) xor
                Codeword(695) xor Codeword(763) xor Codeword(787) xor Codeword(845) xor
                Codeword(916) xor Codeword(964) xor Codeword(1010) xor Codeword(1061) xor
                Codeword(1135) xor Codeword(1168) xor Codeword(1206) xor Codeword(1263) xor
                Codeword(1324) xor Codeword(1405) xor Codeword(1473) xor Codeword(1487) xor
                Codeword(1619) xor Codeword(1658) xor Codeword(1713) xor Codeword(1794);
 
     check289 <= Codeword(21) xor Codeword(89) xor Codeword(134) xor Codeword(192) xor
                Codeword(269) xor Codeword(327) xor Codeword(365) xor Codeword(418) xor
                Codeword(471) xor Codeword(519) xor Codeword(577) xor Codeword(622) xor
                Codeword(717) xor Codeword(774) xor Codeword(778) xor Codeword(913) xor
                Codeword(966) xor Codeword(1021) xor Codeword(1065) xor Codeword(1110) xor
                Codeword(1173) xor Codeword(1227) xor Codeword(1283) xor Codeword(1372) xor
                Codeword(1410) xor Codeword(1441) xor Codeword(1479) xor Codeword(1510) xor
                Codeword(1614) xor Codeword(1654) xor Codeword(1994) xor Codeword(1998);
 
     check290 <= Codeword(20) xor Codeword(60) xor Codeword(131) xor Codeword(187) xor
                Codeword(231) xor Codeword(350) xor Codeword(440) xor Codeword(457) xor
                Codeword(544) xor Codeword(608) xor Codeword(676) xor Codeword(730) xor
                Codeword(811) xor Codeword(872) xor Codeword(992) xor Codeword(1107) xor
                Codeword(1142) xor Codeword(1174) xor Codeword(1247) xor Codeword(1328) xor
                Codeword(1483) xor Codeword(1552) xor Codeword(1558) xor Codeword(1563) xor
                Codeword(1620) xor Codeword(1712) xor Codeword(1783) xor Codeword(1820) xor
                Codeword(1850) xor Codeword(1886) xor Codeword(1972) xor Codeword(1977);
 
     check291 <= Codeword(19) xor Codeword(96) xor Codeword(147) xor Codeword(223) xor
                Codeword(249) xor Codeword(377) xor Codeword(439) xor Codeword(487) xor
                Codeword(558) xor Codeword(590) xor Codeword(629) xor Codeword(673) xor
                Codeword(757) xor Codeword(796) xor Codeword(867) xor Codeword(896) xor
                Codeword(973) xor Codeword(1004) xor Codeword(1089) xor Codeword(1205) xor
                Codeword(1248) xor Codeword(1336) xor Codeword(1409) xor Codeword(1450) xor
                Codeword(1465) xor Codeword(1494) xor Codeword(1512) xor Codeword(1529) xor
                Codeword(1568) xor Codeword(1610) xor Codeword(1767) xor Codeword(1867);
 
     check292 <= Codeword(18) xor Codeword(62) xor Codeword(139) xor Codeword(177) xor
                Codeword(257) xor Codeword(313) xor Codeword(367) xor Codeword(416) xor
                Codeword(453) xor Codeword(554) xor Codeword(592) xor Codeword(633) xor
                Codeword(690) xor Codeword(745) xor Codeword(806) xor Codeword(873) xor
                Codeword(897) xor Codeword(985) xor Codeword(1017) xor Codeword(1074) xor
                Codeword(1122) xor Codeword(1197) xor Codeword(1226) xor Codeword(1321) xor
                Codeword(1365) xor Codeword(1403) xor Codeword(1575) xor Codeword(1594) xor
                Codeword(1630) xor Codeword(1663) xor Codeword(1705) xor Codeword(1795);
 
     check293 <= Codeword(17) xor Codeword(77) xor Codeword(113) xor Codeword(197) xor
                Codeword(306) xor Codeword(354) xor Codeword(397) xor Codeword(479) xor
                Codeword(516) xor Codeword(579) xor Codeword(668) xor Codeword(712) xor
                Codeword(732) xor Codeword(818) xor Codeword(864) xor Codeword(930) xor
                Codeword(993) xor Codeword(1045) xor Codeword(1085) xor Codeword(1119) xor
                Codeword(1214) xor Codeword(1274) xor Codeword(1302) xor Codeword(1379) xor
                Codeword(1448) xor Codeword(1548) xor Codeword(1567) xor Codeword(1582) xor
                Codeword(1636) xor Codeword(1662) xor Codeword(1696) xor Codeword(1796);
 
     check294 <= Codeword(16) xor Codeword(73) xor Codeword(123) xor Codeword(196) xor
                Codeword(258) xor Codeword(284) xor Codeword(373) xor Codeword(400) xor
                Codeword(465) xor Codeword(537) xor Codeword(609) xor Codeword(632) xor
                Codeword(713) xor Codeword(748) xor Codeword(791) xor Codeword(831) xor
                Codeword(922) xor Codeword(965) xor Codeword(1024) xor Codeword(1094) xor
                Codeword(1138) xor Codeword(1217) xor Codeword(1235) xor Codeword(1287) xor
                Codeword(1353) xor Codeword(1393) xor Codeword(1555) xor Codeword(1562) xor
                Codeword(1624) xor Codeword(1686) xor Codeword(1689) xor Codeword(1797);
 
     check295 <= Codeword(15) xor Codeword(92) xor Codeword(117) xor Codeword(175) xor
                Codeword(346) xor Codeword(441) xor Codeword(489) xor Codeword(538) xor
                Codeword(576) xor Codeword(628) xor Codeword(768) xor Codeword(837) xor
                Codeword(938) xor Codeword(1047) xor Codeword(1160) xor Codeword(1169) xor
                Codeword(1299) xor Codeword(1415) xor Codeword(1439) xor Codeword(1519) xor
                Codeword(1535) xor Codeword(1670) xor Codeword(1699) xor Codeword(1737) xor
                Codeword(1756) xor Codeword(1826) xor Codeword(1843) xor Codeword(1931) xor
                Codeword(1975) xor Codeword(1982) xor Codeword(1987) xor Codeword(1989);
 
     check296 <= Codeword(14) xor Codeword(55) xor Codeword(121) xor Codeword(208) xor
                Codeword(286) xor Codeword(343) xor Codeword(417) xor Codeword(481) xor
                Codeword(515) xor Codeword(665) xor Codeword(681) xor Codeword(820) xor
                Codeword(951) xor Codeword(1109) xor Codeword(1161) xor Codeword(1216) xor
                Codeword(1307) xor Codeword(1413) xor Codeword(1469) xor Codeword(1525) xor
                Codeword(1577) xor Codeword(1646) xor Codeword(1671) xor Codeword(1832) xor
                Codeword(1838) xor Codeword(1880) xor Codeword(1882) xor Codeword(1897) xor
                Codeword(1902) xor Codeword(1933) xor Codeword(1950) xor Codeword(1956);
 
     check297 <= Codeword(13) xor Codeword(56) xor Codeword(111) xor Codeword(211) xor
                Codeword(277) xor Codeword(290) xor Codeword(358) xor Codeword(438) xor
                Codeword(469) xor Codeword(508) xor Codeword(587) xor Codeword(620) xor
                Codeword(699) xor Codeword(772) xor Codeword(782) xor Codeword(878) xor
                Codeword(988) xor Codeword(1058) xor Codeword(1096) xor Codeword(1137) xor
                Codeword(1165) xor Codeword(1239) xor Codeword(1284) xor Codeword(1367) xor
                Codeword(1502) xor Codeword(1629) xor Codeword(1734) xor Codeword(1744) xor
                Codeword(1763) xor Codeword(1781) xor Codeword(1784) xor Codeword(1868);
 
     check298 <= Codeword(12) xor Codeword(91) xor Codeword(148) xor Codeword(198) xor
                Codeword(262) xor Codeword(282) xor Codeword(351) xor Codeword(408) xor
                Codeword(485) xor Codeword(523) xor Codeword(611) xor Codeword(639) xor
                Codeword(704) xor Codeword(776) xor Codeword(800) xor Codeword(849) xor
                Codeword(942) xor Codeword(953) xor Codeword(1020) xor Codeword(1129) xor
                Codeword(1194) xor Codeword(1224) xor Codeword(1234) xor Codeword(1323) xor
                Codeword(1495) xor Codeword(1508) xor Codeword(1572) xor Codeword(1602) xor
                Codeword(1639) xor Codeword(1772) xor Codeword(1776) xor Codeword(1869);
 
     check299 <= Codeword(83) xor Codeword(130) xor Codeword(176) xor Codeword(264) xor
                Codeword(314) xor Codeword(385) xor Codeword(393) xor Codeword(462) xor
                Codeword(527) xor Codeword(637) xor Codeword(767) xor Codeword(808) xor
                Codeword(885) xor Codeword(936) xor Codeword(967) xor Codeword(1040) xor
                Codeword(1079) xor Codeword(1146) xor Codeword(1201) xor Codeword(1271) xor
                Codeword(1382) xor Codeword(1451) xor Codeword(1467) xor Codeword(1477) xor
                Codeword(1498) xor Codeword(1538) xor Codeword(1647) xor Codeword(1733) xor
                Codeword(1746) xor Codeword(1883) xor Codeword(1889) xor Codeword(1912);
 
     check300 <= Codeword(11) xor Codeword(99) xor Codeword(143) xor Codeword(195) xor
                Codeword(299) xor Codeword(335) xor Codeword(419) xor Codeword(459) xor
                Codeword(591) xor Codeword(618) xor Codeword(703) xor Codeword(735) xor
                Codeword(804) xor Codeword(841) xor Codeword(920) xor Codeword(1041) xor
                Codeword(1087) xor Codeword(1151) xor Codeword(1326) xor Codeword(1348) xor
                Codeword(1426) xor Codeword(1497) xor Codeword(1518) xor Codeword(1522) xor
                Codeword(1557) xor Codeword(1587) xor Codeword(1625) xor Codeword(1680) xor
                Codeword(1774) xor Codeword(1831) xor Codeword(1859) xor Codeword(1894);
 
     check301 <= Codeword(10) xor Codeword(103) xor Codeword(154) xor Codeword(220) xor
                Codeword(270) xor Codeword(309) xor Codeword(389) xor Codeword(409) xor
                Codeword(474) xor Codeword(526) xor Codeword(697) xor Codeword(741) xor
                Codeword(809) xor Codeword(850) xor Codeword(983) xor Codeword(1019) xor
                Codeword(1082) xor Codeword(1243) xor Codeword(1349) xor Codeword(1428) xor
                Codeword(1514) xor Codeword(1553) xor Codeword(1691) xor Codeword(1773) xor
                Codeword(1812) xor Codeword(1847) xor Codeword(1855) xor Codeword(1856) xor
                Codeword(1903) xor Codeword(1904) xor Codeword(1916) xor Codeword(1920);
 
     check302 <= Codeword(9) xor Codeword(110) xor Codeword(124) xor Codeword(206) xor
                Codeword(227) xor Codeword(321) xor Codeword(398) xor Codeword(521) xor
                Codeword(583) xor Codeword(679) xor Codeword(725) xor Codeword(877) xor
                Codeword(892) xor Codeword(946) xor Codeword(1011) xor Codeword(1150) xor
                Codeword(1199) xor Codeword(1381) xor Codeword(1412) xor Codeword(1443) xor
                Codeword(1573) xor Codeword(1590) xor Codeword(1649) xor Codeword(1759) xor
                Codeword(1769) xor Codeword(1816) xor Codeword(1818) xor Codeword(1821) xor
                Codeword(1823) xor Codeword(1885) xor Codeword(1914) xor Codeword(1917);
 
     check303 <= Codeword(8) xor Codeword(102) xor Codeword(112) xor Codeword(178) xor
                Codeword(235) xor Codeword(293) xor Codeword(382) xor Codeword(415) xor
                Codeword(497) xor Codeword(506) xor Codeword(581) xor Codeword(640) xor
                Codeword(686) xor Codeword(727) xor Codeword(823) xor Codeword(836) xor
                Codeword(890) xor Codeword(947) xor Codeword(1003) xor Codeword(1027) xor
                Codeword(1078) xor Codeword(1144) xor Codeword(1181) xor Codeword(1373) xor
                Codeword(1468) xor Codeword(1520) xor Codeword(1546) xor Codeword(1592) xor
                Codeword(1642) xor Codeword(1681) xor Codeword(1762) xor Codeword(1870);
 
     check304 <= Codeword(7) xor Codeword(97) xor Codeword(157) xor Codeword(222) xor
                Codeword(263) xor Codeword(283) xor Codeword(359) xor Codeword(446) xor
                Codeword(451) xor Codeword(512) xor Codeword(595) xor Codeword(619) xor
                Codeword(709) xor Codeword(751) xor Codeword(828) xor Codeword(865) xor
                Codeword(925) xor Codeword(982) xor Codeword(1031) xor Codeword(1098) xor
                Codeword(1126) xor Codeword(1167) xor Codeword(1184) xor Codeword(1256) xor
                Codeword(1301) xor Codeword(1423) xor Codeword(1571) xor Codeword(1586) xor
                Codeword(1613) xor Codeword(1716) xor Codeword(1809) xor Codeword(1871);
 
     check305 <= Codeword(6) xor Codeword(80) xor Codeword(115) xor Codeword(209) xor
                Codeword(276) xor Codeword(323) xor Codeword(342) xor Codeword(443) xor
                Codeword(501) xor Codeword(533) xor Codeword(588) xor Codeword(636) xor
                Codeword(707) xor Codeword(733) xor Codeword(813) xor Codeword(844) xor
                Codeword(906) xor Codeword(974) xor Codeword(1104) xor Codeword(1112) xor
                Codeword(1133) xor Codeword(1170) xor Codeword(1258) xor Codeword(1292) xor
                Codeword(1338) xor Codeword(1436) xor Codeword(1505) xor Codeword(1604) xor
                Codeword(1626) xor Codeword(1685) xor Codeword(1702) xor Codeword(1798);
 
     check306 <= Codeword(5) xor Codeword(87) xor Codeword(136) xor Codeword(174) xor
                Codeword(402) xor Codeword(448) xor Codeword(531) xor Codeword(564) xor
                Codeword(663) xor Codeword(684) xor Codeword(815) xor Codeword(909) xor
                Codeword(1030) xor Codeword(1156) xor Codeword(1200) xor Codeword(1244) xor
                Codeword(1312) xor Codeword(1387) xor Codeword(1462) xor Codeword(1536) xor
                Codeword(1623) xor Codeword(1667) xor Codeword(1732) xor Codeword(1861) xor
                Codeword(1876) xor Codeword(1878) xor Codeword(1887) xor Codeword(1890) xor
                Codeword(1942) xor Codeword(1944) xor Codeword(2016) xor Codeword(2026);
 
     check307 <= Codeword(4) xor Codeword(107) xor Codeword(145) xor Codeword(202) xor
                Codeword(230) xor Codeword(302) xor Codeword(366) xor Codeword(395) xor
                Codeword(494) xor Codeword(510) xor Codeword(574) xor Codeword(649) xor
                Codeword(719) xor Codeword(752) xor Codeword(785) xor Codeword(879) xor
                Codeword(893) xor Codeword(996) xor Codeword(1025) xor Codeword(1091) xor
                Codeword(1154) xor Codeword(1318) xor Codeword(1470) xor Codeword(1521) xor
                Codeword(1537) xor Codeword(1637) xor Codeword(1665) xor Codeword(1745) xor
                Codeword(1748) xor Codeword(1923) xor Codeword(1932) xor Codeword(1940);
 
     check308 <= Codeword(140) xor Codeword(199) xor Codeword(251) xor Codeword(311) xor
                Codeword(336) xor Codeword(426) xor Codeword(475) xor Codeword(547) xor
                Codeword(568) xor Codeword(669) xor Codeword(726) xor Codeword(821) xor
                Codeword(876) xor Codeword(926) xor Codeword(1008) xor Codeword(1063) xor
                Codeword(1131) xor Codeword(1241) xor Codeword(1280) xor Codeword(1392) xor
                Codeword(1438) xor Codeword(1503) xor Codeword(1597) xor Codeword(1674) xor
                Codeword(1703) xor Codeword(1741) xor Codeword(1930) xor Codeword(1946) xor
                Codeword(1966) xor Codeword(1979) xor Codeword(2018) xor Codeword(2024);
 
     check309 <= Codeword(3) xor Codeword(86) xor Codeword(146) xor Codeword(214) xor
                Codeword(265) xor Codeword(307) xor Codeword(384) xor Codeword(437) xor
                Codeword(458) xor Codeword(550) xor Codeword(571) xor Codeword(664) xor
                Codeword(710) xor Codeword(740) xor Codeword(779) xor Codeword(839) xor
                Codeword(889) xor Codeword(995) xor Codeword(1015) xor Codeword(1097) xor
                Codeword(1177) xor Codeword(1268) xor Codeword(1304) xor Codeword(1370) xor
                Codeword(1420) xor Codeword(1427) xor Codeword(1481) xor Codeword(1513) xor
                Codeword(1715) xor Codeword(1730) xor Codeword(1742) xor Codeword(1872);
 
     check310 <= Codeword(2) xor Codeword(65) xor Codeword(135) xor Codeword(261) xor
                Codeword(312) xor Codeword(369) xor Codeword(430) xor Codeword(470) xor
                Codeword(534) xor Codeword(561) xor Codeword(653) xor Codeword(685) xor
                Codeword(786) xor Codeword(861) xor Codeword(917) xor Codeword(990) xor
                Codeword(1036) xor Codeword(1202) xor Codeword(1219) xor Codeword(1253) xor
                Codeword(1417) xor Codeword(1506) xor Codeword(1527) xor Codeword(1694) xor
                Codeword(1819) xor Codeword(1828) xor Codeword(1860) xor Codeword(1879) xor
                Codeword(1909) xor Codeword(1937) xor Codeword(1957) xor Codeword(1967);
 
     check311 <= Codeword(1) xor Codeword(68) xor Codeword(160) xor Codeword(225) xor
                Codeword(301) xor Codeword(387) xor Codeword(434) xor Codeword(480) xor
                Codeword(511) xor Codeword(596) xor Codeword(617) xor Codeword(706) xor
                Codeword(747) xor Codeword(814) xor Codeword(862) xor Codeword(902) xor
                Codeword(971) xor Codeword(1034) xor Codeword(1064) xor Codeword(1157) xor
                Codeword(1193) xor Codeword(1221) xor Codeword(1310) xor Codeword(1344) xor
                Codeword(1466) xor Codeword(1523) xor Codeword(1660) xor Codeword(1750) xor
                Codeword(1760) xor Codeword(1804) xor Codeword(1899) xor Codeword(1913);
 
     check312 <= Codeword(0) xor Codeword(108) xor Codeword(167) xor Codeword(246) xor
                Codeword(326) xor Codeword(348) xor Codeword(452) xor Codeword(530) xor
                Codeword(580) xor Codeword(645) xor Codeword(770) xor Codeword(827) xor
                Codeword(838) xor Codeword(927) xor Codeword(979) xor Codeword(1090) xor
                Codeword(1132) xor Codeword(1182) xor Codeword(1270) xor Codeword(1322) xor
                Codeword(1342) xor Codeword(1425) xor Codeword(1446) xor Codeword(1482) xor
                Codeword(1645) xor Codeword(1655) xor Codeword(1698) xor Codeword(1729) xor
                Codeword(1925) xor Codeword(1969) xor Codeword(2021) xor Codeword(2027);
 
     check313 <= Codeword(150) xor Codeword(188) xor Codeword(247) xor Codeword(356) xor
                Codeword(403) xor Codeword(496) xor Codeword(642) xor Codeword(728) xor
                Codeword(886) xor Codeword(919) xor Codeword(1001) xor Codeword(1050) xor
                Codeword(1103) xor Codeword(1278) xor Codeword(1376) xor Codeword(1400) xor
                Codeword(1489) xor Codeword(1528) xor Codeword(1596) xor Codeword(1710) xor
                Codeword(1723) xor Codeword(1814) xor Codeword(1830) xor Codeword(1881) xor
                Codeword(1919) xor Codeword(1953) xor Codeword(1973) xor Codeword(1983) xor
                Codeword(2022) xor Codeword(2034) xor Codeword(2038) xor Codeword(2044);
 
     check314 <= Codeword(191) xor Codeword(278) xor Codeword(316) xor Codeword(352) xor
                Codeword(442) xor Codeword(483) xor Codeword(543) xor Codeword(602) xor
                Codeword(656) xor Codeword(687) xor Codeword(781) xor Codeword(848) xor
                Codeword(907) xor Codeword(1053) xor Codeword(1123) xor Codeword(1357) xor
                Codeword(1389) xor Codeword(1411) xor Codeword(1461) xor Codeword(1556) xor
                Codeword(1648) xor Codeword(1651) xor Codeword(1717) xor Codeword(1749) xor
                Codeword(1836) xor Codeword(1853) xor Codeword(1907) xor Codeword(1926) xor
                Codeword(1928) xor Codeword(1938) xor Codeword(1958) xor Codeword(1968);
 
     check315 <= Codeword(78) xor Codeword(119) xor Codeword(183) xor Codeword(271) xor
                Codeword(318) xor Codeword(357) xor Codeword(399) xor Codeword(499) xor
                Codeword(513) xor Codeword(575) xor Codeword(651) xor Codeword(678) xor
                Codeword(743) xor Codeword(802) xor Codeword(853) xor Codeword(924) xor
                Codeword(977) xor Codeword(1037) xor Codeword(1111) xor Codeword(1172) xor
                Codeword(1249) xor Codeword(1317) xor Codeword(1359) xor Codeword(1404) xor
                Codeword(1447) xor Codeword(1457) xor Codeword(1488) xor Codeword(1511) xor
                Codeword(1675) xor Codeword(1714) xor Codeword(1722) xor Codeword(1799);
 
     check316 <= Codeword(61) xor Codeword(158) xor Codeword(234) xor Codeword(288) xor
                Codeword(347) xor Codeword(560) xor Codeword(563) xor Codeword(625) xor
                Codeword(720) xor Codeword(764) xor Codeword(816) xor Codeword(898) xor
                Codeword(956) xor Codeword(1014) xor Codeword(1080) xor Codeword(1134) xor
                Codeword(1186) xor Codeword(1220) xor Codeword(1246) xor Codeword(1293) xor
                Codeword(1345) xor Codeword(1408) xor Codeword(1501) xor Codeword(1569) xor
                Codeword(1664) xor Codeword(1721) xor Codeword(1727) xor Codeword(1754) xor
                Codeword(1961) xor Codeword(2014) xor Codeword(2035) xor Codeword(2039);
 
     check317 <= Codeword(88) xor Codeword(238) xor Codeword(324) xor Codeword(372) xor
                Codeword(472) xor Codeword(548) xor Codeword(604) xor Codeword(634) xor
                Codeword(683) xor Codeword(765) xor Codeword(812) xor Codeword(852) xor
                Codeword(895) xor Codeword(959) xor Codeword(1092) xor Codeword(1125) xor
                Codeword(1179) xor Codeword(1261) xor Codeword(1325) xor Codeword(1332) xor
                Codeword(1377) xor Codeword(1397) xor Codeword(1719) xor Codeword(1775) xor
                Codeword(1811) xor Codeword(1839) xor Codeword(1939) xor Codeword(1952) xor
                Codeword(1960) xor Codeword(1999) xor Codeword(2001) xor Codeword(2012);
 
     check318 <= Codeword(120) xor Codeword(210) xor Codeword(279) xor Codeword(379) xor
                Codeword(425) xor Codeword(467) xor Codeword(566) xor Codeword(742) xor
                Codeword(846) xor Codeword(911) xor Codeword(1002) xor Codeword(1006) xor
                Codeword(1059) xor Codeword(1210) xor Codeword(1295) xor Codeword(1341) xor
                Codeword(1540) xor Codeword(1566) xor Codeword(1598) xor Codeword(1634) xor
                Codeword(1720) xor Codeword(1805) xor Codeword(1837) xor Codeword(1877) xor
                Codeword(1935) xor Codeword(1976) xor Codeword(1980) xor Codeword(2005) xor
                Codeword(2008) xor Codeword(2036) xor Codeword(2037) xor Codeword(2045);
 
     check319 <= Codeword(52) xor Codeword(66) xor Codeword(151) xor Codeword(221) xor
                Codeword(237) xor Codeword(289) xor Codeword(361) xor Codeword(411) xor
                Codeword(473) xor Codeword(539) xor Codeword(585) xor Codeword(631) xor
                Codeword(711) xor Codeword(734) xor Codeword(797) xor Codeword(883) xor
                Codeword(904) xor Codeword(978) xor Codeword(1046) xor Codeword(1106) xor
                Codeword(1130) xor Codeword(1231) xor Codeword(1305) xor Codeword(1368) xor
                Codeword(1416) xor Codeword(1475) xor Codeword(1485) xor Codeword(1515) xor
                Codeword(1595) xor Codeword(1661) xor Codeword(1695) xor Codeword(1800);
 
     check320 <= Codeword(53) xor Codeword(126) xor Codeword(196) xor Codeword(295) xor
                Codeword(338) xor Codeword(439) xor Codeword(454) xor Codeword(531) xor
                Codeword(577) xor Codeword(637) xor Codeword(707) xor Codeword(759) xor
                Codeword(792) xor Codeword(856) xor Codeword(890) xor Codeword(1034) xor
                Codeword(1070) xor Codeword(1154) xor Codeword(1342) xor Codeword(1413) xor
                Codeword(1453) xor Codeword(1484) xor Codeword(1572) xor Codeword(1579) xor
                Codeword(1662) xor Codeword(1725) xor Codeword(1741) xor Codeword(1761) xor
                Codeword(1816) xor Codeword(1836) xor Codeword(1856) xor Codeword(1895);
 
     check321 <= Codeword(51) xor Codeword(65) xor Codeword(150) xor Codeword(220) xor
                Codeword(236) xor Codeword(288) xor Codeword(360) xor Codeword(410) xor
                Codeword(472) xor Codeword(538) xor Codeword(584) xor Codeword(630) xor
                Codeword(733) xor Codeword(882) xor Codeword(903) xor Codeword(977) xor
                Codeword(1045) xor Codeword(1105) xor Codeword(1217) xor Codeword(1230) xor
                Codeword(1304) xor Codeword(1367) xor Codeword(1474) xor Codeword(1558) xor
                Codeword(1594) xor Codeword(1660) xor Codeword(1759) xor Codeword(1831) xor
                Codeword(1929) xor Codeword(1992) xor Codeword(2003) xor Codeword(2013);
 
     check322 <= Codeword(50) xor Codeword(84) xor Codeword(165) xor Codeword(231) xor
                Codeword(316) xor Codeword(362) xor Codeword(427) xor Codeword(462) xor
                Codeword(535) xor Codeword(592) xor Codeword(623) xor Codeword(749) xor
                Codeword(797) xor Codeword(834) xor Codeword(932) xor Codeword(998) xor
                Codeword(1015) xor Codeword(1060) xor Codeword(1075) xor Codeword(1161) xor
                Codeword(1302) xor Codeword(1353) xor Codeword(1463) xor Codeword(1492) xor
                Codeword(1537) xor Codeword(1756) xor Codeword(1813) xor Codeword(1868) xor
                Codeword(1878) xor Codeword(1911) xor Codeword(1953) xor Codeword(1969);
 
     check323 <= Codeword(56) xor Codeword(136) xor Codeword(184) xor Codeword(268) xor
                Codeword(330) xor Codeword(390) xor Codeword(392) xor Codeword(484) xor
                Codeword(552) xor Codeword(588) xor Codeword(656) xor Codeword(717) xor
                Codeword(754) xor Codeword(828) xor Codeword(967) xor Codeword(1007) xor
                Codeword(1076) xor Codeword(1158) xor Codeword(1221) xor Codeword(1234) xor
                Codeword(1319) xor Codeword(1546) xor Codeword(1573) xor Codeword(1583) xor
                Codeword(1631) xor Codeword(1701) xor Codeword(1783) xor Codeword(1832) xor
                Codeword(1833) xor Codeword(1846) xor Codeword(1860) xor Codeword(1896);
 
     check324 <= Codeword(49) xor Codeword(109) xor Codeword(113) xor Codeword(223) xor
                Codeword(273) xor Codeword(302) xor Codeword(369) xor Codeword(400) xor
                Codeword(490) xor Codeword(544) xor Codeword(593) xor Codeword(640) xor
                Codeword(693) xor Codeword(821) xor Codeword(855) xor Codeword(936) xor
                Codeword(951) xor Codeword(1050) xor Codeword(1104) xor Codeword(1116) xor
                Codeword(1169) xor Codeword(1206) xor Codeword(1237) xor Codeword(1288) xor
                Codeword(1369) xor Codeword(1411) xor Codeword(1427) xor Codeword(1499) xor
                Codeword(1614) xor Codeword(1653) xor Codeword(1704) xor Codeword(1801);
 
     check325 <= Codeword(48) xor Codeword(70) xor Codeword(137) xor Codeword(185) xor
                Codeword(242) xor Codeword(284) xor Codeword(382) xor Codeword(395) xor
                Codeword(476) xor Codeword(518) xor Codeword(583) xor Codeword(653) xor
                Codeword(704) xor Codeword(753) xor Codeword(784) xor Codeword(832) xor
                Codeword(940) xor Codeword(979) xor Codeword(1012) xor Codeword(1097) xor
                Codeword(1186) xor Codeword(1227) xor Codeword(1289) xor Codeword(1357) xor
                Codeword(1398) xor Codeword(1436) xor Codeword(1462) xor Codeword(1512) xor
                Codeword(1554) xor Codeword(1617) xor Codeword(1718) xor Codeword(1802);
 
     check326 <= Codeword(47) xor Codeword(62) xor Codeword(203) xor Codeword(241) xor
                Codeword(304) xor Codeword(527) xor Codeword(606) xor Codeword(663) xor
                Codeword(697) xor Codeword(722) xor Codeword(748) xor Codeword(788) xor
                Codeword(867) xor Codeword(969) xor Codeword(1041) xor Codeword(1061) xor
                Codeword(1140) xor Codeword(1170) xor Codeword(1261) xor Codeword(1318) xor
                Codeword(1374) xor Codeword(1485) xor Codeword(1548) xor Codeword(1569) xor
                Codeword(1671) xor Codeword(1764) xor Codeword(1827) xor Codeword(1909) xor
                Codeword(1922) xor Codeword(1926) xor Codeword(1972) xor Codeword(1981);
 
     check327 <= Codeword(46) xor Codeword(94) xor Codeword(148) xor Codeword(211) xor
                Codeword(272) xor Codeword(318) xor Codeword(361) xor Codeword(446) xor
                Codeword(502) xor Codeword(521) xor Codeword(612) xor Codeword(634) xor
                Codeword(701) xor Codeword(777) xor Codeword(870) xor Codeword(911) xor
                Codeword(956) xor Codeword(1038) xor Codeword(1066) xor Codeword(1151) xor
                Codeword(1182) xor Codeword(1244) xor Codeword(1310) xor Codeword(1349) xor
                Codeword(1401) xor Codeword(1456) xor Codeword(1479) xor Codeword(1500) xor
                Codeword(1632) xor Codeword(1699) xor Codeword(1730) xor Codeword(1873);
 
     check328 <= Codeword(45) xor Codeword(103) xor Codeword(168) xor Codeword(314) xor
                Codeword(377) xor Codeword(413) xor Codeword(483) xor Codeword(524) xor
                Codeword(597) xor Codeword(690) xor Codeword(737) xor Codeword(787) xor
                Codeword(857) xor Codeword(893) xor Codeword(975) xor Codeword(1055) xor
                Codeword(1144) xor Codeword(1328) xor Codeword(1346) xor Codeword(1421) xor
                Codeword(1439) xor Codeword(1486) xor Codeword(1491) xor Codeword(1509) xor
                Codeword(1672) xor Codeword(1688) xor Codeword(1742) xor Codeword(1796) xor
                Codeword(1814) xor Codeword(1936) xor Codeword(1946) xor Codeword(1957);
 
     check329 <= Codeword(44) xor Codeword(97) xor Codeword(131) xor Codeword(212) xor
                Codeword(255) xor Codeword(280) xor Codeword(348) xor Codeword(420) xor
                Codeword(494) xor Codeword(516) xor Codeword(599) xor Codeword(665) xor
                Codeword(671) xor Codeword(760) xor Codeword(782) xor Codeword(833) xor
                Codeword(907) xor Codeword(947) xor Codeword(1047) xor Codeword(1065) xor
                Codeword(1148) xor Codeword(1268) xor Codeword(1278) xor Codeword(1361) xor
                Codeword(1515) xor Codeword(1530) xor Codeword(1538) xor Codeword(1560) xor
                Codeword(1607) xor Codeword(1626) xor Codeword(1667) xor Codeword(1803);
 
     check330 <= Codeword(43) xor Codeword(101) xor Codeword(132) xor Codeword(202) xor
                Codeword(243) xor Codeword(385) xor Codeword(404) xor Codeword(503) xor
                Codeword(553) xor Codeword(569) xor Codeword(626) xor Codeword(710) xor
                Codeword(758) xor Codeword(819) xor Codeword(917) xor Codeword(944) xor
                Codeword(1022) xor Codeword(1138) xor Codeword(1208) xor Codeword(1240) xor
                Codeword(1384) xor Codeword(1425) xor Codeword(1483) xor Codeword(1508) xor
                Codeword(1532) xor Codeword(1684) xor Codeword(1747) xor Codeword(1795) xor
                Codeword(1823) xor Codeword(1865) xor Codeword(1867) xor Codeword(1897);
 
     check331 <= Codeword(42) xor Codeword(92) xor Codeword(167) xor Codeword(172) xor
                Codeword(350) xor Codeword(406) xor Codeword(534) xor Codeword(604) xor
                Codeword(646) xor Codeword(720) xor Codeword(736) xor Codeword(826) xor
                Codeword(879) xor Codeword(943) xor Codeword(961) xor Codeword(1031) xor
                Codeword(1117) xor Codeword(1194) xor Codeword(1229) xor Codeword(1428) xor
                Codeword(1449) xor Codeword(1477) xor Codeword(1529) xor Codeword(1533) xor
                Codeword(1634) xor Codeword(1650) xor Codeword(1706) xor Codeword(1753) xor
                Codeword(1862) xor Codeword(1963) xor Codeword(1991) xor Codeword(1993);
 
     check332 <= Codeword(41) xor Codeword(71) xor Codeword(158) xor Codeword(179) xor
                Codeword(240) xor Codeword(363) xor Codeword(431) xor Codeword(489) xor
                Codeword(548) xor Codeword(561) xor Codeword(772) xor Codeword(793) xor
                Codeword(865) xor Codeword(931) xor Codeword(953) xor Codeword(1025) xor
                Codeword(1157) xor Codeword(1211) xor Codeword(1271) xor Codeword(1326) xor
                Codeword(1338) xor Codeword(1389) xor Codeword(1420) xor Codeword(1600) xor
                Codeword(1627) xor Codeword(1676) xor Codeword(1724) xor Codeword(1782) xor
                Codeword(1885) xor Codeword(1925) xor Codeword(2022) xor Codeword(2029);
 
     check333 <= Codeword(108) xor Codeword(117) xor Codeword(215) xor Codeword(265) xor
                Codeword(324) xor Codeword(359) xor Codeword(411) xor Codeword(651) xor
                Codeword(774) xor Codeword(835) xor Codeword(920) xor Codeword(986) xor
                Codeword(1071) xor Codeword(1175) xor Codeword(1232) xor Codeword(1308) xor
                Codeword(1429) xor Codeword(1448) xor Codeword(1458) xor Codeword(1551) xor
                Codeword(1615) xor Codeword(1726) xor Codeword(1776) xor Codeword(1810) xor
                Codeword(1820) xor Codeword(1888) xor Codeword(1961) xor Codeword(1980) xor
                Codeword(2018) xor Codeword(2019) xor Codeword(2020) xor Codeword(2034);
 
     check334 <= Codeword(40) xor Codeword(66) xor Codeword(217) xor Codeword(286) xor
                Codeword(380) xor Codeword(497) xor Codeword(528) xor Codeword(598) xor
                Codeword(654) xor Codeword(692) xor Codeword(761) xor Codeword(824) xor
                Codeword(881) xor Codeword(934) xor Codeword(996) xor Codeword(1020) xor
                Codeword(1069) xor Codeword(1123) xor Codeword(1184) xor Codeword(1250) xor
                Codeword(1314) xor Codeword(1336) xor Codeword(1394) xor Codeword(1443) xor
                Codeword(1630) xor Codeword(1712) xor Codeword(1755) xor Codeword(1852) xor
                Codeword(1913) xor Codeword(1997) xor Codeword(2021) xor Codeword(2026);
 
     check335 <= Codeword(39) xor Codeword(78) xor Codeword(170) xor Codeword(189) xor
                Codeword(274) xor Codeword(291) xor Codeword(343) xor Codeword(432) xor
                Codeword(465) xor Codeword(517) xor Codeword(611) xor Codeword(645) xor
                Codeword(679) xor Codeword(804) xor Codeword(868) xor Codeword(899) xor
                Codeword(990) xor Codeword(1056) xor Codeword(1099) xor Codeword(1152) xor
                Codeword(1179) xor Codeword(1258) xor Codeword(1276) xor Codeword(1285) xor
                Codeword(1382) xor Codeword(1441) xor Codeword(1541) xor Codeword(1578) xor
                Codeword(1682) xor Codeword(1845) xor Codeword(1872) xor Codeword(1898);
 
     check336 <= Codeword(38) xor Codeword(104) xor Codeword(121) xor Codeword(267) xor
                Codeword(332) xor Codeword(344) xor Codeword(405) xor Codeword(477) xor
                Codeword(506) xor Codeword(585) xor Codeword(695) xor Codeword(757) xor
                Codeword(806) xor Codeword(831) xor Codeword(909) xor Codeword(993) xor
                Codeword(1037) xor Codeword(1082) xor Codeword(1139) xor Codeword(1185) xor
                Codeword(1329) xor Codeword(1362) xor Codeword(1471) xor Codeword(1543) xor
                Codeword(1605) xor Codeword(1651) xor Codeword(1692) xor Codeword(1740) xor
                Codeword(1850) xor Codeword(1935) xor Codeword(1951) xor Codeword(1970);
 
     check337 <= Codeword(37) xor Codeword(93) xor Codeword(115) xor Codeword(183) xor
                Codeword(253) xor Codeword(290) xor Codeword(379) xor Codeword(419) xor
                Codeword(475) xor Codeword(519) xor Codeword(564) xor Codeword(714) xor
                Codeword(728) xor Codeword(794) xor Codeword(862) xor Codeword(904) xor
                Codeword(983) xor Codeword(1051) xor Codeword(1085) xor Codeword(1126) xor
                Codeword(1259) xor Codeword(1345) xor Codeword(1405) xor Codeword(1432) xor
                Codeword(1454) xor Codeword(1590) xor Codeword(1620) xor Codeword(1656) xor
                Codeword(1705) xor Codeword(1927) xor Codeword(1947) xor Codeword(1958);
 
     check338 <= Codeword(36) xor Codeword(80) xor Codeword(155) xor Codeword(190) xor
                Codeword(370) xor Codeword(492) xor Codeword(540) xor Codeword(587) xor
                Codeword(658) xor Codeword(669) xor Codeword(825) xor Codeword(859) xor
                Codeword(962) xor Codeword(1006) xor Codeword(1072) xor Codeword(1142) xor
                Codeword(1197) xor Codeword(1249) xor Codeword(1434) xor Codeword(1452) xor
                Codeword(1549) xor Codeword(1613) xor Codeword(1677) xor Codeword(1717) xor
                Codeword(1732) xor Codeword(1770) xor Codeword(1797) xor Codeword(1819) xor
                Codeword(1822) xor Codeword(1870) xor Codeword(1933) xor Codeword(1941);
 
     check339 <= Codeword(35) xor Codeword(96) xor Codeword(163) xor Codeword(216) xor
                Codeword(247) xor Codeword(322) xor Codeword(389) xor Codeword(426) xor
                Codeword(459) xor Codeword(550) xor Codeword(600) xor Codeword(660) xor
                Codeword(718) xor Codeword(738) xor Codeword(791) xor Codeword(873) xor
                Codeword(898) xor Codeword(1002) xor Codeword(1032) xor Codeword(1100) xor
                Codeword(1163) xor Codeword(1203) xor Codeword(1274) xor Codeword(1281) xor
                Codeword(1299) xor Codeword(1368) xor Codeword(1397) xor Codeword(1563) xor
                Codeword(1580) xor Codeword(1640) xor Codeword(1649) xor Codeword(1804);
 
     check340 <= Codeword(34) xor Codeword(58) xor Codeword(127) xor Codeword(178) xor
                Codeword(245) xor Codeword(334) xor Codeword(393) xor Codeword(460) xor
                Codeword(545) xor Codeword(596) xor Codeword(629) xor Codeword(670) xor
                Codeword(730) xor Codeword(816) xor Codeword(922) xor Codeword(957) xor
                Codeword(1021) xor Codeword(1112) xor Codeword(1188) xor Codeword(1339) xor
                Codeword(1406) xor Codeword(1489) xor Codeword(1524) xor Codeword(1606) xor
                Codeword(1693) xor Codeword(1765) xor Codeword(1788) xor Codeword(1828) xor
                Codeword(1887) xor Codeword(1974) xor Codeword(1978) xor Codeword(1982);
 
     check341 <= Codeword(33) xor Codeword(68) xor Codeword(125) xor Codeword(204) xor
                Codeword(258) xor Codeword(296) xor Codeword(491) xor Codeword(551) xor
                Codeword(614) xor Codeword(666) xor Codeword(842) xor Codeword(928) xor
                Codeword(968) xor Codeword(1008) xor Codeword(1092) xor Codeword(1165) xor
                Codeword(1190) xor Codeword(1263) xor Codeword(1313) xor Codeword(1475) xor
                Codeword(1496) xor Codeword(1542) xor Codeword(1577) xor Codeword(1727) xor
                Codeword(1767) xor Codeword(1824) xor Codeword(1864) xor Codeword(1879) xor
                Codeword(1943) xor Codeword(1976) xor Codeword(1977) xor Codeword(1983);
 
     check342 <= Codeword(32) xor Codeword(63) xor Codeword(161) xor Codeword(251) xor
                Codeword(294) xor Codeword(403) xor Codeword(539) xor Codeword(581) xor
                Codeword(624) xor Codeword(681) xor Codeword(735) xor Codeword(853) xor
                Codeword(913) xor Codeword(997) xor Codeword(1024) xor Codeword(1115) xor
                Codeword(1214) xor Codeword(1265) xor Codeword(1284) xor Codeword(1370) xor
                Codeword(1455) xor Codeword(1564) xor Codeword(1598) xor Codeword(1647) xor
                Codeword(1711) xor Codeword(1769) xor Codeword(1773) xor Codeword(1798) xor
                Codeword(1815) xor Codeword(1840) xor Codeword(1853) xor Codeword(1899);
 
     check343 <= Codeword(31) xor Codeword(69) xor Codeword(140) xor Codeword(206) xor
                Codeword(228) xor Codeword(327) xor Codeword(387) xor Codeword(422) xor
                Codeword(501) xor Codeword(508) xor Codeword(582) xor Codeword(688) xor
                Codeword(765) xor Codeword(818) xor Codeword(846) xor Codeword(985) xor
                Codeword(1043) xor Codeword(1101) xor Codeword(1162) xor Codeword(1195) xor
                Codeword(1235) xor Codeword(1282) xor Codeword(1305) xor Codeword(1433) xor
                Codeword(1535) xor Codeword(1637) xor Codeword(1678) xor Codeword(1691) xor
                Codeword(1799) xor Codeword(1825) xor Codeword(1841) xor Codeword(1900);
 
     check344 <= Codeword(30) xor Codeword(57) xor Codeword(143) xor Codeword(218) xor
                Codeword(238) xor Codeword(307) xor Codeword(367) xor Codeword(443) xor
                Codeword(449) xor Codeword(514) xor Codeword(613) xor Codeword(659) xor
                Codeword(673) xor Codeword(763) xor Codeword(805) xor Codeword(850) xor
                Codeword(938) xor Codeword(971) xor Codeword(1053) xor Codeword(1094) xor
                Codeword(1129) xor Codeword(1207) xor Codeword(1272) xor Codeword(1293) xor
                Codeword(1351) xor Codeword(1400) xor Codeword(1451) xor Codeword(1459) xor
                Codeword(1470) xor Codeword(1621) xor Codeword(1675) xor Codeword(1805);
 
     check345 <= Codeword(29) xor Codeword(83) xor Codeword(128) xor Codeword(232) xor
                Codeword(309) xor Codeword(375) xor Codeword(444) xor Codeword(505) xor
                Codeword(554) xor Codeword(605) xor Codeword(674) xor Codeword(776) xor
                Codeword(823) xor Codeword(839) xor Codeword(921) xor Codeword(988) xor
                Codeword(1048) xor Codeword(1083) xor Codeword(1135) xor Codeword(1222) xor
                Codeword(1228) xor Codeword(1315) xor Codeword(1359) xor Codeword(1385) xor
                Codeword(1423) xor Codeword(1493) xor Codeword(1737) xor Codeword(1835) xor
                Codeword(1966) xor Codeword(1994) xor Codeword(2004) xor Codeword(2014);
 
     check346 <= Codeword(28) xor Codeword(89) xor Codeword(162) xor Codeword(181) xor
                Codeword(235) xor Codeword(297) xor Codeword(339) xor Codeword(421) xor
                Codeword(448) xor Codeword(556) xor Codeword(568) xor Codeword(647) xor
                Codeword(699) xor Codeword(770) xor Codeword(798) xor Codeword(874) xor
                Codeword(949) xor Codeword(1054) xor Codeword(1059) xor Codeword(1098) xor
                Codeword(1119) xor Codeword(1189) xor Codeword(1236) xor Codeword(1307) xor
                Codeword(1355) xor Codeword(1457) xor Codeword(1544) xor Codeword(1616) xor
                Codeword(1665) xor Codeword(1746) xor Codeword(1789) xor Codeword(1874);
 
     check347 <= Codeword(27) xor Codeword(73) xor Codeword(124) xor Codeword(199) xor
                Codeword(225) xor Codeword(328) xor Codeword(337) xor Codeword(412) xor
                Codeword(499) xor Codeword(523) xor Codeword(572) xor Codeword(625) xor
                Codeword(680) xor Codeword(745) xor Codeword(796) xor Codeword(858) xor
                Codeword(939) xor Codeword(959) xor Codeword(1042) xor Codeword(1077) xor
                Codeword(1121) xor Codeword(1202) xor Codeword(1264) xor Codeword(1297) xor
                Codeword(1330) xor Codeword(1360) xor Codeword(1387) xor Codeword(1540) xor
                Codeword(1604) xor Codeword(1666) xor Codeword(1710) xor Codeword(1806);
 
     check348 <= Codeword(26) xor Codeword(75) xor Codeword(152) xor Codeword(200) xor
                Codeword(259) xor Codeword(293) xor Codeword(373) xor Codeword(430) xor
                Codeword(481) xor Codeword(507) xor Codeword(616) xor Codeword(649) xor
                Codeword(691) xor Codeword(755) xor Codeword(809) xor Codeword(869) xor
                Codeword(914) xor Codeword(954) xor Codeword(1011) xor Codeword(1074) xor
                Codeword(1146) xor Codeword(1176) xor Codeword(1224) xor Codeword(1312) xor
                Codeword(1350) xor Codeword(1490) xor Codeword(1523) xor Codeword(1584) xor
                Codeword(1696) xor Codeword(1752) xor Codeword(1908) xor Codeword(1918);
 
     check349 <= Codeword(25) xor Codeword(99) xor Codeword(180) xor Codeword(244) xor
                Codeword(319) xor Codeword(352) xor Codeword(435) xor Codeword(487) xor
                Codeword(571) xor Codeword(661) xor Codeword(700) xor Codeword(802) xor
                Codeword(880) xor Codeword(927) xor Codeword(960) xor Codeword(1017) xor
                Codeword(1113) xor Codeword(1127) xor Codeword(1210) xor Codeword(1251) xor
                Codeword(1290) xor Codeword(1373) xor Codeword(1417) xor Codeword(1431) xor
                Codeword(1582) xor Codeword(1639) xor Codeword(1683) xor Codeword(1728) xor
                Codeword(1818) xor Codeword(1842) xor Codeword(1863) xor Codeword(1901);
 
     check350 <= Codeword(24) xor Codeword(81) xor Codeword(164) xor Codeword(171) xor
                Codeword(254) xor Codeword(303) xor Codeword(447) xor Codeword(455) xor
                Codeword(566) xor Codeword(657) xor Codeword(752) xor Codeword(854) xor
                Codeword(900) xor Codeword(948) xor Codeword(1058) xor Codeword(1080) xor
                Codeword(1177) xor Codeword(1231) xor Codeword(1280) xor Codeword(1287) xor
                Codeword(1379) xor Codeword(1418) xor Codeword(1473) xor Codeword(1592) xor
                Codeword(1655) xor Codeword(1700) xor Codeword(1839) xor Codeword(1942) xor
                Codeword(1964) xor Codeword(1987) xor Codeword(2043) xor Codeword(2047);
 
     check351 <= Codeword(23) xor Codeword(154) xor Codeword(188) xor Codeword(266) xor
                Codeword(329) xor Codeword(340) xor Codeword(434) xor Codeword(453) xor
                Codeword(555) xor Codeword(622) xor Codeword(687) xor Codeword(743) xor
                Codeword(789) xor Codeword(830) xor Codeword(841) xor Codeword(933) xor
                Codeword(974) xor Codeword(1004) xor Codeword(1109) xor Codeword(1147) xor
                Codeword(1191) xor Codeword(1253) xor Codeword(1301) xor Codeword(1395) xor
                Codeword(1642) xor Codeword(1658) xor Codeword(1703) xor Codeword(1869) xor
                Codeword(1883) xor Codeword(1996) xor Codeword(2012) xor Codeword(2027);
 
     check352 <= Codeword(22) xor Codeword(100) xor Codeword(141) xor Codeword(192) xor
                Codeword(239) xor Codeword(321) xor Codeword(374) xor Codeword(428) xor
                Codeword(485) xor Codeword(513) xor Codeword(609) xor Codeword(642) xor
                Codeword(715) xor Codeword(723) xor Codeword(783) xor Codeword(883) xor
                Codeword(902) xor Codeword(1027) xor Codeword(1067) xor Codeword(1120) xor
                Codeword(1187) xor Codeword(1266) xor Codeword(1295) xor Codeword(1333) xor
                Codeword(1365) xor Codeword(1550) xor Codeword(1610) xor Codeword(1687) xor
                Codeword(1754) xor Codeword(1784) xor Codeword(1843) xor Codeword(1902);
 
     check353 <= Codeword(21) xor Codeword(74) xor Codeword(160) xor Codeword(224) xor
                Codeword(227) xor Codeword(336) xor Codeword(409) xor Codeword(467) xor
                Codeword(541) xor Codeword(643) xor Codeword(694) xor Codeword(762) xor
                Codeword(786) xor Codeword(844) xor Codeword(915) xor Codeword(1009) xor
                Codeword(1134) xor Codeword(1205) xor Codeword(1262) xor Codeword(1323) xor
                Codeword(1404) xor Codeword(1472) xor Codeword(1576) xor Codeword(1618) xor
                Codeword(1780) xor Codeword(1791) xor Codeword(1871) xor Codeword(1881) xor
                Codeword(1890) xor Codeword(1894) xor Codeword(2011) xor Codeword(2028);
 
     check354 <= Codeword(20) xor Codeword(88) xor Codeword(133) xor Codeword(191) xor
                Codeword(326) xor Codeword(364) xor Codeword(417) xor Codeword(470) xor
                Codeword(576) xor Codeword(621) xor Codeword(773) xor Codeword(864) xor
                Codeword(912) xor Codeword(965) xor Codeword(1064) xor Codeword(1108) xor
                Codeword(1172) xor Codeword(1226) xor Codeword(1371) xor Codeword(1409) xor
                Codeword(1440) xor Codeword(1478) xor Codeword(1531) xor Codeword(1707) xor
                Codeword(1738) xor Codeword(1817) xor Codeword(1877) xor Codeword(1892) xor
                Codeword(1921) xor Codeword(1973) xor Codeword(2002) xor Codeword(2015);
 
     check355 <= Codeword(19) xor Codeword(59) xor Codeword(130) xor Codeword(186) xor
                Codeword(230) xor Codeword(300) xor Codeword(349) xor Codeword(456) xor
                Codeword(543) xor Codeword(667) xor Codeword(675) xor Codeword(729) xor
                Codeword(810) xor Codeword(871) xor Codeword(930) xor Codeword(1028) xor
                Codeword(1106) xor Codeword(1141) xor Codeword(1173) xor Codeword(1246) xor
                Codeword(1327) xor Codeword(1383) xor Codeword(1482) xor Codeword(1552) xor
                Codeword(1557) xor Codeword(1619) xor Codeword(1681) xor Codeword(1847) xor
                Codeword(1990) xor Codeword(2000) xor Codeword(2001) xor Codeword(2016);
 
     check356 <= Codeword(18) xor Codeword(95) xor Codeword(146) xor Codeword(222) xor
                Codeword(299) xor Codeword(376) xor Codeword(438) xor Codeword(486) xor
                Codeword(557) xor Codeword(589) xor Codeword(672) xor Codeword(756) xor
                Codeword(795) xor Codeword(895) xor Codeword(972) xor Codeword(1088) xor
                Codeword(1204) xor Codeword(1247) xor Codeword(1408) xor Codeword(1464) xor
                Codeword(1495) xor Codeword(1504) xor Codeword(1511) xor Codeword(1528) xor
                Codeword(1567) xor Codeword(1609) xor Codeword(1736) xor Codeword(1794) xor
                Codeword(1893) xor Codeword(1931) xor Codeword(2005) xor Codeword(2006);
 
     check357 <= Codeword(17) xor Codeword(61) xor Codeword(138) xor Codeword(176) xor
                Codeword(256) xor Codeword(312) xor Codeword(366) xor Codeword(415) xor
                Codeword(452) xor Codeword(632) xor Codeword(872) xor Codeword(896) xor
                Codeword(984) xor Codeword(1016) xor Codeword(1073) xor Codeword(1196) xor
                Codeword(1225) xor Codeword(1320) xor Codeword(1364) xor Codeword(1402) xor
                Codeword(1444) xor Codeword(1575) xor Codeword(1593) xor Codeword(1760) xor
                Codeword(1792) xor Codeword(1830) xor Codeword(1876) xor Codeword(1962) xor
                Codeword(1975) xor Codeword(2025) xor Codeword(2032) xor Codeword(2041);
 
     check358 <= Codeword(16) xor Codeword(76) xor Codeword(112) xor Codeword(252) xor
                Codeword(305) xor Codeword(353) xor Codeword(396) xor Codeword(478) xor
                Codeword(515) xor Codeword(578) xor Codeword(668) xor Codeword(711) xor
                Codeword(731) xor Codeword(817) xor Codeword(863) xor Codeword(929) xor
                Codeword(992) xor Codeword(1044) xor Codeword(1084) xor Codeword(1118) xor
                Codeword(1213) xor Codeword(1273) xor Codeword(1378) xor Codeword(1447) xor
                Codeword(1566) xor Codeword(1581) xor Codeword(1733) xor Codeword(1812) xor
                Codeword(1866) xor Codeword(1932) xor Codeword(1944) xor Codeword(1959);
 
     check359 <= Codeword(15) xor Codeword(72) xor Codeword(122) xor Codeword(195) xor
                Codeword(257) xor Codeword(283) xor Codeword(372) xor Codeword(399) xor
                Codeword(464) xor Codeword(536) xor Codeword(608) xor Codeword(631) xor
                Codeword(712) xor Codeword(747) xor Codeword(790) xor Codeword(886) xor
                Codeword(964) xor Codeword(1023) xor Codeword(1093) xor Codeword(1137) xor
                Codeword(1216) xor Codeword(1286) xor Codeword(1352) xor Codeword(1561) xor
                Codeword(1591) xor Codeword(1623) xor Codeword(1685) xor Codeword(1743) xor
                Codeword(1771) xor Codeword(1834) xor Codeword(1920) xor Codeword(1924);
 
     check360 <= Codeword(14) xor Codeword(91) xor Codeword(116) xor Codeword(174) xor
                Codeword(248) xor Codeword(292) xor Codeword(345) xor Codeword(440) xor
                Codeword(488) xor Codeword(537) xor Codeword(575) xor Codeword(627) xor
                Codeword(689) xor Codeword(767) xor Codeword(779) xor Codeword(836) xor
                Codeword(937) xor Codeword(980) xor Codeword(1046) xor Codeword(1068) xor
                Codeword(1159) xor Codeword(1168) xor Codeword(1239) xor Codeword(1298) xor
                Codeword(1414) xor Codeword(1438) xor Codeword(1519) xor Codeword(1534) xor
                Codeword(1599) xor Codeword(1625) xor Codeword(1698) xor Codeword(1807);
 
     check361 <= Codeword(13) xor Codeword(54) xor Codeword(120) xor Codeword(207) xor
                Codeword(271) xor Codeword(285) xor Codeword(342) xor Codeword(391) xor
                Codeword(416) xor Codeword(480) xor Codeword(601) xor Codeword(664) xor
                Codeword(775) xor Codeword(876) xor Codeword(942) xor Codeword(950) xor
                Codeword(1005) xor Codeword(1160) xor Codeword(1215) xor Codeword(1306) xor
                Codeword(1354) xor Codeword(1412) xor Codeword(1468) xor Codeword(1487) xor
                Codeword(1506) xor Codeword(1525) xor Codeword(1645) xor Codeword(1774) xor
                Codeword(1811) xor Codeword(1915) xor Codeword(2007) xor Codeword(2009);
 
     check362 <= Codeword(12) xor Codeword(55) xor Codeword(169) xor Codeword(210) xor
                Codeword(276) xor Codeword(289) xor Codeword(357) xor Codeword(468) xor
                Codeword(586) xor Codeword(619) xor Codeword(698) xor Codeword(771) xor
                Codeword(781) xor Codeword(877) xor Codeword(987) xor Codeword(1057) xor
                Codeword(1095) xor Codeword(1136) xor Codeword(1164) xor Codeword(1212) xor
                Codeword(1238) xor Codeword(1283) xor Codeword(1366) xor Codeword(1392) xor
                Codeword(1466) xor Codeword(1502) xor Codeword(1663) xor Codeword(1731) xor
                Codeword(1739) xor Codeword(1829) xor Codeword(1995) xor Codeword(1999);
 
     check363 <= Codeword(90) xor Codeword(147) xor Codeword(197) xor Codeword(261) xor
                Codeword(281) xor Codeword(407) xor Codeword(522) xor Codeword(610) xor
                Codeword(638) xor Codeword(703) xor Codeword(848) xor Codeword(941) xor
                Codeword(952) xor Codeword(1019) xor Codeword(1111) xor Codeword(1128) xor
                Codeword(1193) xor Codeword(1223) xor Codeword(1233) xor Codeword(1322) xor
                Codeword(1363) xor Codeword(1571) xor Codeword(1601) xor Codeword(1638) xor
                Codeword(1686) xor Codeword(1785) xor Codeword(1821) xor Codeword(1858) xor
                Codeword(1889) xor Codeword(1945) xor Codeword(1956) xor Codeword(1965);
 
     check364 <= Codeword(11) xor Codeword(82) xor Codeword(129) xor Codeword(175) xor
                Codeword(263) xor Codeword(313) xor Codeword(384) xor Codeword(461) xor
                Codeword(526) xor Codeword(602) xor Codeword(636) xor Codeword(766) xor
                Codeword(807) xor Codeword(884) xor Codeword(935) xor Codeword(966) xor
                Codeword(1039) xor Codeword(1078) xor Codeword(1145) xor Codeword(1200) xor
                Codeword(1270) xor Codeword(1309) xor Codeword(1381) xor Codeword(1450) xor
                Codeword(1498) xor Codeword(1646) xor Codeword(1661) xor Codeword(1763) xor
                Codeword(1786) xor Codeword(1967) xor Codeword(2035) xor Codeword(2042);
 
     check365 <= Codeword(10) xor Codeword(98) xor Codeword(142) xor Codeword(194) xor
                Codeword(234) xor Codeword(298) xor Codeword(418) xor Codeword(458) xor
                Codeword(590) xor Codeword(617) xor Codeword(702) xor Codeword(734) xor
                Codeword(803) xor Codeword(840) xor Codeword(919) xor Codeword(963) xor
                Codeword(1040) xor Codeword(1086) xor Codeword(1150) xor Codeword(1325) xor
                Codeword(1347) xor Codeword(1390) xor Codeword(1415) xor Codeword(1497) xor
                Codeword(1517) xor Codeword(1521) xor Codeword(1556) xor Codeword(1586) xor
                Codeword(1624) xor Codeword(1679) xor Codeword(1768) xor Codeword(1875);
 
     check366 <= Codeword(9) xor Codeword(102) xor Codeword(153) xor Codeword(219) xor
                Codeword(269) xor Codeword(308) xor Codeword(388) xor Codeword(473) xor
                Codeword(525) xor Codeword(607) xor Codeword(652) xor Codeword(696) xor
                Codeword(740) xor Codeword(808) xor Codeword(849) xor Codeword(926) xor
                Codeword(982) xor Codeword(1018) xor Codeword(1081) xor Codeword(1242) xor
                Codeword(1277) xor Codeword(1292) xor Codeword(1348) xor Codeword(1514) xor
                Codeword(1635) xor Codeword(1668) xor Codeword(1690) xor Codeword(1744) xor
                Codeword(1748) xor Codeword(1986) xor Codeword(2031) xor Codeword(2039);
 
     check367 <= Codeword(8) xor Codeword(110) xor Codeword(123) xor Codeword(205) xor
                Codeword(226) xor Codeword(320) xor Codeword(333) xor Codeword(397) xor
                Codeword(466) xor Codeword(520) xor Codeword(678) xor Codeword(799) xor
                Codeword(891) xor Codeword(945) xor Codeword(1010) xor Codeword(1087) xor
                Codeword(1149) xor Codeword(1241) xor Codeword(1300) xor Codeword(1380) xor
                Codeword(1494) xor Codeword(1589) xor Codeword(1611) xor Codeword(1694) xor
                Codeword(1734) xor Codeword(1735) xor Codeword(1749) xor Codeword(1800) xor
                Codeword(1857) xor Codeword(1919) xor Codeword(1934) xor Codeword(1950);
 
     check368 <= Codeword(7) xor Codeword(177) xor Codeword(381) xor Codeword(414) xor
                Codeword(496) xor Codeword(560) xor Codeword(580) xor Codeword(639) xor
                Codeword(685) xor Codeword(726) xor Codeword(822) xor Codeword(889) xor
                Codeword(946) xor Codeword(1026) xor Codeword(1143) xor Codeword(1180) xor
                Codeword(1296) xor Codeword(1372) xor Codeword(1467) xor Codeword(1545) xor
                Codeword(1641) xor Codeword(1714) xor Codeword(1787) xor Codeword(1837) xor
                Codeword(1859) xor Codeword(1907) xor Codeword(1916) xor Codeword(1940) xor
                Codeword(1952) xor Codeword(1989) xor Codeword(2040) xor Codeword(2046);
 
     check369 <= Codeword(6) xor Codeword(156) xor Codeword(221) xor Codeword(262) xor
                Codeword(358) xor Codeword(445) xor Codeword(450) xor Codeword(511) xor
                Codeword(594) xor Codeword(618) xor Codeword(708) xor Codeword(750) xor
                Codeword(827) xor Codeword(924) xor Codeword(981) xor Codeword(1030) xor
                Codeword(1125) xor Codeword(1166) xor Codeword(1183) xor Codeword(1255) xor
                Codeword(1335) xor Codeword(1422) xor Codeword(1570) xor Codeword(1585) xor
                Codeword(1612) xor Codeword(1670) xor Codeword(1715) xor Codeword(1917) xor
                Codeword(1998) xor Codeword(2008) xor Codeword(2017) xor Codeword(2030);
 
     check370 <= Codeword(5) xor Codeword(114) xor Codeword(208) xor Codeword(275) xor
                Codeword(341) xor Codeword(442) xor Codeword(500) xor Codeword(532) xor
                Codeword(635) xor Codeword(706) xor Codeword(732) xor Codeword(812) xor
                Codeword(843) xor Codeword(905) xor Codeword(973) xor Codeword(1103) xor
                Codeword(1110) xor Codeword(1132) xor Codeword(1257) xor Codeword(1291) xor
                Codeword(1393) xor Codeword(1435) xor Codeword(1505) xor Codeword(1518) xor
                Codeword(1603) xor Codeword(1745) xor Codeword(1757) xor Codeword(1778) xor
                Codeword(1826) xor Codeword(1910) xor Codeword(2033) xor Codeword(2036);
 
     check371 <= Codeword(4) xor Codeword(135) xor Codeword(173) xor Codeword(249) xor
                Codeword(354) xor Codeword(401) xor Codeword(504) xor Codeword(530) xor
                Codeword(563) xor Codeword(662) xor Codeword(683) xor Codeword(744) xor
                Codeword(814) xor Codeword(866) xor Codeword(908) xor Codeword(991) xor
                Codeword(1029) xor Codeword(1155) xor Codeword(1167) xor Codeword(1199) xor
                Codeword(1243) xor Codeword(1311) xor Codeword(1386) xor Codeword(1461) xor
                Codeword(1536) xor Codeword(1547) xor Codeword(1622) xor Codeword(1689) xor
                Codeword(1766) xor Codeword(1988) xor Codeword(2038) xor Codeword(2045);
 
     check372 <= Codeword(106) xor Codeword(144) xor Codeword(201) xor Codeword(229) xor
                Codeword(301) xor Codeword(365) xor Codeword(394) xor Codeword(493) xor
                Codeword(573) xor Codeword(648) xor Codeword(751) xor Codeword(878) xor
                Codeword(887) xor Codeword(892) xor Codeword(995) xor Codeword(1090) xor
                Codeword(1317) xor Codeword(1337) xor Codeword(1469) xor Codeword(1516) xor
                Codeword(1520) xor Codeword(1595) xor Codeword(1664) xor Codeword(1772) xor
                Codeword(1793) xor Codeword(1937) xor Codeword(1985) xor Codeword(2010) xor
                Codeword(2023) xor Codeword(2024) xor Codeword(2037) xor Codeword(2044);
 
     check373 <= Codeword(3) xor Codeword(139) xor Codeword(250) xor Codeword(310) xor
                Codeword(335) xor Codeword(425) xor Codeword(474) xor Codeword(546) xor
                Codeword(567) xor Codeword(620) xor Codeword(721) xor Codeword(725) xor
                Codeword(820) xor Codeword(875) xor Codeword(925) xor Codeword(1062) xor
                Codeword(1130) xor Codeword(1192) xor Codeword(1279) xor Codeword(1303) xor
                Codeword(1391) xor Codeword(1437) xor Codeword(1503) xor Codeword(1596) xor
                Codeword(1608) xor Codeword(1673) xor Codeword(1702) xor Codeword(1884) xor
                Codeword(1906) xor Codeword(1938) xor Codeword(1949) xor Codeword(1960);
 
     check374 <= Codeword(2) xor Codeword(85) xor Codeword(145) xor Codeword(213) xor
                Codeword(264) xor Codeword(306) xor Codeword(383) xor Codeword(436) xor
                Codeword(457) xor Codeword(549) xor Codeword(570) xor Codeword(709) xor
                Codeword(739) xor Codeword(778) xor Codeword(838) xor Codeword(888) xor
                Codeword(994) xor Codeword(1014) xor Codeword(1096) xor Codeword(1267) xor
                Codeword(1332) xor Codeword(1419) xor Codeword(1426) xor Codeword(1480) xor
                Codeword(1669) xor Codeword(1762) xor Codeword(1790) xor Codeword(1844) xor
                Codeword(1891) xor Codeword(1930) xor Codeword(1955) xor Codeword(1968);
 
     check375 <= Codeword(1) xor Codeword(64) xor Codeword(134) xor Codeword(260) xor
                Codeword(311) xor Codeword(368) xor Codeword(429) xor Codeword(469) xor
                Codeword(533) xor Codeword(615) xor Codeword(684) xor Codeword(768) xor
                Codeword(785) xor Codeword(860) xor Codeword(916) xor Codeword(989) xor
                Codeword(1035) xor Codeword(1107) xor Codeword(1114) xor Codeword(1201) xor
                Codeword(1218) xor Codeword(1252) xor Codeword(1377) xor Codeword(1416) xor
                Codeword(1442) xor Codeword(1526) xor Codeword(1602) xor Codeword(1636) xor
                Codeword(1652) xor Codeword(1848) xor Codeword(1854) xor Codeword(1903);
 
     check376 <= Codeword(0) xor Codeword(67) xor Codeword(159) xor Codeword(278) xor
                Codeword(386) xor Codeword(433) xor Codeword(479) xor Codeword(510) xor
                Codeword(595) xor Codeword(705) xor Codeword(746) xor Codeword(813) xor
                Codeword(861) xor Codeword(901) xor Codeword(970) xor Codeword(1063) xor
                Codeword(1156) xor Codeword(1220) xor Codeword(1334) xor Codeword(1343) xor
                Codeword(1465) xor Codeword(1522) xor Codeword(1539) xor Codeword(1629) xor
                Codeword(1659) xor Codeword(1838) xor Codeword(1886) xor Codeword(1912) xor
                Codeword(1939) xor Codeword(1948) xor Codeword(1954) xor Codeword(1971);
 
     check377 <= Codeword(107) xor Codeword(166) xor Codeword(193) xor Codeword(325) xor
                Codeword(347) xor Codeword(423) xor Codeword(451) xor Codeword(529) xor
                Codeword(579) xor Codeword(644) xor Codeword(676) xor Codeword(769) xor
                Codeword(837) xor Codeword(978) xor Codeword(1013) xor Codeword(1131) xor
                Codeword(1181) xor Codeword(1269) xor Codeword(1321) xor Codeword(1341) xor
                Codeword(1424) xor Codeword(1445) xor Codeword(1481) xor Codeword(1574) xor
                Codeword(1644) xor Codeword(1654) xor Codeword(1697) xor Codeword(1723) xor
                Codeword(1758) xor Codeword(1851) xor Codeword(1861) xor Codeword(1904);
 
     check378 <= Codeword(86) xor Codeword(149) xor Codeword(187) xor Codeword(246) xor
                Codeword(331) xor Codeword(355) xor Codeword(402) xor Codeword(495) xor
                Codeword(558) xor Codeword(591) xor Codeword(641) xor Codeword(716) xor
                Codeword(727) xor Codeword(800) xor Codeword(885) xor Codeword(918) xor
                Codeword(1000) xor Codeword(1049) xor Codeword(1102) xor Codeword(1153) xor
                Codeword(1198) xor Codeword(1256) xor Codeword(1375) xor Codeword(1399) xor
                Codeword(1430) xor Codeword(1488) xor Codeword(1527) xor Codeword(1553) xor
                Codeword(1657) xor Codeword(1709) xor Codeword(1923) xor Codeword(1928);
 
     check379 <= Codeword(105) xor Codeword(151) xor Codeword(277) xor Codeword(315) xor
                Codeword(351) xor Codeword(441) xor Codeword(482) xor Codeword(542) xor
                Codeword(655) xor Codeword(686) xor Codeword(724) xor Codeword(780) xor
                Codeword(847) xor Codeword(906) xor Codeword(999) xor Codeword(1052) xor
                Codeword(1079) xor Codeword(1122) xor Codeword(1174) xor Codeword(1275) xor
                Codeword(1356) xor Codeword(1388) xor Codeword(1410) xor Codeword(1460) xor
                Codeword(1555) xor Codeword(1648) xor Codeword(1716) xor Codeword(1722) xor
                Codeword(1777) xor Codeword(1880) xor Codeword(1979) xor Codeword(1984);
 
     check380 <= Codeword(77) xor Codeword(118) xor Codeword(182) xor Codeword(270) xor
                Codeword(317) xor Codeword(356) xor Codeword(398) xor Codeword(498) xor
                Codeword(512) xor Codeword(574) xor Codeword(650) xor Codeword(677) xor
                Codeword(742) xor Codeword(801) xor Codeword(852) xor Codeword(923) xor
                Codeword(976) xor Codeword(1036) xor Codeword(1171) xor Codeword(1248) xor
                Codeword(1316) xor Codeword(1358) xor Codeword(1403) xor Codeword(1446) xor
                Codeword(1507) xor Codeword(1510) xor Codeword(1559) xor Codeword(1587) xor
                Codeword(1674) xor Codeword(1713) xor Codeword(1721) xor Codeword(1808);
 
     check381 <= Codeword(60) xor Codeword(157) xor Codeword(214) xor Codeword(233) xor
                Codeword(287) xor Codeword(346) xor Codeword(408) xor Codeword(463) xor
                Codeword(559) xor Codeword(562) xor Codeword(719) xor Codeword(815) xor
                Codeword(897) xor Codeword(955) xor Codeword(1133) xor Codeword(1219) xor
                Codeword(1245) xor Codeword(1344) xor Codeword(1407) xor Codeword(1476) xor
                Codeword(1501) xor Codeword(1568) xor Codeword(1643) xor Codeword(1695) xor
                Codeword(1719) xor Codeword(1729) xor Codeword(1751) xor Codeword(1779) xor
                Codeword(1781) xor Codeword(1849) xor Codeword(1855) xor Codeword(1905);
 
     check382 <= Codeword(87) xor Codeword(111) xor Codeword(198) xor Codeword(237) xor
                Codeword(323) xor Codeword(371) xor Codeword(437) xor Codeword(471) xor
                Codeword(547) xor Codeword(603) xor Codeword(633) xor Codeword(682) xor
                Codeword(764) xor Codeword(811) xor Codeword(851) xor Codeword(894) xor
                Codeword(958) xor Codeword(1033) xor Codeword(1091) xor Codeword(1124) xor
                Codeword(1178) xor Codeword(1260) xor Codeword(1324) xor Codeword(1331) xor
                Codeword(1376) xor Codeword(1396) xor Codeword(1562) xor Codeword(1588) xor
                Codeword(1628) xor Codeword(1708) xor Codeword(1720) xor Codeword(1809);
 
     check383 <= Codeword(52) xor Codeword(79) xor Codeword(119) xor Codeword(209) xor
                Codeword(279) xor Codeword(282) xor Codeword(378) xor Codeword(424) xor
                Codeword(509) xor Codeword(565) xor Codeword(628) xor Codeword(713) xor
                Codeword(741) xor Codeword(829) xor Codeword(845) xor Codeword(910) xor
                Codeword(1001) xor Codeword(1003) xor Codeword(1089) xor Codeword(1209) xor
                Codeword(1254) xor Codeword(1294) xor Codeword(1340) xor Codeword(1513) xor
                Codeword(1565) xor Codeword(1597) xor Codeword(1633) xor Codeword(1680) xor
                Codeword(1750) xor Codeword(1775) xor Codeword(1882) xor Codeword(1914);
            else
                check0 <= '1';
            end if;
        end if;
    end process;
    check <=     check0 or 
    check1 or    check2 or    check3 or    check4 or    check5 or    check6 or    check7 or    check8 or 
    check9 or    check10 or    check11 or    check12 or    check13 or    check14 or    check15 or    check16 or 
    check17 or    check18 or    check19 or    check20 or    check21 or    check22 or    check23 or    check24 or 
    check25 or    check26 or    check27 or    check28 or    check29 or    check30 or    check31 or    check32 or 
    check33 or    check34 or    check35 or    check36 or    check37 or    check38 or    check39 or    check40 or 
    check41 or    check42 or    check43 or    check44 or    check45 or    check46 or    check47 or    check48 or 
    check49 or    check50 or    check51 or    check52 or    check53 or    check54 or    check55 or    check56 or 
    check57 or    check58 or    check59 or    check60 or    check61 or    check62 or    check63 or    check64 or 
    check65 or    check66 or    check67 or    check68 or    check69 or    check70 or    check71 or    check72 or 
    check73 or    check74 or    check75 or    check76 or    check77 or    check78 or    check79 or    check80 or 
    check81 or    check82 or    check83 or    check84 or    check85 or    check86 or    check87 or    check88 or 
    check89 or    check90 or    check91 or    check92 or    check93 or    check94 or    check95 or    check96 or 
    check97 or    check98 or    check99 or    check100 or    check101 or    check102 or    check103 or    check104 or 
    check105 or    check106 or    check107 or    check108 or    check109 or    check110 or    check111 or    check112 or 
    check113 or    check114 or    check115 or    check116 or    check117 or    check118 or    check119 or    check120 or 
    check121 or    check122 or    check123 or    check124 or    check125 or    check126 or    check127 or    check128 or 
    check129 or    check130 or    check131 or    check132 or    check133 or    check134 or    check135 or    check136 or 
    check137 or    check138 or    check139 or    check140 or    check141 or    check142 or    check143 or    check144 or 
    check145 or    check146 or    check147 or    check148 or    check149 or    check150 or    check151 or    check152 or 
    check153 or    check154 or    check155 or    check156 or    check157 or    check158 or    check159 or    check160 or 
    check161 or    check162 or    check163 or    check164 or    check165 or    check166 or    check167 or    check168 or 
    check169 or    check170 or    check171 or    check172 or    check173 or    check174 or    check175 or    check176 or 
    check177 or    check178 or    check179 or    check180 or    check181 or    check182 or    check183 or    check184 or 
    check185 or    check186 or    check187 or    check188 or    check189 or    check190 or    check191 or    check192 or 
    check193 or    check194 or    check195 or    check196 or    check197 or    check198 or    check199 or    check200 or 
    check201 or    check202 or    check203 or    check204 or    check205 or    check206 or    check207 or    check208 or 
    check209 or    check210 or    check211 or    check212 or    check213 or    check214 or    check215 or    check216 or 
    check217 or    check218 or    check219 or    check220 or    check221 or    check222 or    check223 or    check224 or 
    check225 or    check226 or    check227 or    check228 or    check229 or    check230 or    check231 or    check232 or 
    check233 or    check234 or    check235 or    check236 or    check237 or    check238 or    check239 or    check240 or 
    check241 or    check242 or    check243 or    check244 or    check245 or    check246 or    check247 or    check248 or 
    check249 or    check250 or    check251 or    check252 or    check253 or    check254 or    check255 or    check256 or 
    check257 or    check258 or    check259 or    check260 or    check261 or    check262 or    check263 or    check264 or 
    check265 or    check266 or    check267 or    check268 or    check269 or    check270 or    check271 or    check272 or 
    check273 or    check274 or    check275 or    check276 or    check277 or    check278 or    check279 or    check280 or 
    check281 or    check282 or    check283 or    check284 or    check285 or    check286 or    check287 or    check288 or 
    check289 or    check290 or    check291 or    check292 or    check293 or    check294 or    check295 or    check296 or 
    check297 or    check298 or    check299 or    check300 or    check301 or    check302 or    check303 or    check304 or 
    check305 or    check306 or    check307 or    check308 or    check309 or    check310 or    check311 or    check312 or 
    check313 or    check314 or    check315 or    check316 or    check317 or    check318 or    check319 or    check320 or 
    check321 or    check322 or    check323 or    check324 or    check325 or    check326 or    check327 or    check328 or 
    check329 or    check330 or    check331 or    check332 or    check333 or    check334 or    check335 or    check336 or 
    check337 or    check338 or    check339 or    check340 or    check341 or    check342 or    check343 or    check344 or 
    check345 or    check346 or    check347 or    check348 or    check349 or    check350 or    check351 or    check352 or 
    check353 or    check354 or    check355 or    check356 or    check357 or    check358 or    check359 or    check360 or 
    check361 or    check362 or    check363 or    check364 or    check365 or    check366 or    check367 or    check368 or 
    check369 or    check370 or    check371 or    check372 or    check373 or    check374 or    check375 or    check376 or 
    check377 or    check378 or    check379 or    check380 or    check381 or    check382 or    check383 ;
   

    early_stop : process(clk)
    begin
        if ( clk'event and clk = '1') then
            if( unsigned(Iterations) = 20 or check = '0' ) then        
                DecoderOver <= '1';                                                                      
            else
                DecoderOver <= '0';
            end if;
        end if;
    end process;

end architecture ; -- arch