library ieee;
use ieee.std_logic_1164.all;

entity CNUpdate is
  port (
    rst_n : in std_logic;
    clk : in std_logic;
    CN_sign_in : in std_logic_vector( 12287 downto 0 ); -- 384 * 32 = 12288
    CN_data_in : in std_logic_vector( 12287 downto 0 );
    CN_sign_out : out std_logic_vector( 12287 downto 0 );
    CN_data_out : out std_logic_vector( 12287 downto 0 )
  ) ;
end CNUpdate ;

architecture arch of CNUpdate is
    signal CN_sign_temp : std_logic_vector( 12287 downto 0 );
    signal CN_data_temp : std_logic_vector( 12287 downto 0 );
    
    component CN_Dv32 is
        port(
            VN2CN_bit  : in std_logic_vector( 31 downto 0 );
            VN2CN_sign : in std_logic_vector( 31 downto 0 );
            CN2VN_bit  : out std_logic_vector( 31 downto 0 );
            CN2VN_sign : out std_logic_vector( 31 downto 0)
        );
    end component;


begin
    process(clk, rst_n)
    begin
        if( rst_n = '0' ) then
            CN_sign_out <= ( others => '0' );
            CN_data_out <= ( others => '0' );
        elsif clk'event and clk = '1' then
            CN_sign_out <= CN_sign_temp;
            CN_data_out <= CN_data_temp;
        end if;
    end process;

    -- all CN update at the same time 384
    CN0 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 31 downto 0 ) ,
        VN2CN_bit   => CN_data_in( 31 downto 0 ) ,
        CN2VN_sign  => CN_sign_temp( 31 downto 0),
        CN2VN_bit   => CN_data_temp( 31 downto 0)
    );
    CN1 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 63 downto 32 ) ,
        VN2CN_bit   => CN_data_in( 63 downto 32 ) ,
        CN2VN_sign  => CN_sign_temp( 63 downto 32),
        CN2VN_bit   => CN_data_temp( 63 downto 32)
    );
    CN2 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 95 downto 64 ) ,
        VN2CN_bit   => CN_data_in( 95 downto 64 ) ,
        CN2VN_sign  => CN_sign_temp( 95 downto 64),
        CN2VN_bit   => CN_data_temp( 95 downto 64)
    );
    CN3 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 127 downto 96 ) ,
        VN2CN_bit   => CN_data_in( 127 downto 96 ) ,
        CN2VN_sign  => CN_sign_temp( 127 downto 96),
        CN2VN_bit   => CN_data_temp( 127 downto 96)
    );
    CN4 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 159 downto 128 ) ,
        VN2CN_bit   => CN_data_in( 159 downto 128 ) ,
        CN2VN_sign  => CN_sign_temp( 159 downto 128),
        CN2VN_bit   => CN_data_temp( 159 downto 128)
    );
    CN5 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 191 downto 160 ) ,
        VN2CN_bit   => CN_data_in( 191 downto 160 ) ,
        CN2VN_sign  => CN_sign_temp( 191 downto 160),
        CN2VN_bit   => CN_data_temp( 191 downto 160)
    );
    CN6 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 223 downto 192 ) ,
        VN2CN_bit   => CN_data_in( 223 downto 192 ) ,
        CN2VN_sign  => CN_sign_temp( 223 downto 192),
        CN2VN_bit   => CN_data_temp( 223 downto 192)
    );
    CN7 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 255 downto 224 ) ,
        VN2CN_bit   => CN_data_in( 255 downto 224 ) ,
        CN2VN_sign  => CN_sign_temp( 255 downto 224),
        CN2VN_bit   => CN_data_temp( 255 downto 224)
    );
    CN8 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 287 downto 256 ) ,
        VN2CN_bit   => CN_data_in( 287 downto 256 ) ,
        CN2VN_sign  => CN_sign_temp( 287 downto 256),
        CN2VN_bit   => CN_data_temp( 287 downto 256)
    );
    CN9 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 319 downto 288 ) ,
        VN2CN_bit   => CN_data_in( 319 downto 288 ) ,
        CN2VN_sign  => CN_sign_temp( 319 downto 288),
        CN2VN_bit   => CN_data_temp( 319 downto 288)
    );
    CN10 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 351 downto 320 ) ,
        VN2CN_bit   => CN_data_in( 351 downto 320 ) ,
        CN2VN_sign  => CN_sign_temp( 351 downto 320),
        CN2VN_bit   => CN_data_temp( 351 downto 320)
    );
    CN11 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 383 downto 352 ) ,
        VN2CN_bit   => CN_data_in( 383 downto 352 ) ,
        CN2VN_sign  => CN_sign_temp( 383 downto 352),
        CN2VN_bit   => CN_data_temp( 383 downto 352)
    );
    CN12 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 415 downto 384 ) ,
        VN2CN_bit   => CN_data_in( 415 downto 384 ) ,
        CN2VN_sign  => CN_sign_temp( 415 downto 384),
        CN2VN_bit   => CN_data_temp( 415 downto 384)
    );
    CN13 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 447 downto 416 ) ,
        VN2CN_bit   => CN_data_in( 447 downto 416 ) ,
        CN2VN_sign  => CN_sign_temp( 447 downto 416),
        CN2VN_bit   => CN_data_temp( 447 downto 416)
    );
    CN14 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 479 downto 448 ) ,
        VN2CN_bit   => CN_data_in( 479 downto 448 ) ,
        CN2VN_sign  => CN_sign_temp( 479 downto 448),
        CN2VN_bit   => CN_data_temp( 479 downto 448)
    );
    CN15 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 511 downto 480 ) ,
        VN2CN_bit   => CN_data_in( 511 downto 480 ) ,
        CN2VN_sign  => CN_sign_temp( 511 downto 480),
        CN2VN_bit   => CN_data_temp( 511 downto 480)
    );
    CN16 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 543 downto 512 ) ,
        VN2CN_bit   => CN_data_in( 543 downto 512 ) ,
        CN2VN_sign  => CN_sign_temp( 543 downto 512),
        CN2VN_bit   => CN_data_temp( 543 downto 512)
    );
    CN17 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 575 downto 544 ) ,
        VN2CN_bit   => CN_data_in( 575 downto 544 ) ,
        CN2VN_sign  => CN_sign_temp( 575 downto 544),
        CN2VN_bit   => CN_data_temp( 575 downto 544)
    );
    CN18 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 607 downto 576 ) ,
        VN2CN_bit   => CN_data_in( 607 downto 576 ) ,
        CN2VN_sign  => CN_sign_temp( 607 downto 576),
        CN2VN_bit   => CN_data_temp( 607 downto 576)
    );
    CN19 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 639 downto 608 ) ,
        VN2CN_bit   => CN_data_in( 639 downto 608 ) ,
        CN2VN_sign  => CN_sign_temp( 639 downto 608),
        CN2VN_bit   => CN_data_temp( 639 downto 608)
    );
    CN20 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 671 downto 640 ) ,
        VN2CN_bit   => CN_data_in( 671 downto 640 ) ,
        CN2VN_sign  => CN_sign_temp( 671 downto 640),
        CN2VN_bit   => CN_data_temp( 671 downto 640)
    );
    CN21 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 703 downto 672 ) ,
        VN2CN_bit   => CN_data_in( 703 downto 672 ) ,
        CN2VN_sign  => CN_sign_temp( 703 downto 672),
        CN2VN_bit   => CN_data_temp( 703 downto 672)
    );
    CN22 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 735 downto 704 ) ,
        VN2CN_bit   => CN_data_in( 735 downto 704 ) ,
        CN2VN_sign  => CN_sign_temp( 735 downto 704),
        CN2VN_bit   => CN_data_temp( 735 downto 704)
    );
    CN23 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 767 downto 736 ) ,
        VN2CN_bit   => CN_data_in( 767 downto 736 ) ,
        CN2VN_sign  => CN_sign_temp( 767 downto 736),
        CN2VN_bit   => CN_data_temp( 767 downto 736)
    );
    CN24 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 799 downto 768 ) ,
        VN2CN_bit   => CN_data_in( 799 downto 768 ) ,
        CN2VN_sign  => CN_sign_temp( 799 downto 768),
        CN2VN_bit   => CN_data_temp( 799 downto 768)
    );
    CN25 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 831 downto 800 ) ,
        VN2CN_bit   => CN_data_in( 831 downto 800 ) ,
        CN2VN_sign  => CN_sign_temp( 831 downto 800),
        CN2VN_bit   => CN_data_temp( 831 downto 800)
    );
    CN26 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 863 downto 832 ) ,
        VN2CN_bit   => CN_data_in( 863 downto 832 ) ,
        CN2VN_sign  => CN_sign_temp( 863 downto 832),
        CN2VN_bit   => CN_data_temp( 863 downto 832)
    );
    CN27 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 895 downto 864 ) ,
        VN2CN_bit   => CN_data_in( 895 downto 864 ) ,
        CN2VN_sign  => CN_sign_temp( 895 downto 864),
        CN2VN_bit   => CN_data_temp( 895 downto 864)
    );
    CN28 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 927 downto 896 ) ,
        VN2CN_bit   => CN_data_in( 927 downto 896 ) ,
        CN2VN_sign  => CN_sign_temp( 927 downto 896),
        CN2VN_bit   => CN_data_temp( 927 downto 896)
    );
    CN29 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 959 downto 928 ) ,
        VN2CN_bit   => CN_data_in( 959 downto 928 ) ,
        CN2VN_sign  => CN_sign_temp( 959 downto 928),
        CN2VN_bit   => CN_data_temp( 959 downto 928)
    );
    CN30 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 991 downto 960 ) ,
        VN2CN_bit   => CN_data_in( 991 downto 960 ) ,
        CN2VN_sign  => CN_sign_temp( 991 downto 960),
        CN2VN_bit   => CN_data_temp( 991 downto 960)
    );
    CN31 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1023 downto 992 ) ,
        VN2CN_bit   => CN_data_in( 1023 downto 992 ) ,
        CN2VN_sign  => CN_sign_temp( 1023 downto 992),
        CN2VN_bit   => CN_data_temp( 1023 downto 992)
    );
    CN32 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1055 downto 1024 ) ,
        VN2CN_bit   => CN_data_in( 1055 downto 1024 ) ,
        CN2VN_sign  => CN_sign_temp( 1055 downto 1024),
        CN2VN_bit   => CN_data_temp( 1055 downto 1024)
    );
    CN33 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1087 downto 1056 ) ,
        VN2CN_bit   => CN_data_in( 1087 downto 1056 ) ,
        CN2VN_sign  => CN_sign_temp( 1087 downto 1056),
        CN2VN_bit   => CN_data_temp( 1087 downto 1056)
    );
    CN34 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1119 downto 1088 ) ,
        VN2CN_bit   => CN_data_in( 1119 downto 1088 ) ,
        CN2VN_sign  => CN_sign_temp( 1119 downto 1088),
        CN2VN_bit   => CN_data_temp( 1119 downto 1088)
    );
    CN35 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1151 downto 1120 ) ,
        VN2CN_bit   => CN_data_in( 1151 downto 1120 ) ,
        CN2VN_sign  => CN_sign_temp( 1151 downto 1120),
        CN2VN_bit   => CN_data_temp( 1151 downto 1120)
    );
    CN36 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1183 downto 1152 ) ,
        VN2CN_bit   => CN_data_in( 1183 downto 1152 ) ,
        CN2VN_sign  => CN_sign_temp( 1183 downto 1152),
        CN2VN_bit   => CN_data_temp( 1183 downto 1152)
    );
    CN37 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1215 downto 1184 ) ,
        VN2CN_bit   => CN_data_in( 1215 downto 1184 ) ,
        CN2VN_sign  => CN_sign_temp( 1215 downto 1184),
        CN2VN_bit   => CN_data_temp( 1215 downto 1184)
    );
    CN38 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1247 downto 1216 ) ,
        VN2CN_bit   => CN_data_in( 1247 downto 1216 ) ,
        CN2VN_sign  => CN_sign_temp( 1247 downto 1216),
        CN2VN_bit   => CN_data_temp( 1247 downto 1216)
    );
    CN39 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1279 downto 1248 ) ,
        VN2CN_bit   => CN_data_in( 1279 downto 1248 ) ,
        CN2VN_sign  => CN_sign_temp( 1279 downto 1248),
        CN2VN_bit   => CN_data_temp( 1279 downto 1248)
    );
    CN40 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1311 downto 1280 ) ,
        VN2CN_bit   => CN_data_in( 1311 downto 1280 ) ,
        CN2VN_sign  => CN_sign_temp( 1311 downto 1280),
        CN2VN_bit   => CN_data_temp( 1311 downto 1280)
    );
    CN41 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1343 downto 1312 ) ,
        VN2CN_bit   => CN_data_in( 1343 downto 1312 ) ,
        CN2VN_sign  => CN_sign_temp( 1343 downto 1312),
        CN2VN_bit   => CN_data_temp( 1343 downto 1312)
    );
    CN42 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1375 downto 1344 ) ,
        VN2CN_bit   => CN_data_in( 1375 downto 1344 ) ,
        CN2VN_sign  => CN_sign_temp( 1375 downto 1344),
        CN2VN_bit   => CN_data_temp( 1375 downto 1344)
    );
    CN43 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1407 downto 1376 ) ,
        VN2CN_bit   => CN_data_in( 1407 downto 1376 ) ,
        CN2VN_sign  => CN_sign_temp( 1407 downto 1376),
        CN2VN_bit   => CN_data_temp( 1407 downto 1376)
    );
    CN44 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1439 downto 1408 ) ,
        VN2CN_bit   => CN_data_in( 1439 downto 1408 ) ,
        CN2VN_sign  => CN_sign_temp( 1439 downto 1408),
        CN2VN_bit   => CN_data_temp( 1439 downto 1408)
    );
    CN45 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1471 downto 1440 ) ,
        VN2CN_bit   => CN_data_in( 1471 downto 1440 ) ,
        CN2VN_sign  => CN_sign_temp( 1471 downto 1440),
        CN2VN_bit   => CN_data_temp( 1471 downto 1440)
    );
    CN46 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1503 downto 1472 ) ,
        VN2CN_bit   => CN_data_in( 1503 downto 1472 ) ,
        CN2VN_sign  => CN_sign_temp( 1503 downto 1472),
        CN2VN_bit   => CN_data_temp( 1503 downto 1472)
    );
    CN47 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1535 downto 1504 ) ,
        VN2CN_bit   => CN_data_in( 1535 downto 1504 ) ,
        CN2VN_sign  => CN_sign_temp( 1535 downto 1504),
        CN2VN_bit   => CN_data_temp( 1535 downto 1504)
    );
    CN48 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1567 downto 1536 ) ,
        VN2CN_bit   => CN_data_in( 1567 downto 1536 ) ,
        CN2VN_sign  => CN_sign_temp( 1567 downto 1536),
        CN2VN_bit   => CN_data_temp( 1567 downto 1536)
    );
    CN49 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1599 downto 1568 ) ,
        VN2CN_bit   => CN_data_in( 1599 downto 1568 ) ,
        CN2VN_sign  => CN_sign_temp( 1599 downto 1568),
        CN2VN_bit   => CN_data_temp( 1599 downto 1568)
    );
    CN50 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1631 downto 1600 ) ,
        VN2CN_bit   => CN_data_in( 1631 downto 1600 ) ,
        CN2VN_sign  => CN_sign_temp( 1631 downto 1600),
        CN2VN_bit   => CN_data_temp( 1631 downto 1600)
    );
    CN51 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1663 downto 1632 ) ,
        VN2CN_bit   => CN_data_in( 1663 downto 1632 ) ,
        CN2VN_sign  => CN_sign_temp( 1663 downto 1632),
        CN2VN_bit   => CN_data_temp( 1663 downto 1632)
    );
    CN52 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1695 downto 1664 ) ,
        VN2CN_bit   => CN_data_in( 1695 downto 1664 ) ,
        CN2VN_sign  => CN_sign_temp( 1695 downto 1664),
        CN2VN_bit   => CN_data_temp( 1695 downto 1664)
    );
    CN53 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1727 downto 1696 ) ,
        VN2CN_bit   => CN_data_in( 1727 downto 1696 ) ,
        CN2VN_sign  => CN_sign_temp( 1727 downto 1696),
        CN2VN_bit   => CN_data_temp( 1727 downto 1696)
    );
    CN54 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1759 downto 1728 ) ,
        VN2CN_bit   => CN_data_in( 1759 downto 1728 ) ,
        CN2VN_sign  => CN_sign_temp( 1759 downto 1728),
        CN2VN_bit   => CN_data_temp( 1759 downto 1728)
    );
    CN55 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1791 downto 1760 ) ,
        VN2CN_bit   => CN_data_in( 1791 downto 1760 ) ,
        CN2VN_sign  => CN_sign_temp( 1791 downto 1760),
        CN2VN_bit   => CN_data_temp( 1791 downto 1760)
    );
    CN56 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1823 downto 1792 ) ,
        VN2CN_bit   => CN_data_in( 1823 downto 1792 ) ,
        CN2VN_sign  => CN_sign_temp( 1823 downto 1792),
        CN2VN_bit   => CN_data_temp( 1823 downto 1792)
    );
    CN57 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1855 downto 1824 ) ,
        VN2CN_bit   => CN_data_in( 1855 downto 1824 ) ,
        CN2VN_sign  => CN_sign_temp( 1855 downto 1824),
        CN2VN_bit   => CN_data_temp( 1855 downto 1824)
    );
    CN58 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1887 downto 1856 ) ,
        VN2CN_bit   => CN_data_in( 1887 downto 1856 ) ,
        CN2VN_sign  => CN_sign_temp( 1887 downto 1856),
        CN2VN_bit   => CN_data_temp( 1887 downto 1856)
    );
    CN59 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1919 downto 1888 ) ,
        VN2CN_bit   => CN_data_in( 1919 downto 1888 ) ,
        CN2VN_sign  => CN_sign_temp( 1919 downto 1888),
        CN2VN_bit   => CN_data_temp( 1919 downto 1888)
    );
    CN60 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1951 downto 1920 ) ,
        VN2CN_bit   => CN_data_in( 1951 downto 1920 ) ,
        CN2VN_sign  => CN_sign_temp( 1951 downto 1920),
        CN2VN_bit   => CN_data_temp( 1951 downto 1920)
    );
    CN61 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 1983 downto 1952 ) ,
        VN2CN_bit   => CN_data_in( 1983 downto 1952 ) ,
        CN2VN_sign  => CN_sign_temp( 1983 downto 1952),
        CN2VN_bit   => CN_data_temp( 1983 downto 1952)
    );
    CN62 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2015 downto 1984 ) ,
        VN2CN_bit   => CN_data_in( 2015 downto 1984 ) ,
        CN2VN_sign  => CN_sign_temp( 2015 downto 1984),
        CN2VN_bit   => CN_data_temp( 2015 downto 1984)
    );
    CN63 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2047 downto 2016 ) ,
        VN2CN_bit   => CN_data_in( 2047 downto 2016 ) ,
        CN2VN_sign  => CN_sign_temp( 2047 downto 2016),
        CN2VN_bit   => CN_data_temp( 2047 downto 2016)
    );
    CN64 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2079 downto 2048 ) ,
        VN2CN_bit   => CN_data_in( 2079 downto 2048 ) ,
        CN2VN_sign  => CN_sign_temp( 2079 downto 2048),
        CN2VN_bit   => CN_data_temp( 2079 downto 2048)
    );
    CN65 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2111 downto 2080 ) ,
        VN2CN_bit   => CN_data_in( 2111 downto 2080 ) ,
        CN2VN_sign  => CN_sign_temp( 2111 downto 2080),
        CN2VN_bit   => CN_data_temp( 2111 downto 2080)
    );
    CN66 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2143 downto 2112 ) ,
        VN2CN_bit   => CN_data_in( 2143 downto 2112 ) ,
        CN2VN_sign  => CN_sign_temp( 2143 downto 2112),
        CN2VN_bit   => CN_data_temp( 2143 downto 2112)
    );
    CN67 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2175 downto 2144 ) ,
        VN2CN_bit   => CN_data_in( 2175 downto 2144 ) ,
        CN2VN_sign  => CN_sign_temp( 2175 downto 2144),
        CN2VN_bit   => CN_data_temp( 2175 downto 2144)
    );
    CN68 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2207 downto 2176 ) ,
        VN2CN_bit   => CN_data_in( 2207 downto 2176 ) ,
        CN2VN_sign  => CN_sign_temp( 2207 downto 2176),
        CN2VN_bit   => CN_data_temp( 2207 downto 2176)
    );
    CN69 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2239 downto 2208 ) ,
        VN2CN_bit   => CN_data_in( 2239 downto 2208 ) ,
        CN2VN_sign  => CN_sign_temp( 2239 downto 2208),
        CN2VN_bit   => CN_data_temp( 2239 downto 2208)
    );
    CN70 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2271 downto 2240 ) ,
        VN2CN_bit   => CN_data_in( 2271 downto 2240 ) ,
        CN2VN_sign  => CN_sign_temp( 2271 downto 2240),
        CN2VN_bit   => CN_data_temp( 2271 downto 2240)
    );
    CN71 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2303 downto 2272 ) ,
        VN2CN_bit   => CN_data_in( 2303 downto 2272 ) ,
        CN2VN_sign  => CN_sign_temp( 2303 downto 2272),
        CN2VN_bit   => CN_data_temp( 2303 downto 2272)
    );
    CN72 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2335 downto 2304 ) ,
        VN2CN_bit   => CN_data_in( 2335 downto 2304 ) ,
        CN2VN_sign  => CN_sign_temp( 2335 downto 2304),
        CN2VN_bit   => CN_data_temp( 2335 downto 2304)
    );
    CN73 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2367 downto 2336 ) ,
        VN2CN_bit   => CN_data_in( 2367 downto 2336 ) ,
        CN2VN_sign  => CN_sign_temp( 2367 downto 2336),
        CN2VN_bit   => CN_data_temp( 2367 downto 2336)
    );
    CN74 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2399 downto 2368 ) ,
        VN2CN_bit   => CN_data_in( 2399 downto 2368 ) ,
        CN2VN_sign  => CN_sign_temp( 2399 downto 2368),
        CN2VN_bit   => CN_data_temp( 2399 downto 2368)
    );
    CN75 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2431 downto 2400 ) ,
        VN2CN_bit   => CN_data_in( 2431 downto 2400 ) ,
        CN2VN_sign  => CN_sign_temp( 2431 downto 2400),
        CN2VN_bit   => CN_data_temp( 2431 downto 2400)
    );
    CN76 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2463 downto 2432 ) ,
        VN2CN_bit   => CN_data_in( 2463 downto 2432 ) ,
        CN2VN_sign  => CN_sign_temp( 2463 downto 2432),
        CN2VN_bit   => CN_data_temp( 2463 downto 2432)
    );
    CN77 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2495 downto 2464 ) ,
        VN2CN_bit   => CN_data_in( 2495 downto 2464 ) ,
        CN2VN_sign  => CN_sign_temp( 2495 downto 2464),
        CN2VN_bit   => CN_data_temp( 2495 downto 2464)
    );
    CN78 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2527 downto 2496 ) ,
        VN2CN_bit   => CN_data_in( 2527 downto 2496 ) ,
        CN2VN_sign  => CN_sign_temp( 2527 downto 2496),
        CN2VN_bit   => CN_data_temp( 2527 downto 2496)
    );
    CN79 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2559 downto 2528 ) ,
        VN2CN_bit   => CN_data_in( 2559 downto 2528 ) ,
        CN2VN_sign  => CN_sign_temp( 2559 downto 2528),
        CN2VN_bit   => CN_data_temp( 2559 downto 2528)
    );
    CN80 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2591 downto 2560 ) ,
        VN2CN_bit   => CN_data_in( 2591 downto 2560 ) ,
        CN2VN_sign  => CN_sign_temp( 2591 downto 2560),
        CN2VN_bit   => CN_data_temp( 2591 downto 2560)
    );
    CN81 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2623 downto 2592 ) ,
        VN2CN_bit   => CN_data_in( 2623 downto 2592 ) ,
        CN2VN_sign  => CN_sign_temp( 2623 downto 2592),
        CN2VN_bit   => CN_data_temp( 2623 downto 2592)
    );
    CN82 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2655 downto 2624 ) ,
        VN2CN_bit   => CN_data_in( 2655 downto 2624 ) ,
        CN2VN_sign  => CN_sign_temp( 2655 downto 2624),
        CN2VN_bit   => CN_data_temp( 2655 downto 2624)
    );
    CN83 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2687 downto 2656 ) ,
        VN2CN_bit   => CN_data_in( 2687 downto 2656 ) ,
        CN2VN_sign  => CN_sign_temp( 2687 downto 2656),
        CN2VN_bit   => CN_data_temp( 2687 downto 2656)
    );
    CN84 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2719 downto 2688 ) ,
        VN2CN_bit   => CN_data_in( 2719 downto 2688 ) ,
        CN2VN_sign  => CN_sign_temp( 2719 downto 2688),
        CN2VN_bit   => CN_data_temp( 2719 downto 2688)
    );
    CN85 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2751 downto 2720 ) ,
        VN2CN_bit   => CN_data_in( 2751 downto 2720 ) ,
        CN2VN_sign  => CN_sign_temp( 2751 downto 2720),
        CN2VN_bit   => CN_data_temp( 2751 downto 2720)
    );
    CN86 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2783 downto 2752 ) ,
        VN2CN_bit   => CN_data_in( 2783 downto 2752 ) ,
        CN2VN_sign  => CN_sign_temp( 2783 downto 2752),
        CN2VN_bit   => CN_data_temp( 2783 downto 2752)
    );
    CN87 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2815 downto 2784 ) ,
        VN2CN_bit   => CN_data_in( 2815 downto 2784 ) ,
        CN2VN_sign  => CN_sign_temp( 2815 downto 2784),
        CN2VN_bit   => CN_data_temp( 2815 downto 2784)
    );
    CN88 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2847 downto 2816 ) ,
        VN2CN_bit   => CN_data_in( 2847 downto 2816 ) ,
        CN2VN_sign  => CN_sign_temp( 2847 downto 2816),
        CN2VN_bit   => CN_data_temp( 2847 downto 2816)
    );
    CN89 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2879 downto 2848 ) ,
        VN2CN_bit   => CN_data_in( 2879 downto 2848 ) ,
        CN2VN_sign  => CN_sign_temp( 2879 downto 2848),
        CN2VN_bit   => CN_data_temp( 2879 downto 2848)
    );
    CN90 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2911 downto 2880 ) ,
        VN2CN_bit   => CN_data_in( 2911 downto 2880 ) ,
        CN2VN_sign  => CN_sign_temp( 2911 downto 2880),
        CN2VN_bit   => CN_data_temp( 2911 downto 2880)
    );
    CN91 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2943 downto 2912 ) ,
        VN2CN_bit   => CN_data_in( 2943 downto 2912 ) ,
        CN2VN_sign  => CN_sign_temp( 2943 downto 2912),
        CN2VN_bit   => CN_data_temp( 2943 downto 2912)
    );
    CN92 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 2975 downto 2944 ) ,
        VN2CN_bit   => CN_data_in( 2975 downto 2944 ) ,
        CN2VN_sign  => CN_sign_temp( 2975 downto 2944),
        CN2VN_bit   => CN_data_temp( 2975 downto 2944)
    );
    CN93 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3007 downto 2976 ) ,
        VN2CN_bit   => CN_data_in( 3007 downto 2976 ) ,
        CN2VN_sign  => CN_sign_temp( 3007 downto 2976),
        CN2VN_bit   => CN_data_temp( 3007 downto 2976)
    );
    CN94 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3039 downto 3008 ) ,
        VN2CN_bit   => CN_data_in( 3039 downto 3008 ) ,
        CN2VN_sign  => CN_sign_temp( 3039 downto 3008),
        CN2VN_bit   => CN_data_temp( 3039 downto 3008)
    );
    CN95 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3071 downto 3040 ) ,
        VN2CN_bit   => CN_data_in( 3071 downto 3040 ) ,
        CN2VN_sign  => CN_sign_temp( 3071 downto 3040),
        CN2VN_bit   => CN_data_temp( 3071 downto 3040)
    );
    CN96 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3103 downto 3072 ) ,
        VN2CN_bit   => CN_data_in( 3103 downto 3072 ) ,
        CN2VN_sign  => CN_sign_temp( 3103 downto 3072),
        CN2VN_bit   => CN_data_temp( 3103 downto 3072)
    );
    CN97 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3135 downto 3104 ) ,
        VN2CN_bit   => CN_data_in( 3135 downto 3104 ) ,
        CN2VN_sign  => CN_sign_temp( 3135 downto 3104),
        CN2VN_bit   => CN_data_temp( 3135 downto 3104)
    );
    CN98 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3167 downto 3136 ) ,
        VN2CN_bit   => CN_data_in( 3167 downto 3136 ) ,
        CN2VN_sign  => CN_sign_temp( 3167 downto 3136),
        CN2VN_bit   => CN_data_temp( 3167 downto 3136)
    );
    CN99 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3199 downto 3168 ) ,
        VN2CN_bit   => CN_data_in( 3199 downto 3168 ) ,
        CN2VN_sign  => CN_sign_temp( 3199 downto 3168),
        CN2VN_bit   => CN_data_temp( 3199 downto 3168)
    );
    CN100 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3231 downto 3200 ) ,
        VN2CN_bit   => CN_data_in( 3231 downto 3200 ) ,
        CN2VN_sign  => CN_sign_temp( 3231 downto 3200),
        CN2VN_bit   => CN_data_temp( 3231 downto 3200)
    );
    CN101 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3263 downto 3232 ) ,
        VN2CN_bit   => CN_data_in( 3263 downto 3232 ) ,
        CN2VN_sign  => CN_sign_temp( 3263 downto 3232),
        CN2VN_bit   => CN_data_temp( 3263 downto 3232)
    );
    CN102 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3295 downto 3264 ) ,
        VN2CN_bit   => CN_data_in( 3295 downto 3264 ) ,
        CN2VN_sign  => CN_sign_temp( 3295 downto 3264),
        CN2VN_bit   => CN_data_temp( 3295 downto 3264)
    );
    CN103 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3327 downto 3296 ) ,
        VN2CN_bit   => CN_data_in( 3327 downto 3296 ) ,
        CN2VN_sign  => CN_sign_temp( 3327 downto 3296),
        CN2VN_bit   => CN_data_temp( 3327 downto 3296)
    );
    CN104 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3359 downto 3328 ) ,
        VN2CN_bit   => CN_data_in( 3359 downto 3328 ) ,
        CN2VN_sign  => CN_sign_temp( 3359 downto 3328),
        CN2VN_bit   => CN_data_temp( 3359 downto 3328)
    );
    CN105 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3391 downto 3360 ) ,
        VN2CN_bit   => CN_data_in( 3391 downto 3360 ) ,
        CN2VN_sign  => CN_sign_temp( 3391 downto 3360),
        CN2VN_bit   => CN_data_temp( 3391 downto 3360)
    );
    CN106 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3423 downto 3392 ) ,
        VN2CN_bit   => CN_data_in( 3423 downto 3392 ) ,
        CN2VN_sign  => CN_sign_temp( 3423 downto 3392),
        CN2VN_bit   => CN_data_temp( 3423 downto 3392)
    );
    CN107 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3455 downto 3424 ) ,
        VN2CN_bit   => CN_data_in( 3455 downto 3424 ) ,
        CN2VN_sign  => CN_sign_temp( 3455 downto 3424),
        CN2VN_bit   => CN_data_temp( 3455 downto 3424)
    );
    CN108 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3487 downto 3456 ) ,
        VN2CN_bit   => CN_data_in( 3487 downto 3456 ) ,
        CN2VN_sign  => CN_sign_temp( 3487 downto 3456),
        CN2VN_bit   => CN_data_temp( 3487 downto 3456)
    );
    CN109 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3519 downto 3488 ) ,
        VN2CN_bit   => CN_data_in( 3519 downto 3488 ) ,
        CN2VN_sign  => CN_sign_temp( 3519 downto 3488),
        CN2VN_bit   => CN_data_temp( 3519 downto 3488)
    );
    CN110 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3551 downto 3520 ) ,
        VN2CN_bit   => CN_data_in( 3551 downto 3520 ) ,
        CN2VN_sign  => CN_sign_temp( 3551 downto 3520),
        CN2VN_bit   => CN_data_temp( 3551 downto 3520)
    );
    CN111 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3583 downto 3552 ) ,
        VN2CN_bit   => CN_data_in( 3583 downto 3552 ) ,
        CN2VN_sign  => CN_sign_temp( 3583 downto 3552),
        CN2VN_bit   => CN_data_temp( 3583 downto 3552)
    );
    CN112 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3615 downto 3584 ) ,
        VN2CN_bit   => CN_data_in( 3615 downto 3584 ) ,
        CN2VN_sign  => CN_sign_temp( 3615 downto 3584),
        CN2VN_bit   => CN_data_temp( 3615 downto 3584)
    );
    CN113 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3647 downto 3616 ) ,
        VN2CN_bit   => CN_data_in( 3647 downto 3616 ) ,
        CN2VN_sign  => CN_sign_temp( 3647 downto 3616),
        CN2VN_bit   => CN_data_temp( 3647 downto 3616)
    );
    CN114 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3679 downto 3648 ) ,
        VN2CN_bit   => CN_data_in( 3679 downto 3648 ) ,
        CN2VN_sign  => CN_sign_temp( 3679 downto 3648),
        CN2VN_bit   => CN_data_temp( 3679 downto 3648)
    );
    CN115 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3711 downto 3680 ) ,
        VN2CN_bit   => CN_data_in( 3711 downto 3680 ) ,
        CN2VN_sign  => CN_sign_temp( 3711 downto 3680),
        CN2VN_bit   => CN_data_temp( 3711 downto 3680)
    );
    CN116 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3743 downto 3712 ) ,
        VN2CN_bit   => CN_data_in( 3743 downto 3712 ) ,
        CN2VN_sign  => CN_sign_temp( 3743 downto 3712),
        CN2VN_bit   => CN_data_temp( 3743 downto 3712)
    );
    CN117 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3775 downto 3744 ) ,
        VN2CN_bit   => CN_data_in( 3775 downto 3744 ) ,
        CN2VN_sign  => CN_sign_temp( 3775 downto 3744),
        CN2VN_bit   => CN_data_temp( 3775 downto 3744)
    );
    CN118 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3807 downto 3776 ) ,
        VN2CN_bit   => CN_data_in( 3807 downto 3776 ) ,
        CN2VN_sign  => CN_sign_temp( 3807 downto 3776),
        CN2VN_bit   => CN_data_temp( 3807 downto 3776)
    );
    CN119 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3839 downto 3808 ) ,
        VN2CN_bit   => CN_data_in( 3839 downto 3808 ) ,
        CN2VN_sign  => CN_sign_temp( 3839 downto 3808),
        CN2VN_bit   => CN_data_temp( 3839 downto 3808)
    );
    CN120 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3871 downto 3840 ) ,
        VN2CN_bit   => CN_data_in( 3871 downto 3840 ) ,
        CN2VN_sign  => CN_sign_temp( 3871 downto 3840),
        CN2VN_bit   => CN_data_temp( 3871 downto 3840)
    );
    CN121 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3903 downto 3872 ) ,
        VN2CN_bit   => CN_data_in( 3903 downto 3872 ) ,
        CN2VN_sign  => CN_sign_temp( 3903 downto 3872),
        CN2VN_bit   => CN_data_temp( 3903 downto 3872)
    );
    CN122 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3935 downto 3904 ) ,
        VN2CN_bit   => CN_data_in( 3935 downto 3904 ) ,
        CN2VN_sign  => CN_sign_temp( 3935 downto 3904),
        CN2VN_bit   => CN_data_temp( 3935 downto 3904)
    );
    CN123 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3967 downto 3936 ) ,
        VN2CN_bit   => CN_data_in( 3967 downto 3936 ) ,
        CN2VN_sign  => CN_sign_temp( 3967 downto 3936),
        CN2VN_bit   => CN_data_temp( 3967 downto 3936)
    );
    CN124 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 3999 downto 3968 ) ,
        VN2CN_bit   => CN_data_in( 3999 downto 3968 ) ,
        CN2VN_sign  => CN_sign_temp( 3999 downto 3968),
        CN2VN_bit   => CN_data_temp( 3999 downto 3968)
    );
    CN125 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4031 downto 4000 ) ,
        VN2CN_bit   => CN_data_in( 4031 downto 4000 ) ,
        CN2VN_sign  => CN_sign_temp( 4031 downto 4000),
        CN2VN_bit   => CN_data_temp( 4031 downto 4000)
    );
    CN126 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4063 downto 4032 ) ,
        VN2CN_bit   => CN_data_in( 4063 downto 4032 ) ,
        CN2VN_sign  => CN_sign_temp( 4063 downto 4032),
        CN2VN_bit   => CN_data_temp( 4063 downto 4032)
    );
    CN127 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4095 downto 4064 ) ,
        VN2CN_bit   => CN_data_in( 4095 downto 4064 ) ,
        CN2VN_sign  => CN_sign_temp( 4095 downto 4064),
        CN2VN_bit   => CN_data_temp( 4095 downto 4064)
    );
    CN128 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4127 downto 4096 ) ,
        VN2CN_bit   => CN_data_in( 4127 downto 4096 ) ,
        CN2VN_sign  => CN_sign_temp( 4127 downto 4096),
        CN2VN_bit   => CN_data_temp( 4127 downto 4096)
    );
    CN129 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4159 downto 4128 ) ,
        VN2CN_bit   => CN_data_in( 4159 downto 4128 ) ,
        CN2VN_sign  => CN_sign_temp( 4159 downto 4128),
        CN2VN_bit   => CN_data_temp( 4159 downto 4128)
    );
    CN130 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4191 downto 4160 ) ,
        VN2CN_bit   => CN_data_in( 4191 downto 4160 ) ,
        CN2VN_sign  => CN_sign_temp( 4191 downto 4160),
        CN2VN_bit   => CN_data_temp( 4191 downto 4160)
    );
    CN131 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4223 downto 4192 ) ,
        VN2CN_bit   => CN_data_in( 4223 downto 4192 ) ,
        CN2VN_sign  => CN_sign_temp( 4223 downto 4192),
        CN2VN_bit   => CN_data_temp( 4223 downto 4192)
    );
    CN132 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4255 downto 4224 ) ,
        VN2CN_bit   => CN_data_in( 4255 downto 4224 ) ,
        CN2VN_sign  => CN_sign_temp( 4255 downto 4224),
        CN2VN_bit   => CN_data_temp( 4255 downto 4224)
    );
    CN133 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4287 downto 4256 ) ,
        VN2CN_bit   => CN_data_in( 4287 downto 4256 ) ,
        CN2VN_sign  => CN_sign_temp( 4287 downto 4256),
        CN2VN_bit   => CN_data_temp( 4287 downto 4256)
    );
    CN134 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4319 downto 4288 ) ,
        VN2CN_bit   => CN_data_in( 4319 downto 4288 ) ,
        CN2VN_sign  => CN_sign_temp( 4319 downto 4288),
        CN2VN_bit   => CN_data_temp( 4319 downto 4288)
    );
    CN135 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4351 downto 4320 ) ,
        VN2CN_bit   => CN_data_in( 4351 downto 4320 ) ,
        CN2VN_sign  => CN_sign_temp( 4351 downto 4320),
        CN2VN_bit   => CN_data_temp( 4351 downto 4320)
    );
    CN136 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4383 downto 4352 ) ,
        VN2CN_bit   => CN_data_in( 4383 downto 4352 ) ,
        CN2VN_sign  => CN_sign_temp( 4383 downto 4352),
        CN2VN_bit   => CN_data_temp( 4383 downto 4352)
    );
    CN137 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4415 downto 4384 ) ,
        VN2CN_bit   => CN_data_in( 4415 downto 4384 ) ,
        CN2VN_sign  => CN_sign_temp( 4415 downto 4384),
        CN2VN_bit   => CN_data_temp( 4415 downto 4384)
    );
    CN138 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4447 downto 4416 ) ,
        VN2CN_bit   => CN_data_in( 4447 downto 4416 ) ,
        CN2VN_sign  => CN_sign_temp( 4447 downto 4416),
        CN2VN_bit   => CN_data_temp( 4447 downto 4416)
    );
    CN139 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4479 downto 4448 ) ,
        VN2CN_bit   => CN_data_in( 4479 downto 4448 ) ,
        CN2VN_sign  => CN_sign_temp( 4479 downto 4448),
        CN2VN_bit   => CN_data_temp( 4479 downto 4448)
    );
    CN140 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4511 downto 4480 ) ,
        VN2CN_bit   => CN_data_in( 4511 downto 4480 ) ,
        CN2VN_sign  => CN_sign_temp( 4511 downto 4480),
        CN2VN_bit   => CN_data_temp( 4511 downto 4480)
    );
    CN141 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4543 downto 4512 ) ,
        VN2CN_bit   => CN_data_in( 4543 downto 4512 ) ,
        CN2VN_sign  => CN_sign_temp( 4543 downto 4512),
        CN2VN_bit   => CN_data_temp( 4543 downto 4512)
    );
    CN142 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4575 downto 4544 ) ,
        VN2CN_bit   => CN_data_in( 4575 downto 4544 ) ,
        CN2VN_sign  => CN_sign_temp( 4575 downto 4544),
        CN2VN_bit   => CN_data_temp( 4575 downto 4544)
    );
    CN143 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4607 downto 4576 ) ,
        VN2CN_bit   => CN_data_in( 4607 downto 4576 ) ,
        CN2VN_sign  => CN_sign_temp( 4607 downto 4576),
        CN2VN_bit   => CN_data_temp( 4607 downto 4576)
    );
    CN144 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4639 downto 4608 ) ,
        VN2CN_bit   => CN_data_in( 4639 downto 4608 ) ,
        CN2VN_sign  => CN_sign_temp( 4639 downto 4608),
        CN2VN_bit   => CN_data_temp( 4639 downto 4608)
    );
    CN145 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4671 downto 4640 ) ,
        VN2CN_bit   => CN_data_in( 4671 downto 4640 ) ,
        CN2VN_sign  => CN_sign_temp( 4671 downto 4640),
        CN2VN_bit   => CN_data_temp( 4671 downto 4640)
    );
    CN146 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4703 downto 4672 ) ,
        VN2CN_bit   => CN_data_in( 4703 downto 4672 ) ,
        CN2VN_sign  => CN_sign_temp( 4703 downto 4672),
        CN2VN_bit   => CN_data_temp( 4703 downto 4672)
    );
    CN147 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4735 downto 4704 ) ,
        VN2CN_bit   => CN_data_in( 4735 downto 4704 ) ,
        CN2VN_sign  => CN_sign_temp( 4735 downto 4704),
        CN2VN_bit   => CN_data_temp( 4735 downto 4704)
    );
    CN148 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4767 downto 4736 ) ,
        VN2CN_bit   => CN_data_in( 4767 downto 4736 ) ,
        CN2VN_sign  => CN_sign_temp( 4767 downto 4736),
        CN2VN_bit   => CN_data_temp( 4767 downto 4736)
    );
    CN149 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4799 downto 4768 ) ,
        VN2CN_bit   => CN_data_in( 4799 downto 4768 ) ,
        CN2VN_sign  => CN_sign_temp( 4799 downto 4768),
        CN2VN_bit   => CN_data_temp( 4799 downto 4768)
    );
    CN150 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4831 downto 4800 ) ,
        VN2CN_bit   => CN_data_in( 4831 downto 4800 ) ,
        CN2VN_sign  => CN_sign_temp( 4831 downto 4800),
        CN2VN_bit   => CN_data_temp( 4831 downto 4800)
    );
    CN151 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4863 downto 4832 ) ,
        VN2CN_bit   => CN_data_in( 4863 downto 4832 ) ,
        CN2VN_sign  => CN_sign_temp( 4863 downto 4832),
        CN2VN_bit   => CN_data_temp( 4863 downto 4832)
    );
    CN152 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4895 downto 4864 ) ,
        VN2CN_bit   => CN_data_in( 4895 downto 4864 ) ,
        CN2VN_sign  => CN_sign_temp( 4895 downto 4864),
        CN2VN_bit   => CN_data_temp( 4895 downto 4864)
    );
    CN153 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4927 downto 4896 ) ,
        VN2CN_bit   => CN_data_in( 4927 downto 4896 ) ,
        CN2VN_sign  => CN_sign_temp( 4927 downto 4896),
        CN2VN_bit   => CN_data_temp( 4927 downto 4896)
    );
    CN154 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4959 downto 4928 ) ,
        VN2CN_bit   => CN_data_in( 4959 downto 4928 ) ,
        CN2VN_sign  => CN_sign_temp( 4959 downto 4928),
        CN2VN_bit   => CN_data_temp( 4959 downto 4928)
    );
    CN155 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 4991 downto 4960 ) ,
        VN2CN_bit   => CN_data_in( 4991 downto 4960 ) ,
        CN2VN_sign  => CN_sign_temp( 4991 downto 4960),
        CN2VN_bit   => CN_data_temp( 4991 downto 4960)
    );
    CN156 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5023 downto 4992 ) ,
        VN2CN_bit   => CN_data_in( 5023 downto 4992 ) ,
        CN2VN_sign  => CN_sign_temp( 5023 downto 4992),
        CN2VN_bit   => CN_data_temp( 5023 downto 4992)
    );
    CN157 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5055 downto 5024 ) ,
        VN2CN_bit   => CN_data_in( 5055 downto 5024 ) ,
        CN2VN_sign  => CN_sign_temp( 5055 downto 5024),
        CN2VN_bit   => CN_data_temp( 5055 downto 5024)
    );
    CN158 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5087 downto 5056 ) ,
        VN2CN_bit   => CN_data_in( 5087 downto 5056 ) ,
        CN2VN_sign  => CN_sign_temp( 5087 downto 5056),
        CN2VN_bit   => CN_data_temp( 5087 downto 5056)
    );
    CN159 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5119 downto 5088 ) ,
        VN2CN_bit   => CN_data_in( 5119 downto 5088 ) ,
        CN2VN_sign  => CN_sign_temp( 5119 downto 5088),
        CN2VN_bit   => CN_data_temp( 5119 downto 5088)
    );
    CN160 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5151 downto 5120 ) ,
        VN2CN_bit   => CN_data_in( 5151 downto 5120 ) ,
        CN2VN_sign  => CN_sign_temp( 5151 downto 5120),
        CN2VN_bit   => CN_data_temp( 5151 downto 5120)
    );
    CN161 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5183 downto 5152 ) ,
        VN2CN_bit   => CN_data_in( 5183 downto 5152 ) ,
        CN2VN_sign  => CN_sign_temp( 5183 downto 5152),
        CN2VN_bit   => CN_data_temp( 5183 downto 5152)
    );
    CN162 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5215 downto 5184 ) ,
        VN2CN_bit   => CN_data_in( 5215 downto 5184 ) ,
        CN2VN_sign  => CN_sign_temp( 5215 downto 5184),
        CN2VN_bit   => CN_data_temp( 5215 downto 5184)
    );
    CN163 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5247 downto 5216 ) ,
        VN2CN_bit   => CN_data_in( 5247 downto 5216 ) ,
        CN2VN_sign  => CN_sign_temp( 5247 downto 5216),
        CN2VN_bit   => CN_data_temp( 5247 downto 5216)
    );
    CN164 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5279 downto 5248 ) ,
        VN2CN_bit   => CN_data_in( 5279 downto 5248 ) ,
        CN2VN_sign  => CN_sign_temp( 5279 downto 5248),
        CN2VN_bit   => CN_data_temp( 5279 downto 5248)
    );
    CN165 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5311 downto 5280 ) ,
        VN2CN_bit   => CN_data_in( 5311 downto 5280 ) ,
        CN2VN_sign  => CN_sign_temp( 5311 downto 5280),
        CN2VN_bit   => CN_data_temp( 5311 downto 5280)
    );
    CN166 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5343 downto 5312 ) ,
        VN2CN_bit   => CN_data_in( 5343 downto 5312 ) ,
        CN2VN_sign  => CN_sign_temp( 5343 downto 5312),
        CN2VN_bit   => CN_data_temp( 5343 downto 5312)
    );
    CN167 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5375 downto 5344 ) ,
        VN2CN_bit   => CN_data_in( 5375 downto 5344 ) ,
        CN2VN_sign  => CN_sign_temp( 5375 downto 5344),
        CN2VN_bit   => CN_data_temp( 5375 downto 5344)
    );
    CN168 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5407 downto 5376 ) ,
        VN2CN_bit   => CN_data_in( 5407 downto 5376 ) ,
        CN2VN_sign  => CN_sign_temp( 5407 downto 5376),
        CN2VN_bit   => CN_data_temp( 5407 downto 5376)
    );
    CN169 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5439 downto 5408 ) ,
        VN2CN_bit   => CN_data_in( 5439 downto 5408 ) ,
        CN2VN_sign  => CN_sign_temp( 5439 downto 5408),
        CN2VN_bit   => CN_data_temp( 5439 downto 5408)
    );
    CN170 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5471 downto 5440 ) ,
        VN2CN_bit   => CN_data_in( 5471 downto 5440 ) ,
        CN2VN_sign  => CN_sign_temp( 5471 downto 5440),
        CN2VN_bit   => CN_data_temp( 5471 downto 5440)
    );
    CN171 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5503 downto 5472 ) ,
        VN2CN_bit   => CN_data_in( 5503 downto 5472 ) ,
        CN2VN_sign  => CN_sign_temp( 5503 downto 5472),
        CN2VN_bit   => CN_data_temp( 5503 downto 5472)
    );
    CN172 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5535 downto 5504 ) ,
        VN2CN_bit   => CN_data_in( 5535 downto 5504 ) ,
        CN2VN_sign  => CN_sign_temp( 5535 downto 5504),
        CN2VN_bit   => CN_data_temp( 5535 downto 5504)
    );
    CN173 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5567 downto 5536 ) ,
        VN2CN_bit   => CN_data_in( 5567 downto 5536 ) ,
        CN2VN_sign  => CN_sign_temp( 5567 downto 5536),
        CN2VN_bit   => CN_data_temp( 5567 downto 5536)
    );
    CN174 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5599 downto 5568 ) ,
        VN2CN_bit   => CN_data_in( 5599 downto 5568 ) ,
        CN2VN_sign  => CN_sign_temp( 5599 downto 5568),
        CN2VN_bit   => CN_data_temp( 5599 downto 5568)
    );
    CN175 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5631 downto 5600 ) ,
        VN2CN_bit   => CN_data_in( 5631 downto 5600 ) ,
        CN2VN_sign  => CN_sign_temp( 5631 downto 5600),
        CN2VN_bit   => CN_data_temp( 5631 downto 5600)
    );
    CN176 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5663 downto 5632 ) ,
        VN2CN_bit   => CN_data_in( 5663 downto 5632 ) ,
        CN2VN_sign  => CN_sign_temp( 5663 downto 5632),
        CN2VN_bit   => CN_data_temp( 5663 downto 5632)
    );
    CN177 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5695 downto 5664 ) ,
        VN2CN_bit   => CN_data_in( 5695 downto 5664 ) ,
        CN2VN_sign  => CN_sign_temp( 5695 downto 5664),
        CN2VN_bit   => CN_data_temp( 5695 downto 5664)
    );
    CN178 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5727 downto 5696 ) ,
        VN2CN_bit   => CN_data_in( 5727 downto 5696 ) ,
        CN2VN_sign  => CN_sign_temp( 5727 downto 5696),
        CN2VN_bit   => CN_data_temp( 5727 downto 5696)
    );
    CN179 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5759 downto 5728 ) ,
        VN2CN_bit   => CN_data_in( 5759 downto 5728 ) ,
        CN2VN_sign  => CN_sign_temp( 5759 downto 5728),
        CN2VN_bit   => CN_data_temp( 5759 downto 5728)
    );
    CN180 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5791 downto 5760 ) ,
        VN2CN_bit   => CN_data_in( 5791 downto 5760 ) ,
        CN2VN_sign  => CN_sign_temp( 5791 downto 5760),
        CN2VN_bit   => CN_data_temp( 5791 downto 5760)
    );
    CN181 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5823 downto 5792 ) ,
        VN2CN_bit   => CN_data_in( 5823 downto 5792 ) ,
        CN2VN_sign  => CN_sign_temp( 5823 downto 5792),
        CN2VN_bit   => CN_data_temp( 5823 downto 5792)
    );
    CN182 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5855 downto 5824 ) ,
        VN2CN_bit   => CN_data_in( 5855 downto 5824 ) ,
        CN2VN_sign  => CN_sign_temp( 5855 downto 5824),
        CN2VN_bit   => CN_data_temp( 5855 downto 5824)
    );
    CN183 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5887 downto 5856 ) ,
        VN2CN_bit   => CN_data_in( 5887 downto 5856 ) ,
        CN2VN_sign  => CN_sign_temp( 5887 downto 5856),
        CN2VN_bit   => CN_data_temp( 5887 downto 5856)
    );
    CN184 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5919 downto 5888 ) ,
        VN2CN_bit   => CN_data_in( 5919 downto 5888 ) ,
        CN2VN_sign  => CN_sign_temp( 5919 downto 5888),
        CN2VN_bit   => CN_data_temp( 5919 downto 5888)
    );
    CN185 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5951 downto 5920 ) ,
        VN2CN_bit   => CN_data_in( 5951 downto 5920 ) ,
        CN2VN_sign  => CN_sign_temp( 5951 downto 5920),
        CN2VN_bit   => CN_data_temp( 5951 downto 5920)
    );
    CN186 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 5983 downto 5952 ) ,
        VN2CN_bit   => CN_data_in( 5983 downto 5952 ) ,
        CN2VN_sign  => CN_sign_temp( 5983 downto 5952),
        CN2VN_bit   => CN_data_temp( 5983 downto 5952)
    );
    CN187 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6015 downto 5984 ) ,
        VN2CN_bit   => CN_data_in( 6015 downto 5984 ) ,
        CN2VN_sign  => CN_sign_temp( 6015 downto 5984),
        CN2VN_bit   => CN_data_temp( 6015 downto 5984)
    );
    CN188 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6047 downto 6016 ) ,
        VN2CN_bit   => CN_data_in( 6047 downto 6016 ) ,
        CN2VN_sign  => CN_sign_temp( 6047 downto 6016),
        CN2VN_bit   => CN_data_temp( 6047 downto 6016)
    );
    CN189 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6079 downto 6048 ) ,
        VN2CN_bit   => CN_data_in( 6079 downto 6048 ) ,
        CN2VN_sign  => CN_sign_temp( 6079 downto 6048),
        CN2VN_bit   => CN_data_temp( 6079 downto 6048)
    );
    CN190 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6111 downto 6080 ) ,
        VN2CN_bit   => CN_data_in( 6111 downto 6080 ) ,
        CN2VN_sign  => CN_sign_temp( 6111 downto 6080),
        CN2VN_bit   => CN_data_temp( 6111 downto 6080)
    );
    CN191 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6143 downto 6112 ) ,
        VN2CN_bit   => CN_data_in( 6143 downto 6112 ) ,
        CN2VN_sign  => CN_sign_temp( 6143 downto 6112),
        CN2VN_bit   => CN_data_temp( 6143 downto 6112)
    );
    CN192 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6175 downto 6144 ) ,
        VN2CN_bit   => CN_data_in( 6175 downto 6144 ) ,
        CN2VN_sign  => CN_sign_temp( 6175 downto 6144),
        CN2VN_bit   => CN_data_temp( 6175 downto 6144)
    );
    CN193 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6207 downto 6176 ) ,
        VN2CN_bit   => CN_data_in( 6207 downto 6176 ) ,
        CN2VN_sign  => CN_sign_temp( 6207 downto 6176),
        CN2VN_bit   => CN_data_temp( 6207 downto 6176)
    );
    CN194 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6239 downto 6208 ) ,
        VN2CN_bit   => CN_data_in( 6239 downto 6208 ) ,
        CN2VN_sign  => CN_sign_temp( 6239 downto 6208),
        CN2VN_bit   => CN_data_temp( 6239 downto 6208)
    );
    CN195 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6271 downto 6240 ) ,
        VN2CN_bit   => CN_data_in( 6271 downto 6240 ) ,
        CN2VN_sign  => CN_sign_temp( 6271 downto 6240),
        CN2VN_bit   => CN_data_temp( 6271 downto 6240)
    );
    CN196 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6303 downto 6272 ) ,
        VN2CN_bit   => CN_data_in( 6303 downto 6272 ) ,
        CN2VN_sign  => CN_sign_temp( 6303 downto 6272),
        CN2VN_bit   => CN_data_temp( 6303 downto 6272)
    );
    CN197 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6335 downto 6304 ) ,
        VN2CN_bit   => CN_data_in( 6335 downto 6304 ) ,
        CN2VN_sign  => CN_sign_temp( 6335 downto 6304),
        CN2VN_bit   => CN_data_temp( 6335 downto 6304)
    );
    CN198 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6367 downto 6336 ) ,
        VN2CN_bit   => CN_data_in( 6367 downto 6336 ) ,
        CN2VN_sign  => CN_sign_temp( 6367 downto 6336),
        CN2VN_bit   => CN_data_temp( 6367 downto 6336)
    );
    CN199 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6399 downto 6368 ) ,
        VN2CN_bit   => CN_data_in( 6399 downto 6368 ) ,
        CN2VN_sign  => CN_sign_temp( 6399 downto 6368),
        CN2VN_bit   => CN_data_temp( 6399 downto 6368)
    );
    CN200 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6431 downto 6400 ) ,
        VN2CN_bit   => CN_data_in( 6431 downto 6400 ) ,
        CN2VN_sign  => CN_sign_temp( 6431 downto 6400),
        CN2VN_bit   => CN_data_temp( 6431 downto 6400)
    );
    CN201 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6463 downto 6432 ) ,
        VN2CN_bit   => CN_data_in( 6463 downto 6432 ) ,
        CN2VN_sign  => CN_sign_temp( 6463 downto 6432),
        CN2VN_bit   => CN_data_temp( 6463 downto 6432)
    );
    CN202 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6495 downto 6464 ) ,
        VN2CN_bit   => CN_data_in( 6495 downto 6464 ) ,
        CN2VN_sign  => CN_sign_temp( 6495 downto 6464),
        CN2VN_bit   => CN_data_temp( 6495 downto 6464)
    );
    CN203 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6527 downto 6496 ) ,
        VN2CN_bit   => CN_data_in( 6527 downto 6496 ) ,
        CN2VN_sign  => CN_sign_temp( 6527 downto 6496),
        CN2VN_bit   => CN_data_temp( 6527 downto 6496)
    );
    CN204 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6559 downto 6528 ) ,
        VN2CN_bit   => CN_data_in( 6559 downto 6528 ) ,
        CN2VN_sign  => CN_sign_temp( 6559 downto 6528),
        CN2VN_bit   => CN_data_temp( 6559 downto 6528)
    );
    CN205 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6591 downto 6560 ) ,
        VN2CN_bit   => CN_data_in( 6591 downto 6560 ) ,
        CN2VN_sign  => CN_sign_temp( 6591 downto 6560),
        CN2VN_bit   => CN_data_temp( 6591 downto 6560)
    );
    CN206 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6623 downto 6592 ) ,
        VN2CN_bit   => CN_data_in( 6623 downto 6592 ) ,
        CN2VN_sign  => CN_sign_temp( 6623 downto 6592),
        CN2VN_bit   => CN_data_temp( 6623 downto 6592)
    );
    CN207 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6655 downto 6624 ) ,
        VN2CN_bit   => CN_data_in( 6655 downto 6624 ) ,
        CN2VN_sign  => CN_sign_temp( 6655 downto 6624),
        CN2VN_bit   => CN_data_temp( 6655 downto 6624)
    );
    CN208 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6687 downto 6656 ) ,
        VN2CN_bit   => CN_data_in( 6687 downto 6656 ) ,
        CN2VN_sign  => CN_sign_temp( 6687 downto 6656),
        CN2VN_bit   => CN_data_temp( 6687 downto 6656)
    );
    CN209 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6719 downto 6688 ) ,
        VN2CN_bit   => CN_data_in( 6719 downto 6688 ) ,
        CN2VN_sign  => CN_sign_temp( 6719 downto 6688),
        CN2VN_bit   => CN_data_temp( 6719 downto 6688)
    );
    CN210 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6751 downto 6720 ) ,
        VN2CN_bit   => CN_data_in( 6751 downto 6720 ) ,
        CN2VN_sign  => CN_sign_temp( 6751 downto 6720),
        CN2VN_bit   => CN_data_temp( 6751 downto 6720)
    );
    CN211 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6783 downto 6752 ) ,
        VN2CN_bit   => CN_data_in( 6783 downto 6752 ) ,
        CN2VN_sign  => CN_sign_temp( 6783 downto 6752),
        CN2VN_bit   => CN_data_temp( 6783 downto 6752)
    );
    CN212 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6815 downto 6784 ) ,
        VN2CN_bit   => CN_data_in( 6815 downto 6784 ) ,
        CN2VN_sign  => CN_sign_temp( 6815 downto 6784),
        CN2VN_bit   => CN_data_temp( 6815 downto 6784)
    );
    CN213 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6847 downto 6816 ) ,
        VN2CN_bit   => CN_data_in( 6847 downto 6816 ) ,
        CN2VN_sign  => CN_sign_temp( 6847 downto 6816),
        CN2VN_bit   => CN_data_temp( 6847 downto 6816)
    );
    CN214 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6879 downto 6848 ) ,
        VN2CN_bit   => CN_data_in( 6879 downto 6848 ) ,
        CN2VN_sign  => CN_sign_temp( 6879 downto 6848),
        CN2VN_bit   => CN_data_temp( 6879 downto 6848)
    );
    CN215 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6911 downto 6880 ) ,
        VN2CN_bit   => CN_data_in( 6911 downto 6880 ) ,
        CN2VN_sign  => CN_sign_temp( 6911 downto 6880),
        CN2VN_bit   => CN_data_temp( 6911 downto 6880)
    );
    CN216 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6943 downto 6912 ) ,
        VN2CN_bit   => CN_data_in( 6943 downto 6912 ) ,
        CN2VN_sign  => CN_sign_temp( 6943 downto 6912),
        CN2VN_bit   => CN_data_temp( 6943 downto 6912)
    );
    CN217 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 6975 downto 6944 ) ,
        VN2CN_bit   => CN_data_in( 6975 downto 6944 ) ,
        CN2VN_sign  => CN_sign_temp( 6975 downto 6944),
        CN2VN_bit   => CN_data_temp( 6975 downto 6944)
    );
    CN218 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7007 downto 6976 ) ,
        VN2CN_bit   => CN_data_in( 7007 downto 6976 ) ,
        CN2VN_sign  => CN_sign_temp( 7007 downto 6976),
        CN2VN_bit   => CN_data_temp( 7007 downto 6976)
    );
    CN219 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7039 downto 7008 ) ,
        VN2CN_bit   => CN_data_in( 7039 downto 7008 ) ,
        CN2VN_sign  => CN_sign_temp( 7039 downto 7008),
        CN2VN_bit   => CN_data_temp( 7039 downto 7008)
    );
    CN220 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7071 downto 7040 ) ,
        VN2CN_bit   => CN_data_in( 7071 downto 7040 ) ,
        CN2VN_sign  => CN_sign_temp( 7071 downto 7040),
        CN2VN_bit   => CN_data_temp( 7071 downto 7040)
    );
    CN221 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7103 downto 7072 ) ,
        VN2CN_bit   => CN_data_in( 7103 downto 7072 ) ,
        CN2VN_sign  => CN_sign_temp( 7103 downto 7072),
        CN2VN_bit   => CN_data_temp( 7103 downto 7072)
    );
    CN222 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7135 downto 7104 ) ,
        VN2CN_bit   => CN_data_in( 7135 downto 7104 ) ,
        CN2VN_sign  => CN_sign_temp( 7135 downto 7104),
        CN2VN_bit   => CN_data_temp( 7135 downto 7104)
    );
    CN223 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7167 downto 7136 ) ,
        VN2CN_bit   => CN_data_in( 7167 downto 7136 ) ,
        CN2VN_sign  => CN_sign_temp( 7167 downto 7136),
        CN2VN_bit   => CN_data_temp( 7167 downto 7136)
    );
    CN224 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7199 downto 7168 ) ,
        VN2CN_bit   => CN_data_in( 7199 downto 7168 ) ,
        CN2VN_sign  => CN_sign_temp( 7199 downto 7168),
        CN2VN_bit   => CN_data_temp( 7199 downto 7168)
    );
    CN225 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7231 downto 7200 ) ,
        VN2CN_bit   => CN_data_in( 7231 downto 7200 ) ,
        CN2VN_sign  => CN_sign_temp( 7231 downto 7200),
        CN2VN_bit   => CN_data_temp( 7231 downto 7200)
    );
    CN226 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7263 downto 7232 ) ,
        VN2CN_bit   => CN_data_in( 7263 downto 7232 ) ,
        CN2VN_sign  => CN_sign_temp( 7263 downto 7232),
        CN2VN_bit   => CN_data_temp( 7263 downto 7232)
    );
    CN227 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7295 downto 7264 ) ,
        VN2CN_bit   => CN_data_in( 7295 downto 7264 ) ,
        CN2VN_sign  => CN_sign_temp( 7295 downto 7264),
        CN2VN_bit   => CN_data_temp( 7295 downto 7264)
    );
    CN228 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7327 downto 7296 ) ,
        VN2CN_bit   => CN_data_in( 7327 downto 7296 ) ,
        CN2VN_sign  => CN_sign_temp( 7327 downto 7296),
        CN2VN_bit   => CN_data_temp( 7327 downto 7296)
    );
    CN229 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7359 downto 7328 ) ,
        VN2CN_bit   => CN_data_in( 7359 downto 7328 ) ,
        CN2VN_sign  => CN_sign_temp( 7359 downto 7328),
        CN2VN_bit   => CN_data_temp( 7359 downto 7328)
    );
    CN230 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7391 downto 7360 ) ,
        VN2CN_bit   => CN_data_in( 7391 downto 7360 ) ,
        CN2VN_sign  => CN_sign_temp( 7391 downto 7360),
        CN2VN_bit   => CN_data_temp( 7391 downto 7360)
    );
    CN231 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7423 downto 7392 ) ,
        VN2CN_bit   => CN_data_in( 7423 downto 7392 ) ,
        CN2VN_sign  => CN_sign_temp( 7423 downto 7392),
        CN2VN_bit   => CN_data_temp( 7423 downto 7392)
    );
    CN232 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7455 downto 7424 ) ,
        VN2CN_bit   => CN_data_in( 7455 downto 7424 ) ,
        CN2VN_sign  => CN_sign_temp( 7455 downto 7424),
        CN2VN_bit   => CN_data_temp( 7455 downto 7424)
    );
    CN233 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7487 downto 7456 ) ,
        VN2CN_bit   => CN_data_in( 7487 downto 7456 ) ,
        CN2VN_sign  => CN_sign_temp( 7487 downto 7456),
        CN2VN_bit   => CN_data_temp( 7487 downto 7456)
    );
    CN234 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7519 downto 7488 ) ,
        VN2CN_bit   => CN_data_in( 7519 downto 7488 ) ,
        CN2VN_sign  => CN_sign_temp( 7519 downto 7488),
        CN2VN_bit   => CN_data_temp( 7519 downto 7488)
    );
    CN235 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7551 downto 7520 ) ,
        VN2CN_bit   => CN_data_in( 7551 downto 7520 ) ,
        CN2VN_sign  => CN_sign_temp( 7551 downto 7520),
        CN2VN_bit   => CN_data_temp( 7551 downto 7520)
    );
    CN236 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7583 downto 7552 ) ,
        VN2CN_bit   => CN_data_in( 7583 downto 7552 ) ,
        CN2VN_sign  => CN_sign_temp( 7583 downto 7552),
        CN2VN_bit   => CN_data_temp( 7583 downto 7552)
    );
    CN237 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7615 downto 7584 ) ,
        VN2CN_bit   => CN_data_in( 7615 downto 7584 ) ,
        CN2VN_sign  => CN_sign_temp( 7615 downto 7584),
        CN2VN_bit   => CN_data_temp( 7615 downto 7584)
    );
    CN238 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7647 downto 7616 ) ,
        VN2CN_bit   => CN_data_in( 7647 downto 7616 ) ,
        CN2VN_sign  => CN_sign_temp( 7647 downto 7616),
        CN2VN_bit   => CN_data_temp( 7647 downto 7616)
    );
    CN239 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7679 downto 7648 ) ,
        VN2CN_bit   => CN_data_in( 7679 downto 7648 ) ,
        CN2VN_sign  => CN_sign_temp( 7679 downto 7648),
        CN2VN_bit   => CN_data_temp( 7679 downto 7648)
    );
    CN240 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7711 downto 7680 ) ,
        VN2CN_bit   => CN_data_in( 7711 downto 7680 ) ,
        CN2VN_sign  => CN_sign_temp( 7711 downto 7680),
        CN2VN_bit   => CN_data_temp( 7711 downto 7680)
    );
    CN241 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7743 downto 7712 ) ,
        VN2CN_bit   => CN_data_in( 7743 downto 7712 ) ,
        CN2VN_sign  => CN_sign_temp( 7743 downto 7712),
        CN2VN_bit   => CN_data_temp( 7743 downto 7712)
    );
    CN242 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7775 downto 7744 ) ,
        VN2CN_bit   => CN_data_in( 7775 downto 7744 ) ,
        CN2VN_sign  => CN_sign_temp( 7775 downto 7744),
        CN2VN_bit   => CN_data_temp( 7775 downto 7744)
    );
    CN243 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7807 downto 7776 ) ,
        VN2CN_bit   => CN_data_in( 7807 downto 7776 ) ,
        CN2VN_sign  => CN_sign_temp( 7807 downto 7776),
        CN2VN_bit   => CN_data_temp( 7807 downto 7776)
    );
    CN244 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7839 downto 7808 ) ,
        VN2CN_bit   => CN_data_in( 7839 downto 7808 ) ,
        CN2VN_sign  => CN_sign_temp( 7839 downto 7808),
        CN2VN_bit   => CN_data_temp( 7839 downto 7808)
    );
    CN245 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7871 downto 7840 ) ,
        VN2CN_bit   => CN_data_in( 7871 downto 7840 ) ,
        CN2VN_sign  => CN_sign_temp( 7871 downto 7840),
        CN2VN_bit   => CN_data_temp( 7871 downto 7840)
    );
    CN246 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7903 downto 7872 ) ,
        VN2CN_bit   => CN_data_in( 7903 downto 7872 ) ,
        CN2VN_sign  => CN_sign_temp( 7903 downto 7872),
        CN2VN_bit   => CN_data_temp( 7903 downto 7872)
    );
    CN247 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7935 downto 7904 ) ,
        VN2CN_bit   => CN_data_in( 7935 downto 7904 ) ,
        CN2VN_sign  => CN_sign_temp( 7935 downto 7904),
        CN2VN_bit   => CN_data_temp( 7935 downto 7904)
    );
    CN248 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7967 downto 7936 ) ,
        VN2CN_bit   => CN_data_in( 7967 downto 7936 ) ,
        CN2VN_sign  => CN_sign_temp( 7967 downto 7936),
        CN2VN_bit   => CN_data_temp( 7967 downto 7936)
    );
    CN249 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 7999 downto 7968 ) ,
        VN2CN_bit   => CN_data_in( 7999 downto 7968 ) ,
        CN2VN_sign  => CN_sign_temp( 7999 downto 7968),
        CN2VN_bit   => CN_data_temp( 7999 downto 7968)
    );
    CN250 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8031 downto 8000 ) ,
        VN2CN_bit   => CN_data_in( 8031 downto 8000 ) ,
        CN2VN_sign  => CN_sign_temp( 8031 downto 8000),
        CN2VN_bit   => CN_data_temp( 8031 downto 8000)
    );
    CN251 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8063 downto 8032 ) ,
        VN2CN_bit   => CN_data_in( 8063 downto 8032 ) ,
        CN2VN_sign  => CN_sign_temp( 8063 downto 8032),
        CN2VN_bit   => CN_data_temp( 8063 downto 8032)
    );
    CN252 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8095 downto 8064 ) ,
        VN2CN_bit   => CN_data_in( 8095 downto 8064 ) ,
        CN2VN_sign  => CN_sign_temp( 8095 downto 8064),
        CN2VN_bit   => CN_data_temp( 8095 downto 8064)
    );
    CN253 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8127 downto 8096 ) ,
        VN2CN_bit   => CN_data_in( 8127 downto 8096 ) ,
        CN2VN_sign  => CN_sign_temp( 8127 downto 8096),
        CN2VN_bit   => CN_data_temp( 8127 downto 8096)
    );
    CN254 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8159 downto 8128 ) ,
        VN2CN_bit   => CN_data_in( 8159 downto 8128 ) ,
        CN2VN_sign  => CN_sign_temp( 8159 downto 8128),
        CN2VN_bit   => CN_data_temp( 8159 downto 8128)
    );
    CN255 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8191 downto 8160 ) ,
        VN2CN_bit   => CN_data_in( 8191 downto 8160 ) ,
        CN2VN_sign  => CN_sign_temp( 8191 downto 8160),
        CN2VN_bit   => CN_data_temp( 8191 downto 8160)
    );
    CN256 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8223 downto 8192 ) ,
        VN2CN_bit   => CN_data_in( 8223 downto 8192 ) ,
        CN2VN_sign  => CN_sign_temp( 8223 downto 8192),
        CN2VN_bit   => CN_data_temp( 8223 downto 8192)
    );
    CN257 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8255 downto 8224 ) ,
        VN2CN_bit   => CN_data_in( 8255 downto 8224 ) ,
        CN2VN_sign  => CN_sign_temp( 8255 downto 8224),
        CN2VN_bit   => CN_data_temp( 8255 downto 8224)
    );
    CN258 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8287 downto 8256 ) ,
        VN2CN_bit   => CN_data_in( 8287 downto 8256 ) ,
        CN2VN_sign  => CN_sign_temp( 8287 downto 8256),
        CN2VN_bit   => CN_data_temp( 8287 downto 8256)
    );
    CN259 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8319 downto 8288 ) ,
        VN2CN_bit   => CN_data_in( 8319 downto 8288 ) ,
        CN2VN_sign  => CN_sign_temp( 8319 downto 8288),
        CN2VN_bit   => CN_data_temp( 8319 downto 8288)
    );
    CN260 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8351 downto 8320 ) ,
        VN2CN_bit   => CN_data_in( 8351 downto 8320 ) ,
        CN2VN_sign  => CN_sign_temp( 8351 downto 8320),
        CN2VN_bit   => CN_data_temp( 8351 downto 8320)
    );
    CN261 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8383 downto 8352 ) ,
        VN2CN_bit   => CN_data_in( 8383 downto 8352 ) ,
        CN2VN_sign  => CN_sign_temp( 8383 downto 8352),
        CN2VN_bit   => CN_data_temp( 8383 downto 8352)
    );
    CN262 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8415 downto 8384 ) ,
        VN2CN_bit   => CN_data_in( 8415 downto 8384 ) ,
        CN2VN_sign  => CN_sign_temp( 8415 downto 8384),
        CN2VN_bit   => CN_data_temp( 8415 downto 8384)
    );
    CN263 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8447 downto 8416 ) ,
        VN2CN_bit   => CN_data_in( 8447 downto 8416 ) ,
        CN2VN_sign  => CN_sign_temp( 8447 downto 8416),
        CN2VN_bit   => CN_data_temp( 8447 downto 8416)
    );
    CN264 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8479 downto 8448 ) ,
        VN2CN_bit   => CN_data_in( 8479 downto 8448 ) ,
        CN2VN_sign  => CN_sign_temp( 8479 downto 8448),
        CN2VN_bit   => CN_data_temp( 8479 downto 8448)
    );
    CN265 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8511 downto 8480 ) ,
        VN2CN_bit   => CN_data_in( 8511 downto 8480 ) ,
        CN2VN_sign  => CN_sign_temp( 8511 downto 8480),
        CN2VN_bit   => CN_data_temp( 8511 downto 8480)
    );
    CN266 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8543 downto 8512 ) ,
        VN2CN_bit   => CN_data_in( 8543 downto 8512 ) ,
        CN2VN_sign  => CN_sign_temp( 8543 downto 8512),
        CN2VN_bit   => CN_data_temp( 8543 downto 8512)
    );
    CN267 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8575 downto 8544 ) ,
        VN2CN_bit   => CN_data_in( 8575 downto 8544 ) ,
        CN2VN_sign  => CN_sign_temp( 8575 downto 8544),
        CN2VN_bit   => CN_data_temp( 8575 downto 8544)
    );
    CN268 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8607 downto 8576 ) ,
        VN2CN_bit   => CN_data_in( 8607 downto 8576 ) ,
        CN2VN_sign  => CN_sign_temp( 8607 downto 8576),
        CN2VN_bit   => CN_data_temp( 8607 downto 8576)
    );
    CN269 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8639 downto 8608 ) ,
        VN2CN_bit   => CN_data_in( 8639 downto 8608 ) ,
        CN2VN_sign  => CN_sign_temp( 8639 downto 8608),
        CN2VN_bit   => CN_data_temp( 8639 downto 8608)
    );
    CN270 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8671 downto 8640 ) ,
        VN2CN_bit   => CN_data_in( 8671 downto 8640 ) ,
        CN2VN_sign  => CN_sign_temp( 8671 downto 8640),
        CN2VN_bit   => CN_data_temp( 8671 downto 8640)
    );
    CN271 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8703 downto 8672 ) ,
        VN2CN_bit   => CN_data_in( 8703 downto 8672 ) ,
        CN2VN_sign  => CN_sign_temp( 8703 downto 8672),
        CN2VN_bit   => CN_data_temp( 8703 downto 8672)
    );
    CN272 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8735 downto 8704 ) ,
        VN2CN_bit   => CN_data_in( 8735 downto 8704 ) ,
        CN2VN_sign  => CN_sign_temp( 8735 downto 8704),
        CN2VN_bit   => CN_data_temp( 8735 downto 8704)
    );
    CN273 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8767 downto 8736 ) ,
        VN2CN_bit   => CN_data_in( 8767 downto 8736 ) ,
        CN2VN_sign  => CN_sign_temp( 8767 downto 8736),
        CN2VN_bit   => CN_data_temp( 8767 downto 8736)
    );
    CN274 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8799 downto 8768 ) ,
        VN2CN_bit   => CN_data_in( 8799 downto 8768 ) ,
        CN2VN_sign  => CN_sign_temp( 8799 downto 8768),
        CN2VN_bit   => CN_data_temp( 8799 downto 8768)
    );
    CN275 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8831 downto 8800 ) ,
        VN2CN_bit   => CN_data_in( 8831 downto 8800 ) ,
        CN2VN_sign  => CN_sign_temp( 8831 downto 8800),
        CN2VN_bit   => CN_data_temp( 8831 downto 8800)
    );
    CN276 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8863 downto 8832 ) ,
        VN2CN_bit   => CN_data_in( 8863 downto 8832 ) ,
        CN2VN_sign  => CN_sign_temp( 8863 downto 8832),
        CN2VN_bit   => CN_data_temp( 8863 downto 8832)
    );
    CN277 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8895 downto 8864 ) ,
        VN2CN_bit   => CN_data_in( 8895 downto 8864 ) ,
        CN2VN_sign  => CN_sign_temp( 8895 downto 8864),
        CN2VN_bit   => CN_data_temp( 8895 downto 8864)
    );
    CN278 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8927 downto 8896 ) ,
        VN2CN_bit   => CN_data_in( 8927 downto 8896 ) ,
        CN2VN_sign  => CN_sign_temp( 8927 downto 8896),
        CN2VN_bit   => CN_data_temp( 8927 downto 8896)
    );
    CN279 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8959 downto 8928 ) ,
        VN2CN_bit   => CN_data_in( 8959 downto 8928 ) ,
        CN2VN_sign  => CN_sign_temp( 8959 downto 8928),
        CN2VN_bit   => CN_data_temp( 8959 downto 8928)
    );
    CN280 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 8991 downto 8960 ) ,
        VN2CN_bit   => CN_data_in( 8991 downto 8960 ) ,
        CN2VN_sign  => CN_sign_temp( 8991 downto 8960),
        CN2VN_bit   => CN_data_temp( 8991 downto 8960)
    );
    CN281 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9023 downto 8992 ) ,
        VN2CN_bit   => CN_data_in( 9023 downto 8992 ) ,
        CN2VN_sign  => CN_sign_temp( 9023 downto 8992),
        CN2VN_bit   => CN_data_temp( 9023 downto 8992)
    );
    CN282 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9055 downto 9024 ) ,
        VN2CN_bit   => CN_data_in( 9055 downto 9024 ) ,
        CN2VN_sign  => CN_sign_temp( 9055 downto 9024),
        CN2VN_bit   => CN_data_temp( 9055 downto 9024)
    );
    CN283 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9087 downto 9056 ) ,
        VN2CN_bit   => CN_data_in( 9087 downto 9056 ) ,
        CN2VN_sign  => CN_sign_temp( 9087 downto 9056),
        CN2VN_bit   => CN_data_temp( 9087 downto 9056)
    );
    CN284 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9119 downto 9088 ) ,
        VN2CN_bit   => CN_data_in( 9119 downto 9088 ) ,
        CN2VN_sign  => CN_sign_temp( 9119 downto 9088),
        CN2VN_bit   => CN_data_temp( 9119 downto 9088)
    );
    CN285 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9151 downto 9120 ) ,
        VN2CN_bit   => CN_data_in( 9151 downto 9120 ) ,
        CN2VN_sign  => CN_sign_temp( 9151 downto 9120),
        CN2VN_bit   => CN_data_temp( 9151 downto 9120)
    );
    CN286 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9183 downto 9152 ) ,
        VN2CN_bit   => CN_data_in( 9183 downto 9152 ) ,
        CN2VN_sign  => CN_sign_temp( 9183 downto 9152),
        CN2VN_bit   => CN_data_temp( 9183 downto 9152)
    );
    CN287 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9215 downto 9184 ) ,
        VN2CN_bit   => CN_data_in( 9215 downto 9184 ) ,
        CN2VN_sign  => CN_sign_temp( 9215 downto 9184),
        CN2VN_bit   => CN_data_temp( 9215 downto 9184)
    );
    CN288 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9247 downto 9216 ) ,
        VN2CN_bit   => CN_data_in( 9247 downto 9216 ) ,
        CN2VN_sign  => CN_sign_temp( 9247 downto 9216),
        CN2VN_bit   => CN_data_temp( 9247 downto 9216)
    );
    CN289 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9279 downto 9248 ) ,
        VN2CN_bit   => CN_data_in( 9279 downto 9248 ) ,
        CN2VN_sign  => CN_sign_temp( 9279 downto 9248),
        CN2VN_bit   => CN_data_temp( 9279 downto 9248)
    );
    CN290 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9311 downto 9280 ) ,
        VN2CN_bit   => CN_data_in( 9311 downto 9280 ) ,
        CN2VN_sign  => CN_sign_temp( 9311 downto 9280),
        CN2VN_bit   => CN_data_temp( 9311 downto 9280)
    );
    CN291 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9343 downto 9312 ) ,
        VN2CN_bit   => CN_data_in( 9343 downto 9312 ) ,
        CN2VN_sign  => CN_sign_temp( 9343 downto 9312),
        CN2VN_bit   => CN_data_temp( 9343 downto 9312)
    );
    CN292 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9375 downto 9344 ) ,
        VN2CN_bit   => CN_data_in( 9375 downto 9344 ) ,
        CN2VN_sign  => CN_sign_temp( 9375 downto 9344),
        CN2VN_bit   => CN_data_temp( 9375 downto 9344)
    );
    CN293 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9407 downto 9376 ) ,
        VN2CN_bit   => CN_data_in( 9407 downto 9376 ) ,
        CN2VN_sign  => CN_sign_temp( 9407 downto 9376),
        CN2VN_bit   => CN_data_temp( 9407 downto 9376)
    );
    CN294 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9439 downto 9408 ) ,
        VN2CN_bit   => CN_data_in( 9439 downto 9408 ) ,
        CN2VN_sign  => CN_sign_temp( 9439 downto 9408),
        CN2VN_bit   => CN_data_temp( 9439 downto 9408)
    );
    CN295 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9471 downto 9440 ) ,
        VN2CN_bit   => CN_data_in( 9471 downto 9440 ) ,
        CN2VN_sign  => CN_sign_temp( 9471 downto 9440),
        CN2VN_bit   => CN_data_temp( 9471 downto 9440)
    );
    CN296 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9503 downto 9472 ) ,
        VN2CN_bit   => CN_data_in( 9503 downto 9472 ) ,
        CN2VN_sign  => CN_sign_temp( 9503 downto 9472),
        CN2VN_bit   => CN_data_temp( 9503 downto 9472)
    );
    CN297 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9535 downto 9504 ) ,
        VN2CN_bit   => CN_data_in( 9535 downto 9504 ) ,
        CN2VN_sign  => CN_sign_temp( 9535 downto 9504),
        CN2VN_bit   => CN_data_temp( 9535 downto 9504)
    );
    CN298 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9567 downto 9536 ) ,
        VN2CN_bit   => CN_data_in( 9567 downto 9536 ) ,
        CN2VN_sign  => CN_sign_temp( 9567 downto 9536),
        CN2VN_bit   => CN_data_temp( 9567 downto 9536)
    );
    CN299 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9599 downto 9568 ) ,
        VN2CN_bit   => CN_data_in( 9599 downto 9568 ) ,
        CN2VN_sign  => CN_sign_temp( 9599 downto 9568),
        CN2VN_bit   => CN_data_temp( 9599 downto 9568)
    );
    CN300 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9631 downto 9600 ) ,
        VN2CN_bit   => CN_data_in( 9631 downto 9600 ) ,
        CN2VN_sign  => CN_sign_temp( 9631 downto 9600),
        CN2VN_bit   => CN_data_temp( 9631 downto 9600)
    );
    CN301 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9663 downto 9632 ) ,
        VN2CN_bit   => CN_data_in( 9663 downto 9632 ) ,
        CN2VN_sign  => CN_sign_temp( 9663 downto 9632),
        CN2VN_bit   => CN_data_temp( 9663 downto 9632)
    );
    CN302 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9695 downto 9664 ) ,
        VN2CN_bit   => CN_data_in( 9695 downto 9664 ) ,
        CN2VN_sign  => CN_sign_temp( 9695 downto 9664),
        CN2VN_bit   => CN_data_temp( 9695 downto 9664)
    );
    CN303 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9727 downto 9696 ) ,
        VN2CN_bit   => CN_data_in( 9727 downto 9696 ) ,
        CN2VN_sign  => CN_sign_temp( 9727 downto 9696),
        CN2VN_bit   => CN_data_temp( 9727 downto 9696)
    );
    CN304 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9759 downto 9728 ) ,
        VN2CN_bit   => CN_data_in( 9759 downto 9728 ) ,
        CN2VN_sign  => CN_sign_temp( 9759 downto 9728),
        CN2VN_bit   => CN_data_temp( 9759 downto 9728)
    );
    CN305 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9791 downto 9760 ) ,
        VN2CN_bit   => CN_data_in( 9791 downto 9760 ) ,
        CN2VN_sign  => CN_sign_temp( 9791 downto 9760),
        CN2VN_bit   => CN_data_temp( 9791 downto 9760)
    );
    CN306 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9823 downto 9792 ) ,
        VN2CN_bit   => CN_data_in( 9823 downto 9792 ) ,
        CN2VN_sign  => CN_sign_temp( 9823 downto 9792),
        CN2VN_bit   => CN_data_temp( 9823 downto 9792)
    );
    CN307 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9855 downto 9824 ) ,
        VN2CN_bit   => CN_data_in( 9855 downto 9824 ) ,
        CN2VN_sign  => CN_sign_temp( 9855 downto 9824),
        CN2VN_bit   => CN_data_temp( 9855 downto 9824)
    );
    CN308 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9887 downto 9856 ) ,
        VN2CN_bit   => CN_data_in( 9887 downto 9856 ) ,
        CN2VN_sign  => CN_sign_temp( 9887 downto 9856),
        CN2VN_bit   => CN_data_temp( 9887 downto 9856)
    );
    CN309 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9919 downto 9888 ) ,
        VN2CN_bit   => CN_data_in( 9919 downto 9888 ) ,
        CN2VN_sign  => CN_sign_temp( 9919 downto 9888),
        CN2VN_bit   => CN_data_temp( 9919 downto 9888)
    );
    CN310 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9951 downto 9920 ) ,
        VN2CN_bit   => CN_data_in( 9951 downto 9920 ) ,
        CN2VN_sign  => CN_sign_temp( 9951 downto 9920),
        CN2VN_bit   => CN_data_temp( 9951 downto 9920)
    );
    CN311 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 9983 downto 9952 ) ,
        VN2CN_bit   => CN_data_in( 9983 downto 9952 ) ,
        CN2VN_sign  => CN_sign_temp( 9983 downto 9952),
        CN2VN_bit   => CN_data_temp( 9983 downto 9952)
    );
    CN312 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10015 downto 9984 ) ,
        VN2CN_bit   => CN_data_in( 10015 downto 9984 ) ,
        CN2VN_sign  => CN_sign_temp( 10015 downto 9984),
        CN2VN_bit   => CN_data_temp( 10015 downto 9984)
    );
    CN313 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10047 downto 10016 ) ,
        VN2CN_bit   => CN_data_in( 10047 downto 10016 ) ,
        CN2VN_sign  => CN_sign_temp( 10047 downto 10016),
        CN2VN_bit   => CN_data_temp( 10047 downto 10016)
    );
    CN314 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10079 downto 10048 ) ,
        VN2CN_bit   => CN_data_in( 10079 downto 10048 ) ,
        CN2VN_sign  => CN_sign_temp( 10079 downto 10048),
        CN2VN_bit   => CN_data_temp( 10079 downto 10048)
    );
    CN315 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10111 downto 10080 ) ,
        VN2CN_bit   => CN_data_in( 10111 downto 10080 ) ,
        CN2VN_sign  => CN_sign_temp( 10111 downto 10080),
        CN2VN_bit   => CN_data_temp( 10111 downto 10080)
    );
    CN316 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10143 downto 10112 ) ,
        VN2CN_bit   => CN_data_in( 10143 downto 10112 ) ,
        CN2VN_sign  => CN_sign_temp( 10143 downto 10112),
        CN2VN_bit   => CN_data_temp( 10143 downto 10112)
    );
    CN317 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10175 downto 10144 ) ,
        VN2CN_bit   => CN_data_in( 10175 downto 10144 ) ,
        CN2VN_sign  => CN_sign_temp( 10175 downto 10144),
        CN2VN_bit   => CN_data_temp( 10175 downto 10144)
    );
    CN318 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10207 downto 10176 ) ,
        VN2CN_bit   => CN_data_in( 10207 downto 10176 ) ,
        CN2VN_sign  => CN_sign_temp( 10207 downto 10176),
        CN2VN_bit   => CN_data_temp( 10207 downto 10176)
    );
    CN319 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10239 downto 10208 ) ,
        VN2CN_bit   => CN_data_in( 10239 downto 10208 ) ,
        CN2VN_sign  => CN_sign_temp( 10239 downto 10208),
        CN2VN_bit   => CN_data_temp( 10239 downto 10208)
    );
    CN320 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10271 downto 10240 ) ,
        VN2CN_bit   => CN_data_in( 10271 downto 10240 ) ,
        CN2VN_sign  => CN_sign_temp( 10271 downto 10240),
        CN2VN_bit   => CN_data_temp( 10271 downto 10240)
    );
    CN321 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10303 downto 10272 ) ,
        VN2CN_bit   => CN_data_in( 10303 downto 10272 ) ,
        CN2VN_sign  => CN_sign_temp( 10303 downto 10272),
        CN2VN_bit   => CN_data_temp( 10303 downto 10272)
    );
    CN322 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10335 downto 10304 ) ,
        VN2CN_bit   => CN_data_in( 10335 downto 10304 ) ,
        CN2VN_sign  => CN_sign_temp( 10335 downto 10304),
        CN2VN_bit   => CN_data_temp( 10335 downto 10304)
    );
    CN323 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10367 downto 10336 ) ,
        VN2CN_bit   => CN_data_in( 10367 downto 10336 ) ,
        CN2VN_sign  => CN_sign_temp( 10367 downto 10336),
        CN2VN_bit   => CN_data_temp( 10367 downto 10336)
    );
    CN324 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10399 downto 10368 ) ,
        VN2CN_bit   => CN_data_in( 10399 downto 10368 ) ,
        CN2VN_sign  => CN_sign_temp( 10399 downto 10368),
        CN2VN_bit   => CN_data_temp( 10399 downto 10368)
    );
    CN325 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10431 downto 10400 ) ,
        VN2CN_bit   => CN_data_in( 10431 downto 10400 ) ,
        CN2VN_sign  => CN_sign_temp( 10431 downto 10400),
        CN2VN_bit   => CN_data_temp( 10431 downto 10400)
    );
    CN326 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10463 downto 10432 ) ,
        VN2CN_bit   => CN_data_in( 10463 downto 10432 ) ,
        CN2VN_sign  => CN_sign_temp( 10463 downto 10432),
        CN2VN_bit   => CN_data_temp( 10463 downto 10432)
    );
    CN327 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10495 downto 10464 ) ,
        VN2CN_bit   => CN_data_in( 10495 downto 10464 ) ,
        CN2VN_sign  => CN_sign_temp( 10495 downto 10464),
        CN2VN_bit   => CN_data_temp( 10495 downto 10464)
    );
    CN328 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10527 downto 10496 ) ,
        VN2CN_bit   => CN_data_in( 10527 downto 10496 ) ,
        CN2VN_sign  => CN_sign_temp( 10527 downto 10496),
        CN2VN_bit   => CN_data_temp( 10527 downto 10496)
    );
    CN329 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10559 downto 10528 ) ,
        VN2CN_bit   => CN_data_in( 10559 downto 10528 ) ,
        CN2VN_sign  => CN_sign_temp( 10559 downto 10528),
        CN2VN_bit   => CN_data_temp( 10559 downto 10528)
    );
    CN330 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10591 downto 10560 ) ,
        VN2CN_bit   => CN_data_in( 10591 downto 10560 ) ,
        CN2VN_sign  => CN_sign_temp( 10591 downto 10560),
        CN2VN_bit   => CN_data_temp( 10591 downto 10560)
    );
    CN331 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10623 downto 10592 ) ,
        VN2CN_bit   => CN_data_in( 10623 downto 10592 ) ,
        CN2VN_sign  => CN_sign_temp( 10623 downto 10592),
        CN2VN_bit   => CN_data_temp( 10623 downto 10592)
    );
    CN332 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10655 downto 10624 ) ,
        VN2CN_bit   => CN_data_in( 10655 downto 10624 ) ,
        CN2VN_sign  => CN_sign_temp( 10655 downto 10624),
        CN2VN_bit   => CN_data_temp( 10655 downto 10624)
    );
    CN333 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10687 downto 10656 ) ,
        VN2CN_bit   => CN_data_in( 10687 downto 10656 ) ,
        CN2VN_sign  => CN_sign_temp( 10687 downto 10656),
        CN2VN_bit   => CN_data_temp( 10687 downto 10656)
    );
    CN334 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10719 downto 10688 ) ,
        VN2CN_bit   => CN_data_in( 10719 downto 10688 ) ,
        CN2VN_sign  => CN_sign_temp( 10719 downto 10688),
        CN2VN_bit   => CN_data_temp( 10719 downto 10688)
    );
    CN335 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10751 downto 10720 ) ,
        VN2CN_bit   => CN_data_in( 10751 downto 10720 ) ,
        CN2VN_sign  => CN_sign_temp( 10751 downto 10720),
        CN2VN_bit   => CN_data_temp( 10751 downto 10720)
    );
    CN336 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10783 downto 10752 ) ,
        VN2CN_bit   => CN_data_in( 10783 downto 10752 ) ,
        CN2VN_sign  => CN_sign_temp( 10783 downto 10752),
        CN2VN_bit   => CN_data_temp( 10783 downto 10752)
    );
    CN337 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10815 downto 10784 ) ,
        VN2CN_bit   => CN_data_in( 10815 downto 10784 ) ,
        CN2VN_sign  => CN_sign_temp( 10815 downto 10784),
        CN2VN_bit   => CN_data_temp( 10815 downto 10784)
    );
    CN338 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10847 downto 10816 ) ,
        VN2CN_bit   => CN_data_in( 10847 downto 10816 ) ,
        CN2VN_sign  => CN_sign_temp( 10847 downto 10816),
        CN2VN_bit   => CN_data_temp( 10847 downto 10816)
    );
    CN339 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10879 downto 10848 ) ,
        VN2CN_bit   => CN_data_in( 10879 downto 10848 ) ,
        CN2VN_sign  => CN_sign_temp( 10879 downto 10848),
        CN2VN_bit   => CN_data_temp( 10879 downto 10848)
    );
    CN340 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10911 downto 10880 ) ,
        VN2CN_bit   => CN_data_in( 10911 downto 10880 ) ,
        CN2VN_sign  => CN_sign_temp( 10911 downto 10880),
        CN2VN_bit   => CN_data_temp( 10911 downto 10880)
    );
    CN341 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10943 downto 10912 ) ,
        VN2CN_bit   => CN_data_in( 10943 downto 10912 ) ,
        CN2VN_sign  => CN_sign_temp( 10943 downto 10912),
        CN2VN_bit   => CN_data_temp( 10943 downto 10912)
    );
    CN342 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 10975 downto 10944 ) ,
        VN2CN_bit   => CN_data_in( 10975 downto 10944 ) ,
        CN2VN_sign  => CN_sign_temp( 10975 downto 10944),
        CN2VN_bit   => CN_data_temp( 10975 downto 10944)
    );
    CN343 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11007 downto 10976 ) ,
        VN2CN_bit   => CN_data_in( 11007 downto 10976 ) ,
        CN2VN_sign  => CN_sign_temp( 11007 downto 10976),
        CN2VN_bit   => CN_data_temp( 11007 downto 10976)
    );
    CN344 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11039 downto 11008 ) ,
        VN2CN_bit   => CN_data_in( 11039 downto 11008 ) ,
        CN2VN_sign  => CN_sign_temp( 11039 downto 11008),
        CN2VN_bit   => CN_data_temp( 11039 downto 11008)
    );
    CN345 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11071 downto 11040 ) ,
        VN2CN_bit   => CN_data_in( 11071 downto 11040 ) ,
        CN2VN_sign  => CN_sign_temp( 11071 downto 11040),
        CN2VN_bit   => CN_data_temp( 11071 downto 11040)
    );
    CN346 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11103 downto 11072 ) ,
        VN2CN_bit   => CN_data_in( 11103 downto 11072 ) ,
        CN2VN_sign  => CN_sign_temp( 11103 downto 11072),
        CN2VN_bit   => CN_data_temp( 11103 downto 11072)
    );
    CN347 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11135 downto 11104 ) ,
        VN2CN_bit   => CN_data_in( 11135 downto 11104 ) ,
        CN2VN_sign  => CN_sign_temp( 11135 downto 11104),
        CN2VN_bit   => CN_data_temp( 11135 downto 11104)
    );
    CN348 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11167 downto 11136 ) ,
        VN2CN_bit   => CN_data_in( 11167 downto 11136 ) ,
        CN2VN_sign  => CN_sign_temp( 11167 downto 11136),
        CN2VN_bit   => CN_data_temp( 11167 downto 11136)
    );
    CN349 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11199 downto 11168 ) ,
        VN2CN_bit   => CN_data_in( 11199 downto 11168 ) ,
        CN2VN_sign  => CN_sign_temp( 11199 downto 11168),
        CN2VN_bit   => CN_data_temp( 11199 downto 11168)
    );
    CN350 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11231 downto 11200 ) ,
        VN2CN_bit   => CN_data_in( 11231 downto 11200 ) ,
        CN2VN_sign  => CN_sign_temp( 11231 downto 11200),
        CN2VN_bit   => CN_data_temp( 11231 downto 11200)
    );
    CN351 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11263 downto 11232 ) ,
        VN2CN_bit   => CN_data_in( 11263 downto 11232 ) ,
        CN2VN_sign  => CN_sign_temp( 11263 downto 11232),
        CN2VN_bit   => CN_data_temp( 11263 downto 11232)
    );
    CN352 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11295 downto 11264 ) ,
        VN2CN_bit   => CN_data_in( 11295 downto 11264 ) ,
        CN2VN_sign  => CN_sign_temp( 11295 downto 11264),
        CN2VN_bit   => CN_data_temp( 11295 downto 11264)
    );
    CN353 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11327 downto 11296 ) ,
        VN2CN_bit   => CN_data_in( 11327 downto 11296 ) ,
        CN2VN_sign  => CN_sign_temp( 11327 downto 11296),
        CN2VN_bit   => CN_data_temp( 11327 downto 11296)
    );
    CN354 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11359 downto 11328 ) ,
        VN2CN_bit   => CN_data_in( 11359 downto 11328 ) ,
        CN2VN_sign  => CN_sign_temp( 11359 downto 11328),
        CN2VN_bit   => CN_data_temp( 11359 downto 11328)
    );
    CN355 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11391 downto 11360 ) ,
        VN2CN_bit   => CN_data_in( 11391 downto 11360 ) ,
        CN2VN_sign  => CN_sign_temp( 11391 downto 11360),
        CN2VN_bit   => CN_data_temp( 11391 downto 11360)
    );
    CN356 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11423 downto 11392 ) ,
        VN2CN_bit   => CN_data_in( 11423 downto 11392 ) ,
        CN2VN_sign  => CN_sign_temp( 11423 downto 11392),
        CN2VN_bit   => CN_data_temp( 11423 downto 11392)
    );
    CN357 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11455 downto 11424 ) ,
        VN2CN_bit   => CN_data_in( 11455 downto 11424 ) ,
        CN2VN_sign  => CN_sign_temp( 11455 downto 11424),
        CN2VN_bit   => CN_data_temp( 11455 downto 11424)
    );
    CN358 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11487 downto 11456 ) ,
        VN2CN_bit   => CN_data_in( 11487 downto 11456 ) ,
        CN2VN_sign  => CN_sign_temp( 11487 downto 11456),
        CN2VN_bit   => CN_data_temp( 11487 downto 11456)
    );
    CN359 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11519 downto 11488 ) ,
        VN2CN_bit   => CN_data_in( 11519 downto 11488 ) ,
        CN2VN_sign  => CN_sign_temp( 11519 downto 11488),
        CN2VN_bit   => CN_data_temp( 11519 downto 11488)
    );
    CN360 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11551 downto 11520 ) ,
        VN2CN_bit   => CN_data_in( 11551 downto 11520 ) ,
        CN2VN_sign  => CN_sign_temp( 11551 downto 11520),
        CN2VN_bit   => CN_data_temp( 11551 downto 11520)
    );
    CN361 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11583 downto 11552 ) ,
        VN2CN_bit   => CN_data_in( 11583 downto 11552 ) ,
        CN2VN_sign  => CN_sign_temp( 11583 downto 11552),
        CN2VN_bit   => CN_data_temp( 11583 downto 11552)
    );
    CN362 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11615 downto 11584 ) ,
        VN2CN_bit   => CN_data_in( 11615 downto 11584 ) ,
        CN2VN_sign  => CN_sign_temp( 11615 downto 11584),
        CN2VN_bit   => CN_data_temp( 11615 downto 11584)
    );
    CN363 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11647 downto 11616 ) ,
        VN2CN_bit   => CN_data_in( 11647 downto 11616 ) ,
        CN2VN_sign  => CN_sign_temp( 11647 downto 11616),
        CN2VN_bit   => CN_data_temp( 11647 downto 11616)
    );
    CN364 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11679 downto 11648 ) ,
        VN2CN_bit   => CN_data_in( 11679 downto 11648 ) ,
        CN2VN_sign  => CN_sign_temp( 11679 downto 11648),
        CN2VN_bit   => CN_data_temp( 11679 downto 11648)
    );
    CN365 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11711 downto 11680 ) ,
        VN2CN_bit   => CN_data_in( 11711 downto 11680 ) ,
        CN2VN_sign  => CN_sign_temp( 11711 downto 11680),
        CN2VN_bit   => CN_data_temp( 11711 downto 11680)
    );
    CN366 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11743 downto 11712 ) ,
        VN2CN_bit   => CN_data_in( 11743 downto 11712 ) ,
        CN2VN_sign  => CN_sign_temp( 11743 downto 11712),
        CN2VN_bit   => CN_data_temp( 11743 downto 11712)
    );
    CN367 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11775 downto 11744 ) ,
        VN2CN_bit   => CN_data_in( 11775 downto 11744 ) ,
        CN2VN_sign  => CN_sign_temp( 11775 downto 11744),
        CN2VN_bit   => CN_data_temp( 11775 downto 11744)
    );
    CN368 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11807 downto 11776 ) ,
        VN2CN_bit   => CN_data_in( 11807 downto 11776 ) ,
        CN2VN_sign  => CN_sign_temp( 11807 downto 11776),
        CN2VN_bit   => CN_data_temp( 11807 downto 11776)
    );
    CN369 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11839 downto 11808 ) ,
        VN2CN_bit   => CN_data_in( 11839 downto 11808 ) ,
        CN2VN_sign  => CN_sign_temp( 11839 downto 11808),
        CN2VN_bit   => CN_data_temp( 11839 downto 11808)
    );
    CN370 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11871 downto 11840 ) ,
        VN2CN_bit   => CN_data_in( 11871 downto 11840 ) ,
        CN2VN_sign  => CN_sign_temp( 11871 downto 11840),
        CN2VN_bit   => CN_data_temp( 11871 downto 11840)
    );
    CN371 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11903 downto 11872 ) ,
        VN2CN_bit   => CN_data_in( 11903 downto 11872 ) ,
        CN2VN_sign  => CN_sign_temp( 11903 downto 11872),
        CN2VN_bit   => CN_data_temp( 11903 downto 11872)
    );
    CN372 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11935 downto 11904 ) ,
        VN2CN_bit   => CN_data_in( 11935 downto 11904 ) ,
        CN2VN_sign  => CN_sign_temp( 11935 downto 11904),
        CN2VN_bit   => CN_data_temp( 11935 downto 11904)
    );
    CN373 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11967 downto 11936 ) ,
        VN2CN_bit   => CN_data_in( 11967 downto 11936 ) ,
        CN2VN_sign  => CN_sign_temp( 11967 downto 11936),
        CN2VN_bit   => CN_data_temp( 11967 downto 11936)
    );
    CN374 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 11999 downto 11968 ) ,
        VN2CN_bit   => CN_data_in( 11999 downto 11968 ) ,
        CN2VN_sign  => CN_sign_temp( 11999 downto 11968),
        CN2VN_bit   => CN_data_temp( 11999 downto 11968)
    );
    CN375 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12031 downto 12000 ) ,
        VN2CN_bit   => CN_data_in( 12031 downto 12000 ) ,
        CN2VN_sign  => CN_sign_temp( 12031 downto 12000),
        CN2VN_bit   => CN_data_temp( 12031 downto 12000)
    );
    CN376 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12063 downto 12032 ) ,
        VN2CN_bit   => CN_data_in( 12063 downto 12032 ) ,
        CN2VN_sign  => CN_sign_temp( 12063 downto 12032),
        CN2VN_bit   => CN_data_temp( 12063 downto 12032)
    );
    CN377 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12095 downto 12064 ) ,
        VN2CN_bit   => CN_data_in( 12095 downto 12064 ) ,
        CN2VN_sign  => CN_sign_temp( 12095 downto 12064),
        CN2VN_bit   => CN_data_temp( 12095 downto 12064)
    );
    CN378 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12127 downto 12096 ) ,
        VN2CN_bit   => CN_data_in( 12127 downto 12096 ) ,
        CN2VN_sign  => CN_sign_temp( 12127 downto 12096),
        CN2VN_bit   => CN_data_temp( 12127 downto 12096)
    );
    CN379 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12159 downto 12128 ) ,
        VN2CN_bit   => CN_data_in( 12159 downto 12128 ) ,
        CN2VN_sign  => CN_sign_temp( 12159 downto 12128),
        CN2VN_bit   => CN_data_temp( 12159 downto 12128)
    );
    CN380 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12191 downto 12160 ) ,
        VN2CN_bit   => CN_data_in( 12191 downto 12160 ) ,
        CN2VN_sign  => CN_sign_temp( 12191 downto 12160),
        CN2VN_bit   => CN_data_temp( 12191 downto 12160)
    );
    CN381 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12223 downto 12192 ) ,
        VN2CN_bit   => CN_data_in( 12223 downto 12192 ) ,
        CN2VN_sign  => CN_sign_temp( 12223 downto 12192),
        CN2VN_bit   => CN_data_temp( 12223 downto 12192)
    );
    CN382 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12255 downto 12224 ) ,
        VN2CN_bit   => CN_data_in( 12255 downto 12224 ) ,
        CN2VN_sign  => CN_sign_temp( 12255 downto 12224),
        CN2VN_bit   => CN_data_temp( 12255 downto 12224)
    );
    CN383 : CN_Dv32 port map(
        VN2CN_sign  => CN_sign_in( 12287 downto 12256 ) ,
        VN2CN_bit   => CN_data_in( 12287 downto 12256 ) ,
        CN2VN_sign  => CN_sign_temp( 12287 downto 12256),
        CN2VN_bit   => CN_data_temp( 12287 downto 12256)
    );






end architecture ; -- arch