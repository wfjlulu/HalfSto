library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity VNUpdate is
  port (
    clk :         in std_logic;
    rst_n :       in std_logic;
    LLR :         in std_logic_vector(12287 downto 0);  --2048*6 = 12288
    VN_data_in :  in std_logic_vector(12287 downto 0);--2048*6 = 12288
    VN_sign_in :  in std_logic_vector(12287 downto 0);
    RandomNum :   in std_logic_vector(3 downto 0);
    New_LLR   :   in std_logic;
    DecoderOver : in std_logic;
    --DV_in :       in std_logic;
    VN_data_out : out std_logic_vector(12287 downto 0);
    VN_sign_out : out std_logic_vector(12287 downto 0);
    codeword :    out std_logic_vector(0 to 2047);
    Iterations :  inout std_logic_vector(4 downto 0);
    DV_out :      out std_logic;
    DecodeState : out std_logic_vector( 1 downto 0 )
  ) ;
end VNUpdate ;

architecture arch of VNUpdate is
    component VN_Dv6 is
        port(
            clk : in std_logic;
            rst_n : in std_logic;
            New_LLR : in std_logic;
            DecoderOver : in std_logic;
            --DV_in : in std_logic;
            RandomNum : in std_logic_vector( 3 downto 0 ); --unsigned number
            LLR  : in std_logic_vector( 5 downto 0);  -- input LLR is 5 bits signed number +-15
            Din0 : in std_logic_vector( 1 downto 0);  -- one bit for sign 4 bits for AM 
            Din1 : in std_logic_vector( 1 downto 0);
            Din2 : in std_logic_vector( 1 downto 0);
            Din3 : in std_logic_vector( 1 downto 0);
            Din4 : in std_logic_vector( 1 downto 0);
            Din5 : in std_logic_vector( 1 downto 0);
            VN2CN0_bit : out std_logic;
            VN2CN1_bit : out std_logic;
            VN2CN2_bit : out std_logic;
            VN2CN3_bit : out std_logic;
            VN2CN4_bit : out std_logic;
            VN2CN5_bit : out std_logic;
            VN2CN0_sign : out std_logic;
            VN2CN1_sign : out std_logic;
            VN2CN2_sign : out std_logic;
            VN2CN3_sign : out std_logic;
            VN2CN4_sign : out std_logic;
            VN2CN5_sign : out std_logic;
    
            codeword    : out std_logic;
            Iterations  : inout std_logic_vector(4 downto 0 );
    
            DV_out : out std_logic;  -- data valid flag
            DecodeState : out std_logic_vector( 1 downto 0 )
        );
    end component;
    
    signal VN0_in0 : std_logic_vector(1 downto 0);
    signal VN0_in1 : std_logic_vector(1 downto 0);
    signal VN0_in2 : std_logic_vector(1 downto 0);
    signal VN0_in3 : std_logic_vector(1 downto 0);
    signal VN0_in4 : std_logic_vector(1 downto 0);
    signal VN0_in5 : std_logic_vector(1 downto 0);

    signal VN1_in0 : std_logic_vector(1 downto 0);
    signal VN1_in1 : std_logic_vector(1 downto 0);
    signal VN1_in2 : std_logic_vector(1 downto 0);
    signal VN1_in3 : std_logic_vector(1 downto 0);
    signal VN1_in4 : std_logic_vector(1 downto 0);
    signal VN1_in5 : std_logic_vector(1 downto 0);
    signal VN2_in0 : std_logic_vector(1 downto 0);
    signal VN2_in1 : std_logic_vector(1 downto 0);
    signal VN2_in2 : std_logic_vector(1 downto 0);
    signal VN2_in3 : std_logic_vector(1 downto 0);
    signal VN2_in4 : std_logic_vector(1 downto 0);
    signal VN2_in5 : std_logic_vector(1 downto 0);
    signal VN3_in0 : std_logic_vector(1 downto 0);
    signal VN3_in1 : std_logic_vector(1 downto 0);
    signal VN3_in2 : std_logic_vector(1 downto 0);
    signal VN3_in3 : std_logic_vector(1 downto 0);
    signal VN3_in4 : std_logic_vector(1 downto 0);
    signal VN3_in5 : std_logic_vector(1 downto 0);
    signal VN4_in0 : std_logic_vector(1 downto 0);
    signal VN4_in1 : std_logic_vector(1 downto 0);
    signal VN4_in2 : std_logic_vector(1 downto 0);
    signal VN4_in3 : std_logic_vector(1 downto 0);
    signal VN4_in4 : std_logic_vector(1 downto 0);
    signal VN4_in5 : std_logic_vector(1 downto 0);
    signal VN5_in0 : std_logic_vector(1 downto 0);
    signal VN5_in1 : std_logic_vector(1 downto 0);
    signal VN5_in2 : std_logic_vector(1 downto 0);
    signal VN5_in3 : std_logic_vector(1 downto 0);
    signal VN5_in4 : std_logic_vector(1 downto 0);
    signal VN5_in5 : std_logic_vector(1 downto 0);
    signal VN6_in0 : std_logic_vector(1 downto 0);
    signal VN6_in1 : std_logic_vector(1 downto 0);
    signal VN6_in2 : std_logic_vector(1 downto 0);
    signal VN6_in3 : std_logic_vector(1 downto 0);
    signal VN6_in4 : std_logic_vector(1 downto 0);
    signal VN6_in5 : std_logic_vector(1 downto 0);
    signal VN7_in0 : std_logic_vector(1 downto 0);
    signal VN7_in1 : std_logic_vector(1 downto 0);
    signal VN7_in2 : std_logic_vector(1 downto 0);
    signal VN7_in3 : std_logic_vector(1 downto 0);
    signal VN7_in4 : std_logic_vector(1 downto 0);
    signal VN7_in5 : std_logic_vector(1 downto 0);
    signal VN8_in0 : std_logic_vector(1 downto 0);
    signal VN8_in1 : std_logic_vector(1 downto 0);
    signal VN8_in2 : std_logic_vector(1 downto 0);
    signal VN8_in3 : std_logic_vector(1 downto 0);
    signal VN8_in4 : std_logic_vector(1 downto 0);
    signal VN8_in5 : std_logic_vector(1 downto 0);
    signal VN9_in0 : std_logic_vector(1 downto 0);
    signal VN9_in1 : std_logic_vector(1 downto 0);
    signal VN9_in2 : std_logic_vector(1 downto 0);
    signal VN9_in3 : std_logic_vector(1 downto 0);
    signal VN9_in4 : std_logic_vector(1 downto 0);
    signal VN9_in5 : std_logic_vector(1 downto 0);
    signal VN10_in0 : std_logic_vector(1 downto 0);
    signal VN10_in1 : std_logic_vector(1 downto 0);
    signal VN10_in2 : std_logic_vector(1 downto 0);
    signal VN10_in3 : std_logic_vector(1 downto 0);
    signal VN10_in4 : std_logic_vector(1 downto 0);
    signal VN10_in5 : std_logic_vector(1 downto 0);
    signal VN11_in0 : std_logic_vector(1 downto 0);
    signal VN11_in1 : std_logic_vector(1 downto 0);
    signal VN11_in2 : std_logic_vector(1 downto 0);
    signal VN11_in3 : std_logic_vector(1 downto 0);
    signal VN11_in4 : std_logic_vector(1 downto 0);
    signal VN11_in5 : std_logic_vector(1 downto 0);
    signal VN12_in0 : std_logic_vector(1 downto 0);
    signal VN12_in1 : std_logic_vector(1 downto 0);
    signal VN12_in2 : std_logic_vector(1 downto 0);
    signal VN12_in3 : std_logic_vector(1 downto 0);
    signal VN12_in4 : std_logic_vector(1 downto 0);
    signal VN12_in5 : std_logic_vector(1 downto 0);
    signal VN13_in0 : std_logic_vector(1 downto 0);
    signal VN13_in1 : std_logic_vector(1 downto 0);
    signal VN13_in2 : std_logic_vector(1 downto 0);
    signal VN13_in3 : std_logic_vector(1 downto 0);
    signal VN13_in4 : std_logic_vector(1 downto 0);
    signal VN13_in5 : std_logic_vector(1 downto 0);
    signal VN14_in0 : std_logic_vector(1 downto 0);
    signal VN14_in1 : std_logic_vector(1 downto 0);
    signal VN14_in2 : std_logic_vector(1 downto 0);
    signal VN14_in3 : std_logic_vector(1 downto 0);
    signal VN14_in4 : std_logic_vector(1 downto 0);
    signal VN14_in5 : std_logic_vector(1 downto 0);
    signal VN15_in0 : std_logic_vector(1 downto 0);
    signal VN15_in1 : std_logic_vector(1 downto 0);
    signal VN15_in2 : std_logic_vector(1 downto 0);
    signal VN15_in3 : std_logic_vector(1 downto 0);
    signal VN15_in4 : std_logic_vector(1 downto 0);
    signal VN15_in5 : std_logic_vector(1 downto 0);
    signal VN16_in0 : std_logic_vector(1 downto 0);
    signal VN16_in1 : std_logic_vector(1 downto 0);
    signal VN16_in2 : std_logic_vector(1 downto 0);
    signal VN16_in3 : std_logic_vector(1 downto 0);
    signal VN16_in4 : std_logic_vector(1 downto 0);
    signal VN16_in5 : std_logic_vector(1 downto 0);
    signal VN17_in0 : std_logic_vector(1 downto 0);
    signal VN17_in1 : std_logic_vector(1 downto 0);
    signal VN17_in2 : std_logic_vector(1 downto 0);
    signal VN17_in3 : std_logic_vector(1 downto 0);
    signal VN17_in4 : std_logic_vector(1 downto 0);
    signal VN17_in5 : std_logic_vector(1 downto 0);
    signal VN18_in0 : std_logic_vector(1 downto 0);
    signal VN18_in1 : std_logic_vector(1 downto 0);
    signal VN18_in2 : std_logic_vector(1 downto 0);
    signal VN18_in3 : std_logic_vector(1 downto 0);
    signal VN18_in4 : std_logic_vector(1 downto 0);
    signal VN18_in5 : std_logic_vector(1 downto 0);
    signal VN19_in0 : std_logic_vector(1 downto 0);
    signal VN19_in1 : std_logic_vector(1 downto 0);
    signal VN19_in2 : std_logic_vector(1 downto 0);
    signal VN19_in3 : std_logic_vector(1 downto 0);
    signal VN19_in4 : std_logic_vector(1 downto 0);
    signal VN19_in5 : std_logic_vector(1 downto 0);
    signal VN20_in0 : std_logic_vector(1 downto 0);
    signal VN20_in1 : std_logic_vector(1 downto 0);
    signal VN20_in2 : std_logic_vector(1 downto 0);
    signal VN20_in3 : std_logic_vector(1 downto 0);
    signal VN20_in4 : std_logic_vector(1 downto 0);
    signal VN20_in5 : std_logic_vector(1 downto 0);
    signal VN21_in0 : std_logic_vector(1 downto 0);
    signal VN21_in1 : std_logic_vector(1 downto 0);
    signal VN21_in2 : std_logic_vector(1 downto 0);
    signal VN21_in3 : std_logic_vector(1 downto 0);
    signal VN21_in4 : std_logic_vector(1 downto 0);
    signal VN21_in5 : std_logic_vector(1 downto 0);
    signal VN22_in0 : std_logic_vector(1 downto 0);
    signal VN22_in1 : std_logic_vector(1 downto 0);
    signal VN22_in2 : std_logic_vector(1 downto 0);
    signal VN22_in3 : std_logic_vector(1 downto 0);
    signal VN22_in4 : std_logic_vector(1 downto 0);
    signal VN22_in5 : std_logic_vector(1 downto 0);
    signal VN23_in0 : std_logic_vector(1 downto 0);
    signal VN23_in1 : std_logic_vector(1 downto 0);
    signal VN23_in2 : std_logic_vector(1 downto 0);
    signal VN23_in3 : std_logic_vector(1 downto 0);
    signal VN23_in4 : std_logic_vector(1 downto 0);
    signal VN23_in5 : std_logic_vector(1 downto 0);
    signal VN24_in0 : std_logic_vector(1 downto 0);
    signal VN24_in1 : std_logic_vector(1 downto 0);
    signal VN24_in2 : std_logic_vector(1 downto 0);
    signal VN24_in3 : std_logic_vector(1 downto 0);
    signal VN24_in4 : std_logic_vector(1 downto 0);
    signal VN24_in5 : std_logic_vector(1 downto 0);
    signal VN25_in0 : std_logic_vector(1 downto 0);
    signal VN25_in1 : std_logic_vector(1 downto 0);
    signal VN25_in2 : std_logic_vector(1 downto 0);
    signal VN25_in3 : std_logic_vector(1 downto 0);
    signal VN25_in4 : std_logic_vector(1 downto 0);
    signal VN25_in5 : std_logic_vector(1 downto 0);
    signal VN26_in0 : std_logic_vector(1 downto 0);
    signal VN26_in1 : std_logic_vector(1 downto 0);
    signal VN26_in2 : std_logic_vector(1 downto 0);
    signal VN26_in3 : std_logic_vector(1 downto 0);
    signal VN26_in4 : std_logic_vector(1 downto 0);
    signal VN26_in5 : std_logic_vector(1 downto 0);
    signal VN27_in0 : std_logic_vector(1 downto 0);
    signal VN27_in1 : std_logic_vector(1 downto 0);
    signal VN27_in2 : std_logic_vector(1 downto 0);
    signal VN27_in3 : std_logic_vector(1 downto 0);
    signal VN27_in4 : std_logic_vector(1 downto 0);
    signal VN27_in5 : std_logic_vector(1 downto 0);
    signal VN28_in0 : std_logic_vector(1 downto 0);
    signal VN28_in1 : std_logic_vector(1 downto 0);
    signal VN28_in2 : std_logic_vector(1 downto 0);
    signal VN28_in3 : std_logic_vector(1 downto 0);
    signal VN28_in4 : std_logic_vector(1 downto 0);
    signal VN28_in5 : std_logic_vector(1 downto 0);
    signal VN29_in0 : std_logic_vector(1 downto 0);
    signal VN29_in1 : std_logic_vector(1 downto 0);
    signal VN29_in2 : std_logic_vector(1 downto 0);
    signal VN29_in3 : std_logic_vector(1 downto 0);
    signal VN29_in4 : std_logic_vector(1 downto 0);
    signal VN29_in5 : std_logic_vector(1 downto 0);
    signal VN30_in0 : std_logic_vector(1 downto 0);
    signal VN30_in1 : std_logic_vector(1 downto 0);
    signal VN30_in2 : std_logic_vector(1 downto 0);
    signal VN30_in3 : std_logic_vector(1 downto 0);
    signal VN30_in4 : std_logic_vector(1 downto 0);
    signal VN30_in5 : std_logic_vector(1 downto 0);
    signal VN31_in0 : std_logic_vector(1 downto 0);
    signal VN31_in1 : std_logic_vector(1 downto 0);
    signal VN31_in2 : std_logic_vector(1 downto 0);
    signal VN31_in3 : std_logic_vector(1 downto 0);
    signal VN31_in4 : std_logic_vector(1 downto 0);
    signal VN31_in5 : std_logic_vector(1 downto 0);
    signal VN32_in0 : std_logic_vector(1 downto 0);
    signal VN32_in1 : std_logic_vector(1 downto 0);
    signal VN32_in2 : std_logic_vector(1 downto 0);
    signal VN32_in3 : std_logic_vector(1 downto 0);
    signal VN32_in4 : std_logic_vector(1 downto 0);
    signal VN32_in5 : std_logic_vector(1 downto 0);
    signal VN33_in0 : std_logic_vector(1 downto 0);
    signal VN33_in1 : std_logic_vector(1 downto 0);
    signal VN33_in2 : std_logic_vector(1 downto 0);
    signal VN33_in3 : std_logic_vector(1 downto 0);
    signal VN33_in4 : std_logic_vector(1 downto 0);
    signal VN33_in5 : std_logic_vector(1 downto 0);
    signal VN34_in0 : std_logic_vector(1 downto 0);
    signal VN34_in1 : std_logic_vector(1 downto 0);
    signal VN34_in2 : std_logic_vector(1 downto 0);
    signal VN34_in3 : std_logic_vector(1 downto 0);
    signal VN34_in4 : std_logic_vector(1 downto 0);
    signal VN34_in5 : std_logic_vector(1 downto 0);
    signal VN35_in0 : std_logic_vector(1 downto 0);
    signal VN35_in1 : std_logic_vector(1 downto 0);
    signal VN35_in2 : std_logic_vector(1 downto 0);
    signal VN35_in3 : std_logic_vector(1 downto 0);
    signal VN35_in4 : std_logic_vector(1 downto 0);
    signal VN35_in5 : std_logic_vector(1 downto 0);
    signal VN36_in0 : std_logic_vector(1 downto 0);
    signal VN36_in1 : std_logic_vector(1 downto 0);
    signal VN36_in2 : std_logic_vector(1 downto 0);
    signal VN36_in3 : std_logic_vector(1 downto 0);
    signal VN36_in4 : std_logic_vector(1 downto 0);
    signal VN36_in5 : std_logic_vector(1 downto 0);
    signal VN37_in0 : std_logic_vector(1 downto 0);
    signal VN37_in1 : std_logic_vector(1 downto 0);
    signal VN37_in2 : std_logic_vector(1 downto 0);
    signal VN37_in3 : std_logic_vector(1 downto 0);
    signal VN37_in4 : std_logic_vector(1 downto 0);
    signal VN37_in5 : std_logic_vector(1 downto 0);
    signal VN38_in0 : std_logic_vector(1 downto 0);
    signal VN38_in1 : std_logic_vector(1 downto 0);
    signal VN38_in2 : std_logic_vector(1 downto 0);
    signal VN38_in3 : std_logic_vector(1 downto 0);
    signal VN38_in4 : std_logic_vector(1 downto 0);
    signal VN38_in5 : std_logic_vector(1 downto 0);
    signal VN39_in0 : std_logic_vector(1 downto 0);
    signal VN39_in1 : std_logic_vector(1 downto 0);
    signal VN39_in2 : std_logic_vector(1 downto 0);
    signal VN39_in3 : std_logic_vector(1 downto 0);
    signal VN39_in4 : std_logic_vector(1 downto 0);
    signal VN39_in5 : std_logic_vector(1 downto 0);
    signal VN40_in0 : std_logic_vector(1 downto 0);
    signal VN40_in1 : std_logic_vector(1 downto 0);
    signal VN40_in2 : std_logic_vector(1 downto 0);
    signal VN40_in3 : std_logic_vector(1 downto 0);
    signal VN40_in4 : std_logic_vector(1 downto 0);
    signal VN40_in5 : std_logic_vector(1 downto 0);
    signal VN41_in0 : std_logic_vector(1 downto 0);
    signal VN41_in1 : std_logic_vector(1 downto 0);
    signal VN41_in2 : std_logic_vector(1 downto 0);
    signal VN41_in3 : std_logic_vector(1 downto 0);
    signal VN41_in4 : std_logic_vector(1 downto 0);
    signal VN41_in5 : std_logic_vector(1 downto 0);
    signal VN42_in0 : std_logic_vector(1 downto 0);
    signal VN42_in1 : std_logic_vector(1 downto 0);
    signal VN42_in2 : std_logic_vector(1 downto 0);
    signal VN42_in3 : std_logic_vector(1 downto 0);
    signal VN42_in4 : std_logic_vector(1 downto 0);
    signal VN42_in5 : std_logic_vector(1 downto 0);
    signal VN43_in0 : std_logic_vector(1 downto 0);
    signal VN43_in1 : std_logic_vector(1 downto 0);
    signal VN43_in2 : std_logic_vector(1 downto 0);
    signal VN43_in3 : std_logic_vector(1 downto 0);
    signal VN43_in4 : std_logic_vector(1 downto 0);
    signal VN43_in5 : std_logic_vector(1 downto 0);
    signal VN44_in0 : std_logic_vector(1 downto 0);
    signal VN44_in1 : std_logic_vector(1 downto 0);
    signal VN44_in2 : std_logic_vector(1 downto 0);
    signal VN44_in3 : std_logic_vector(1 downto 0);
    signal VN44_in4 : std_logic_vector(1 downto 0);
    signal VN44_in5 : std_logic_vector(1 downto 0);
    signal VN45_in0 : std_logic_vector(1 downto 0);
    signal VN45_in1 : std_logic_vector(1 downto 0);
    signal VN45_in2 : std_logic_vector(1 downto 0);
    signal VN45_in3 : std_logic_vector(1 downto 0);
    signal VN45_in4 : std_logic_vector(1 downto 0);
    signal VN45_in5 : std_logic_vector(1 downto 0);
    signal VN46_in0 : std_logic_vector(1 downto 0);
    signal VN46_in1 : std_logic_vector(1 downto 0);
    signal VN46_in2 : std_logic_vector(1 downto 0);
    signal VN46_in3 : std_logic_vector(1 downto 0);
    signal VN46_in4 : std_logic_vector(1 downto 0);
    signal VN46_in5 : std_logic_vector(1 downto 0);
    signal VN47_in0 : std_logic_vector(1 downto 0);
    signal VN47_in1 : std_logic_vector(1 downto 0);
    signal VN47_in2 : std_logic_vector(1 downto 0);
    signal VN47_in3 : std_logic_vector(1 downto 0);
    signal VN47_in4 : std_logic_vector(1 downto 0);
    signal VN47_in5 : std_logic_vector(1 downto 0);
    signal VN48_in0 : std_logic_vector(1 downto 0);
    signal VN48_in1 : std_logic_vector(1 downto 0);
    signal VN48_in2 : std_logic_vector(1 downto 0);
    signal VN48_in3 : std_logic_vector(1 downto 0);
    signal VN48_in4 : std_logic_vector(1 downto 0);
    signal VN48_in5 : std_logic_vector(1 downto 0);
    signal VN49_in0 : std_logic_vector(1 downto 0);
    signal VN49_in1 : std_logic_vector(1 downto 0);
    signal VN49_in2 : std_logic_vector(1 downto 0);
    signal VN49_in3 : std_logic_vector(1 downto 0);
    signal VN49_in4 : std_logic_vector(1 downto 0);
    signal VN49_in5 : std_logic_vector(1 downto 0);
    signal VN50_in0 : std_logic_vector(1 downto 0);
    signal VN50_in1 : std_logic_vector(1 downto 0);
    signal VN50_in2 : std_logic_vector(1 downto 0);
    signal VN50_in3 : std_logic_vector(1 downto 0);
    signal VN50_in4 : std_logic_vector(1 downto 0);
    signal VN50_in5 : std_logic_vector(1 downto 0);
    signal VN51_in0 : std_logic_vector(1 downto 0);
    signal VN51_in1 : std_logic_vector(1 downto 0);
    signal VN51_in2 : std_logic_vector(1 downto 0);
    signal VN51_in3 : std_logic_vector(1 downto 0);
    signal VN51_in4 : std_logic_vector(1 downto 0);
    signal VN51_in5 : std_logic_vector(1 downto 0);
    signal VN52_in0 : std_logic_vector(1 downto 0);
    signal VN52_in1 : std_logic_vector(1 downto 0);
    signal VN52_in2 : std_logic_vector(1 downto 0);
    signal VN52_in3 : std_logic_vector(1 downto 0);
    signal VN52_in4 : std_logic_vector(1 downto 0);
    signal VN52_in5 : std_logic_vector(1 downto 0);
    signal VN53_in0 : std_logic_vector(1 downto 0);
    signal VN53_in1 : std_logic_vector(1 downto 0);
    signal VN53_in2 : std_logic_vector(1 downto 0);
    signal VN53_in3 : std_logic_vector(1 downto 0);
    signal VN53_in4 : std_logic_vector(1 downto 0);
    signal VN53_in5 : std_logic_vector(1 downto 0);
    signal VN54_in0 : std_logic_vector(1 downto 0);
    signal VN54_in1 : std_logic_vector(1 downto 0);
    signal VN54_in2 : std_logic_vector(1 downto 0);
    signal VN54_in3 : std_logic_vector(1 downto 0);
    signal VN54_in4 : std_logic_vector(1 downto 0);
    signal VN54_in5 : std_logic_vector(1 downto 0);
    signal VN55_in0 : std_logic_vector(1 downto 0);
    signal VN55_in1 : std_logic_vector(1 downto 0);
    signal VN55_in2 : std_logic_vector(1 downto 0);
    signal VN55_in3 : std_logic_vector(1 downto 0);
    signal VN55_in4 : std_logic_vector(1 downto 0);
    signal VN55_in5 : std_logic_vector(1 downto 0);
    signal VN56_in0 : std_logic_vector(1 downto 0);
    signal VN56_in1 : std_logic_vector(1 downto 0);
    signal VN56_in2 : std_logic_vector(1 downto 0);
    signal VN56_in3 : std_logic_vector(1 downto 0);
    signal VN56_in4 : std_logic_vector(1 downto 0);
    signal VN56_in5 : std_logic_vector(1 downto 0);
    signal VN57_in0 : std_logic_vector(1 downto 0);
    signal VN57_in1 : std_logic_vector(1 downto 0);
    signal VN57_in2 : std_logic_vector(1 downto 0);
    signal VN57_in3 : std_logic_vector(1 downto 0);
    signal VN57_in4 : std_logic_vector(1 downto 0);
    signal VN57_in5 : std_logic_vector(1 downto 0);
    signal VN58_in0 : std_logic_vector(1 downto 0);
    signal VN58_in1 : std_logic_vector(1 downto 0);
    signal VN58_in2 : std_logic_vector(1 downto 0);
    signal VN58_in3 : std_logic_vector(1 downto 0);
    signal VN58_in4 : std_logic_vector(1 downto 0);
    signal VN58_in5 : std_logic_vector(1 downto 0);
    signal VN59_in0 : std_logic_vector(1 downto 0);
    signal VN59_in1 : std_logic_vector(1 downto 0);
    signal VN59_in2 : std_logic_vector(1 downto 0);
    signal VN59_in3 : std_logic_vector(1 downto 0);
    signal VN59_in4 : std_logic_vector(1 downto 0);
    signal VN59_in5 : std_logic_vector(1 downto 0);
    signal VN60_in0 : std_logic_vector(1 downto 0);
    signal VN60_in1 : std_logic_vector(1 downto 0);
    signal VN60_in2 : std_logic_vector(1 downto 0);
    signal VN60_in3 : std_logic_vector(1 downto 0);
    signal VN60_in4 : std_logic_vector(1 downto 0);
    signal VN60_in5 : std_logic_vector(1 downto 0);
    signal VN61_in0 : std_logic_vector(1 downto 0);
    signal VN61_in1 : std_logic_vector(1 downto 0);
    signal VN61_in2 : std_logic_vector(1 downto 0);
    signal VN61_in3 : std_logic_vector(1 downto 0);
    signal VN61_in4 : std_logic_vector(1 downto 0);
    signal VN61_in5 : std_logic_vector(1 downto 0);
    signal VN62_in0 : std_logic_vector(1 downto 0);
    signal VN62_in1 : std_logic_vector(1 downto 0);
    signal VN62_in2 : std_logic_vector(1 downto 0);
    signal VN62_in3 : std_logic_vector(1 downto 0);
    signal VN62_in4 : std_logic_vector(1 downto 0);
    signal VN62_in5 : std_logic_vector(1 downto 0);
    signal VN63_in0 : std_logic_vector(1 downto 0);
    signal VN63_in1 : std_logic_vector(1 downto 0);
    signal VN63_in2 : std_logic_vector(1 downto 0);
    signal VN63_in3 : std_logic_vector(1 downto 0);
    signal VN63_in4 : std_logic_vector(1 downto 0);
    signal VN63_in5 : std_logic_vector(1 downto 0);
    signal VN64_in0 : std_logic_vector(1 downto 0);
    signal VN64_in1 : std_logic_vector(1 downto 0);
    signal VN64_in2 : std_logic_vector(1 downto 0);
    signal VN64_in3 : std_logic_vector(1 downto 0);
    signal VN64_in4 : std_logic_vector(1 downto 0);
    signal VN64_in5 : std_logic_vector(1 downto 0);
    signal VN65_in0 : std_logic_vector(1 downto 0);
    signal VN65_in1 : std_logic_vector(1 downto 0);
    signal VN65_in2 : std_logic_vector(1 downto 0);
    signal VN65_in3 : std_logic_vector(1 downto 0);
    signal VN65_in4 : std_logic_vector(1 downto 0);
    signal VN65_in5 : std_logic_vector(1 downto 0);
    signal VN66_in0 : std_logic_vector(1 downto 0);
    signal VN66_in1 : std_logic_vector(1 downto 0);
    signal VN66_in2 : std_logic_vector(1 downto 0);
    signal VN66_in3 : std_logic_vector(1 downto 0);
    signal VN66_in4 : std_logic_vector(1 downto 0);
    signal VN66_in5 : std_logic_vector(1 downto 0);
    signal VN67_in0 : std_logic_vector(1 downto 0);
    signal VN67_in1 : std_logic_vector(1 downto 0);
    signal VN67_in2 : std_logic_vector(1 downto 0);
    signal VN67_in3 : std_logic_vector(1 downto 0);
    signal VN67_in4 : std_logic_vector(1 downto 0);
    signal VN67_in5 : std_logic_vector(1 downto 0);
    signal VN68_in0 : std_logic_vector(1 downto 0);
    signal VN68_in1 : std_logic_vector(1 downto 0);
    signal VN68_in2 : std_logic_vector(1 downto 0);
    signal VN68_in3 : std_logic_vector(1 downto 0);
    signal VN68_in4 : std_logic_vector(1 downto 0);
    signal VN68_in5 : std_logic_vector(1 downto 0);
    signal VN69_in0 : std_logic_vector(1 downto 0);
    signal VN69_in1 : std_logic_vector(1 downto 0);
    signal VN69_in2 : std_logic_vector(1 downto 0);
    signal VN69_in3 : std_logic_vector(1 downto 0);
    signal VN69_in4 : std_logic_vector(1 downto 0);
    signal VN69_in5 : std_logic_vector(1 downto 0);
    signal VN70_in0 : std_logic_vector(1 downto 0);
    signal VN70_in1 : std_logic_vector(1 downto 0);
    signal VN70_in2 : std_logic_vector(1 downto 0);
    signal VN70_in3 : std_logic_vector(1 downto 0);
    signal VN70_in4 : std_logic_vector(1 downto 0);
    signal VN70_in5 : std_logic_vector(1 downto 0);
    signal VN71_in0 : std_logic_vector(1 downto 0);
    signal VN71_in1 : std_logic_vector(1 downto 0);
    signal VN71_in2 : std_logic_vector(1 downto 0);
    signal VN71_in3 : std_logic_vector(1 downto 0);
    signal VN71_in4 : std_logic_vector(1 downto 0);
    signal VN71_in5 : std_logic_vector(1 downto 0);
    signal VN72_in0 : std_logic_vector(1 downto 0);
    signal VN72_in1 : std_logic_vector(1 downto 0);
    signal VN72_in2 : std_logic_vector(1 downto 0);
    signal VN72_in3 : std_logic_vector(1 downto 0);
    signal VN72_in4 : std_logic_vector(1 downto 0);
    signal VN72_in5 : std_logic_vector(1 downto 0);
    signal VN73_in0 : std_logic_vector(1 downto 0);
    signal VN73_in1 : std_logic_vector(1 downto 0);
    signal VN73_in2 : std_logic_vector(1 downto 0);
    signal VN73_in3 : std_logic_vector(1 downto 0);
    signal VN73_in4 : std_logic_vector(1 downto 0);
    signal VN73_in5 : std_logic_vector(1 downto 0);
    signal VN74_in0 : std_logic_vector(1 downto 0);
    signal VN74_in1 : std_logic_vector(1 downto 0);
    signal VN74_in2 : std_logic_vector(1 downto 0);
    signal VN74_in3 : std_logic_vector(1 downto 0);
    signal VN74_in4 : std_logic_vector(1 downto 0);
    signal VN74_in5 : std_logic_vector(1 downto 0);
    signal VN75_in0 : std_logic_vector(1 downto 0);
    signal VN75_in1 : std_logic_vector(1 downto 0);
    signal VN75_in2 : std_logic_vector(1 downto 0);
    signal VN75_in3 : std_logic_vector(1 downto 0);
    signal VN75_in4 : std_logic_vector(1 downto 0);
    signal VN75_in5 : std_logic_vector(1 downto 0);
    signal VN76_in0 : std_logic_vector(1 downto 0);
    signal VN76_in1 : std_logic_vector(1 downto 0);
    signal VN76_in2 : std_logic_vector(1 downto 0);
    signal VN76_in3 : std_logic_vector(1 downto 0);
    signal VN76_in4 : std_logic_vector(1 downto 0);
    signal VN76_in5 : std_logic_vector(1 downto 0);
    signal VN77_in0 : std_logic_vector(1 downto 0);
    signal VN77_in1 : std_logic_vector(1 downto 0);
    signal VN77_in2 : std_logic_vector(1 downto 0);
    signal VN77_in3 : std_logic_vector(1 downto 0);
    signal VN77_in4 : std_logic_vector(1 downto 0);
    signal VN77_in5 : std_logic_vector(1 downto 0);
    signal VN78_in0 : std_logic_vector(1 downto 0);
    signal VN78_in1 : std_logic_vector(1 downto 0);
    signal VN78_in2 : std_logic_vector(1 downto 0);
    signal VN78_in3 : std_logic_vector(1 downto 0);
    signal VN78_in4 : std_logic_vector(1 downto 0);
    signal VN78_in5 : std_logic_vector(1 downto 0);
    signal VN79_in0 : std_logic_vector(1 downto 0);
    signal VN79_in1 : std_logic_vector(1 downto 0);
    signal VN79_in2 : std_logic_vector(1 downto 0);
    signal VN79_in3 : std_logic_vector(1 downto 0);
    signal VN79_in4 : std_logic_vector(1 downto 0);
    signal VN79_in5 : std_logic_vector(1 downto 0);
    signal VN80_in0 : std_logic_vector(1 downto 0);
    signal VN80_in1 : std_logic_vector(1 downto 0);
    signal VN80_in2 : std_logic_vector(1 downto 0);
    signal VN80_in3 : std_logic_vector(1 downto 0);
    signal VN80_in4 : std_logic_vector(1 downto 0);
    signal VN80_in5 : std_logic_vector(1 downto 0);
    signal VN81_in0 : std_logic_vector(1 downto 0);
    signal VN81_in1 : std_logic_vector(1 downto 0);
    signal VN81_in2 : std_logic_vector(1 downto 0);
    signal VN81_in3 : std_logic_vector(1 downto 0);
    signal VN81_in4 : std_logic_vector(1 downto 0);
    signal VN81_in5 : std_logic_vector(1 downto 0);
    signal VN82_in0 : std_logic_vector(1 downto 0);
    signal VN82_in1 : std_logic_vector(1 downto 0);
    signal VN82_in2 : std_logic_vector(1 downto 0);
    signal VN82_in3 : std_logic_vector(1 downto 0);
    signal VN82_in4 : std_logic_vector(1 downto 0);
    signal VN82_in5 : std_logic_vector(1 downto 0);
    signal VN83_in0 : std_logic_vector(1 downto 0);
    signal VN83_in1 : std_logic_vector(1 downto 0);
    signal VN83_in2 : std_logic_vector(1 downto 0);
    signal VN83_in3 : std_logic_vector(1 downto 0);
    signal VN83_in4 : std_logic_vector(1 downto 0);
    signal VN83_in5 : std_logic_vector(1 downto 0);
    signal VN84_in0 : std_logic_vector(1 downto 0);
    signal VN84_in1 : std_logic_vector(1 downto 0);
    signal VN84_in2 : std_logic_vector(1 downto 0);
    signal VN84_in3 : std_logic_vector(1 downto 0);
    signal VN84_in4 : std_logic_vector(1 downto 0);
    signal VN84_in5 : std_logic_vector(1 downto 0);
    signal VN85_in0 : std_logic_vector(1 downto 0);
    signal VN85_in1 : std_logic_vector(1 downto 0);
    signal VN85_in2 : std_logic_vector(1 downto 0);
    signal VN85_in3 : std_logic_vector(1 downto 0);
    signal VN85_in4 : std_logic_vector(1 downto 0);
    signal VN85_in5 : std_logic_vector(1 downto 0);
    signal VN86_in0 : std_logic_vector(1 downto 0);
    signal VN86_in1 : std_logic_vector(1 downto 0);
    signal VN86_in2 : std_logic_vector(1 downto 0);
    signal VN86_in3 : std_logic_vector(1 downto 0);
    signal VN86_in4 : std_logic_vector(1 downto 0);
    signal VN86_in5 : std_logic_vector(1 downto 0);
    signal VN87_in0 : std_logic_vector(1 downto 0);
    signal VN87_in1 : std_logic_vector(1 downto 0);
    signal VN87_in2 : std_logic_vector(1 downto 0);
    signal VN87_in3 : std_logic_vector(1 downto 0);
    signal VN87_in4 : std_logic_vector(1 downto 0);
    signal VN87_in5 : std_logic_vector(1 downto 0);
    signal VN88_in0 : std_logic_vector(1 downto 0);
    signal VN88_in1 : std_logic_vector(1 downto 0);
    signal VN88_in2 : std_logic_vector(1 downto 0);
    signal VN88_in3 : std_logic_vector(1 downto 0);
    signal VN88_in4 : std_logic_vector(1 downto 0);
    signal VN88_in5 : std_logic_vector(1 downto 0);
    signal VN89_in0 : std_logic_vector(1 downto 0);
    signal VN89_in1 : std_logic_vector(1 downto 0);
    signal VN89_in2 : std_logic_vector(1 downto 0);
    signal VN89_in3 : std_logic_vector(1 downto 0);
    signal VN89_in4 : std_logic_vector(1 downto 0);
    signal VN89_in5 : std_logic_vector(1 downto 0);
    signal VN90_in0 : std_logic_vector(1 downto 0);
    signal VN90_in1 : std_logic_vector(1 downto 0);
    signal VN90_in2 : std_logic_vector(1 downto 0);
    signal VN90_in3 : std_logic_vector(1 downto 0);
    signal VN90_in4 : std_logic_vector(1 downto 0);
    signal VN90_in5 : std_logic_vector(1 downto 0);
    signal VN91_in0 : std_logic_vector(1 downto 0);
    signal VN91_in1 : std_logic_vector(1 downto 0);
    signal VN91_in2 : std_logic_vector(1 downto 0);
    signal VN91_in3 : std_logic_vector(1 downto 0);
    signal VN91_in4 : std_logic_vector(1 downto 0);
    signal VN91_in5 : std_logic_vector(1 downto 0);
    signal VN92_in0 : std_logic_vector(1 downto 0);
    signal VN92_in1 : std_logic_vector(1 downto 0);
    signal VN92_in2 : std_logic_vector(1 downto 0);
    signal VN92_in3 : std_logic_vector(1 downto 0);
    signal VN92_in4 : std_logic_vector(1 downto 0);
    signal VN92_in5 : std_logic_vector(1 downto 0);
    signal VN93_in0 : std_logic_vector(1 downto 0);
    signal VN93_in1 : std_logic_vector(1 downto 0);
    signal VN93_in2 : std_logic_vector(1 downto 0);
    signal VN93_in3 : std_logic_vector(1 downto 0);
    signal VN93_in4 : std_logic_vector(1 downto 0);
    signal VN93_in5 : std_logic_vector(1 downto 0);
    signal VN94_in0 : std_logic_vector(1 downto 0);
    signal VN94_in1 : std_logic_vector(1 downto 0);
    signal VN94_in2 : std_logic_vector(1 downto 0);
    signal VN94_in3 : std_logic_vector(1 downto 0);
    signal VN94_in4 : std_logic_vector(1 downto 0);
    signal VN94_in5 : std_logic_vector(1 downto 0);
    signal VN95_in0 : std_logic_vector(1 downto 0);
    signal VN95_in1 : std_logic_vector(1 downto 0);
    signal VN95_in2 : std_logic_vector(1 downto 0);
    signal VN95_in3 : std_logic_vector(1 downto 0);
    signal VN95_in4 : std_logic_vector(1 downto 0);
    signal VN95_in5 : std_logic_vector(1 downto 0);
    signal VN96_in0 : std_logic_vector(1 downto 0);
    signal VN96_in1 : std_logic_vector(1 downto 0);
    signal VN96_in2 : std_logic_vector(1 downto 0);
    signal VN96_in3 : std_logic_vector(1 downto 0);
    signal VN96_in4 : std_logic_vector(1 downto 0);
    signal VN96_in5 : std_logic_vector(1 downto 0);
    signal VN97_in0 : std_logic_vector(1 downto 0);
    signal VN97_in1 : std_logic_vector(1 downto 0);
    signal VN97_in2 : std_logic_vector(1 downto 0);
    signal VN97_in3 : std_logic_vector(1 downto 0);
    signal VN97_in4 : std_logic_vector(1 downto 0);
    signal VN97_in5 : std_logic_vector(1 downto 0);
    signal VN98_in0 : std_logic_vector(1 downto 0);
    signal VN98_in1 : std_logic_vector(1 downto 0);
    signal VN98_in2 : std_logic_vector(1 downto 0);
    signal VN98_in3 : std_logic_vector(1 downto 0);
    signal VN98_in4 : std_logic_vector(1 downto 0);
    signal VN98_in5 : std_logic_vector(1 downto 0);
    signal VN99_in0 : std_logic_vector(1 downto 0);
    signal VN99_in1 : std_logic_vector(1 downto 0);
    signal VN99_in2 : std_logic_vector(1 downto 0);
    signal VN99_in3 : std_logic_vector(1 downto 0);
    signal VN99_in4 : std_logic_vector(1 downto 0);
    signal VN99_in5 : std_logic_vector(1 downto 0);
    signal VN100_in0 : std_logic_vector(1 downto 0);
    signal VN100_in1 : std_logic_vector(1 downto 0);
    signal VN100_in2 : std_logic_vector(1 downto 0);
    signal VN100_in3 : std_logic_vector(1 downto 0);
    signal VN100_in4 : std_logic_vector(1 downto 0);
    signal VN100_in5 : std_logic_vector(1 downto 0);
    signal VN101_in0 : std_logic_vector(1 downto 0);
    signal VN101_in1 : std_logic_vector(1 downto 0);
    signal VN101_in2 : std_logic_vector(1 downto 0);
    signal VN101_in3 : std_logic_vector(1 downto 0);
    signal VN101_in4 : std_logic_vector(1 downto 0);
    signal VN101_in5 : std_logic_vector(1 downto 0);
    signal VN102_in0 : std_logic_vector(1 downto 0);
    signal VN102_in1 : std_logic_vector(1 downto 0);
    signal VN102_in2 : std_logic_vector(1 downto 0);
    signal VN102_in3 : std_logic_vector(1 downto 0);
    signal VN102_in4 : std_logic_vector(1 downto 0);
    signal VN102_in5 : std_logic_vector(1 downto 0);
    signal VN103_in0 : std_logic_vector(1 downto 0);
    signal VN103_in1 : std_logic_vector(1 downto 0);
    signal VN103_in2 : std_logic_vector(1 downto 0);
    signal VN103_in3 : std_logic_vector(1 downto 0);
    signal VN103_in4 : std_logic_vector(1 downto 0);
    signal VN103_in5 : std_logic_vector(1 downto 0);
    signal VN104_in0 : std_logic_vector(1 downto 0);
    signal VN104_in1 : std_logic_vector(1 downto 0);
    signal VN104_in2 : std_logic_vector(1 downto 0);
    signal VN104_in3 : std_logic_vector(1 downto 0);
    signal VN104_in4 : std_logic_vector(1 downto 0);
    signal VN104_in5 : std_logic_vector(1 downto 0);
    signal VN105_in0 : std_logic_vector(1 downto 0);
    signal VN105_in1 : std_logic_vector(1 downto 0);
    signal VN105_in2 : std_logic_vector(1 downto 0);
    signal VN105_in3 : std_logic_vector(1 downto 0);
    signal VN105_in4 : std_logic_vector(1 downto 0);
    signal VN105_in5 : std_logic_vector(1 downto 0);
    signal VN106_in0 : std_logic_vector(1 downto 0);
    signal VN106_in1 : std_logic_vector(1 downto 0);
    signal VN106_in2 : std_logic_vector(1 downto 0);
    signal VN106_in3 : std_logic_vector(1 downto 0);
    signal VN106_in4 : std_logic_vector(1 downto 0);
    signal VN106_in5 : std_logic_vector(1 downto 0);
    signal VN107_in0 : std_logic_vector(1 downto 0);
    signal VN107_in1 : std_logic_vector(1 downto 0);
    signal VN107_in2 : std_logic_vector(1 downto 0);
    signal VN107_in3 : std_logic_vector(1 downto 0);
    signal VN107_in4 : std_logic_vector(1 downto 0);
    signal VN107_in5 : std_logic_vector(1 downto 0);
    signal VN108_in0 : std_logic_vector(1 downto 0);
    signal VN108_in1 : std_logic_vector(1 downto 0);
    signal VN108_in2 : std_logic_vector(1 downto 0);
    signal VN108_in3 : std_logic_vector(1 downto 0);
    signal VN108_in4 : std_logic_vector(1 downto 0);
    signal VN108_in5 : std_logic_vector(1 downto 0);
    signal VN109_in0 : std_logic_vector(1 downto 0);
    signal VN109_in1 : std_logic_vector(1 downto 0);
    signal VN109_in2 : std_logic_vector(1 downto 0);
    signal VN109_in3 : std_logic_vector(1 downto 0);
    signal VN109_in4 : std_logic_vector(1 downto 0);
    signal VN109_in5 : std_logic_vector(1 downto 0);
    signal VN110_in0 : std_logic_vector(1 downto 0);
    signal VN110_in1 : std_logic_vector(1 downto 0);
    signal VN110_in2 : std_logic_vector(1 downto 0);
    signal VN110_in3 : std_logic_vector(1 downto 0);
    signal VN110_in4 : std_logic_vector(1 downto 0);
    signal VN110_in5 : std_logic_vector(1 downto 0);
    signal VN111_in0 : std_logic_vector(1 downto 0);
    signal VN111_in1 : std_logic_vector(1 downto 0);
    signal VN111_in2 : std_logic_vector(1 downto 0);
    signal VN111_in3 : std_logic_vector(1 downto 0);
    signal VN111_in4 : std_logic_vector(1 downto 0);
    signal VN111_in5 : std_logic_vector(1 downto 0);
    signal VN112_in0 : std_logic_vector(1 downto 0);
    signal VN112_in1 : std_logic_vector(1 downto 0);
    signal VN112_in2 : std_logic_vector(1 downto 0);
    signal VN112_in3 : std_logic_vector(1 downto 0);
    signal VN112_in4 : std_logic_vector(1 downto 0);
    signal VN112_in5 : std_logic_vector(1 downto 0);
    signal VN113_in0 : std_logic_vector(1 downto 0);
    signal VN113_in1 : std_logic_vector(1 downto 0);
    signal VN113_in2 : std_logic_vector(1 downto 0);
    signal VN113_in3 : std_logic_vector(1 downto 0);
    signal VN113_in4 : std_logic_vector(1 downto 0);
    signal VN113_in5 : std_logic_vector(1 downto 0);
    signal VN114_in0 : std_logic_vector(1 downto 0);
    signal VN114_in1 : std_logic_vector(1 downto 0);
    signal VN114_in2 : std_logic_vector(1 downto 0);
    signal VN114_in3 : std_logic_vector(1 downto 0);
    signal VN114_in4 : std_logic_vector(1 downto 0);
    signal VN114_in5 : std_logic_vector(1 downto 0);
    signal VN115_in0 : std_logic_vector(1 downto 0);
    signal VN115_in1 : std_logic_vector(1 downto 0);
    signal VN115_in2 : std_logic_vector(1 downto 0);
    signal VN115_in3 : std_logic_vector(1 downto 0);
    signal VN115_in4 : std_logic_vector(1 downto 0);
    signal VN115_in5 : std_logic_vector(1 downto 0);
    signal VN116_in0 : std_logic_vector(1 downto 0);
    signal VN116_in1 : std_logic_vector(1 downto 0);
    signal VN116_in2 : std_logic_vector(1 downto 0);
    signal VN116_in3 : std_logic_vector(1 downto 0);
    signal VN116_in4 : std_logic_vector(1 downto 0);
    signal VN116_in5 : std_logic_vector(1 downto 0);
    signal VN117_in0 : std_logic_vector(1 downto 0);
    signal VN117_in1 : std_logic_vector(1 downto 0);
    signal VN117_in2 : std_logic_vector(1 downto 0);
    signal VN117_in3 : std_logic_vector(1 downto 0);
    signal VN117_in4 : std_logic_vector(1 downto 0);
    signal VN117_in5 : std_logic_vector(1 downto 0);
    signal VN118_in0 : std_logic_vector(1 downto 0);
    signal VN118_in1 : std_logic_vector(1 downto 0);
    signal VN118_in2 : std_logic_vector(1 downto 0);
    signal VN118_in3 : std_logic_vector(1 downto 0);
    signal VN118_in4 : std_logic_vector(1 downto 0);
    signal VN118_in5 : std_logic_vector(1 downto 0);
    signal VN119_in0 : std_logic_vector(1 downto 0);
    signal VN119_in1 : std_logic_vector(1 downto 0);
    signal VN119_in2 : std_logic_vector(1 downto 0);
    signal VN119_in3 : std_logic_vector(1 downto 0);
    signal VN119_in4 : std_logic_vector(1 downto 0);
    signal VN119_in5 : std_logic_vector(1 downto 0);
    signal VN120_in0 : std_logic_vector(1 downto 0);
    signal VN120_in1 : std_logic_vector(1 downto 0);
    signal VN120_in2 : std_logic_vector(1 downto 0);
    signal VN120_in3 : std_logic_vector(1 downto 0);
    signal VN120_in4 : std_logic_vector(1 downto 0);
    signal VN120_in5 : std_logic_vector(1 downto 0);
    signal VN121_in0 : std_logic_vector(1 downto 0);
    signal VN121_in1 : std_logic_vector(1 downto 0);
    signal VN121_in2 : std_logic_vector(1 downto 0);
    signal VN121_in3 : std_logic_vector(1 downto 0);
    signal VN121_in4 : std_logic_vector(1 downto 0);
    signal VN121_in5 : std_logic_vector(1 downto 0);
    signal VN122_in0 : std_logic_vector(1 downto 0);
    signal VN122_in1 : std_logic_vector(1 downto 0);
    signal VN122_in2 : std_logic_vector(1 downto 0);
    signal VN122_in3 : std_logic_vector(1 downto 0);
    signal VN122_in4 : std_logic_vector(1 downto 0);
    signal VN122_in5 : std_logic_vector(1 downto 0);
    signal VN123_in0 : std_logic_vector(1 downto 0);
    signal VN123_in1 : std_logic_vector(1 downto 0);
    signal VN123_in2 : std_logic_vector(1 downto 0);
    signal VN123_in3 : std_logic_vector(1 downto 0);
    signal VN123_in4 : std_logic_vector(1 downto 0);
    signal VN123_in5 : std_logic_vector(1 downto 0);
    signal VN124_in0 : std_logic_vector(1 downto 0);
    signal VN124_in1 : std_logic_vector(1 downto 0);
    signal VN124_in2 : std_logic_vector(1 downto 0);
    signal VN124_in3 : std_logic_vector(1 downto 0);
    signal VN124_in4 : std_logic_vector(1 downto 0);
    signal VN124_in5 : std_logic_vector(1 downto 0);
    signal VN125_in0 : std_logic_vector(1 downto 0);
    signal VN125_in1 : std_logic_vector(1 downto 0);
    signal VN125_in2 : std_logic_vector(1 downto 0);
    signal VN125_in3 : std_logic_vector(1 downto 0);
    signal VN125_in4 : std_logic_vector(1 downto 0);
    signal VN125_in5 : std_logic_vector(1 downto 0);
    signal VN126_in0 : std_logic_vector(1 downto 0);
    signal VN126_in1 : std_logic_vector(1 downto 0);
    signal VN126_in2 : std_logic_vector(1 downto 0);
    signal VN126_in3 : std_logic_vector(1 downto 0);
    signal VN126_in4 : std_logic_vector(1 downto 0);
    signal VN126_in5 : std_logic_vector(1 downto 0);
    signal VN127_in0 : std_logic_vector(1 downto 0);
    signal VN127_in1 : std_logic_vector(1 downto 0);
    signal VN127_in2 : std_logic_vector(1 downto 0);
    signal VN127_in3 : std_logic_vector(1 downto 0);
    signal VN127_in4 : std_logic_vector(1 downto 0);
    signal VN127_in5 : std_logic_vector(1 downto 0);
    signal VN128_in0 : std_logic_vector(1 downto 0);
    signal VN128_in1 : std_logic_vector(1 downto 0);
    signal VN128_in2 : std_logic_vector(1 downto 0);
    signal VN128_in3 : std_logic_vector(1 downto 0);
    signal VN128_in4 : std_logic_vector(1 downto 0);
    signal VN128_in5 : std_logic_vector(1 downto 0);
    signal VN129_in0 : std_logic_vector(1 downto 0);
    signal VN129_in1 : std_logic_vector(1 downto 0);
    signal VN129_in2 : std_logic_vector(1 downto 0);
    signal VN129_in3 : std_logic_vector(1 downto 0);
    signal VN129_in4 : std_logic_vector(1 downto 0);
    signal VN129_in5 : std_logic_vector(1 downto 0);
    signal VN130_in0 : std_logic_vector(1 downto 0);
    signal VN130_in1 : std_logic_vector(1 downto 0);
    signal VN130_in2 : std_logic_vector(1 downto 0);
    signal VN130_in3 : std_logic_vector(1 downto 0);
    signal VN130_in4 : std_logic_vector(1 downto 0);
    signal VN130_in5 : std_logic_vector(1 downto 0);
    signal VN131_in0 : std_logic_vector(1 downto 0);
    signal VN131_in1 : std_logic_vector(1 downto 0);
    signal VN131_in2 : std_logic_vector(1 downto 0);
    signal VN131_in3 : std_logic_vector(1 downto 0);
    signal VN131_in4 : std_logic_vector(1 downto 0);
    signal VN131_in5 : std_logic_vector(1 downto 0);
    signal VN132_in0 : std_logic_vector(1 downto 0);
    signal VN132_in1 : std_logic_vector(1 downto 0);
    signal VN132_in2 : std_logic_vector(1 downto 0);
    signal VN132_in3 : std_logic_vector(1 downto 0);
    signal VN132_in4 : std_logic_vector(1 downto 0);
    signal VN132_in5 : std_logic_vector(1 downto 0);
    signal VN133_in0 : std_logic_vector(1 downto 0);
    signal VN133_in1 : std_logic_vector(1 downto 0);
    signal VN133_in2 : std_logic_vector(1 downto 0);
    signal VN133_in3 : std_logic_vector(1 downto 0);
    signal VN133_in4 : std_logic_vector(1 downto 0);
    signal VN133_in5 : std_logic_vector(1 downto 0);
    signal VN134_in0 : std_logic_vector(1 downto 0);
    signal VN134_in1 : std_logic_vector(1 downto 0);
    signal VN134_in2 : std_logic_vector(1 downto 0);
    signal VN134_in3 : std_logic_vector(1 downto 0);
    signal VN134_in4 : std_logic_vector(1 downto 0);
    signal VN134_in5 : std_logic_vector(1 downto 0);
    signal VN135_in0 : std_logic_vector(1 downto 0);
    signal VN135_in1 : std_logic_vector(1 downto 0);
    signal VN135_in2 : std_logic_vector(1 downto 0);
    signal VN135_in3 : std_logic_vector(1 downto 0);
    signal VN135_in4 : std_logic_vector(1 downto 0);
    signal VN135_in5 : std_logic_vector(1 downto 0);
    signal VN136_in0 : std_logic_vector(1 downto 0);
    signal VN136_in1 : std_logic_vector(1 downto 0);
    signal VN136_in2 : std_logic_vector(1 downto 0);
    signal VN136_in3 : std_logic_vector(1 downto 0);
    signal VN136_in4 : std_logic_vector(1 downto 0);
    signal VN136_in5 : std_logic_vector(1 downto 0);
    signal VN137_in0 : std_logic_vector(1 downto 0);
    signal VN137_in1 : std_logic_vector(1 downto 0);
    signal VN137_in2 : std_logic_vector(1 downto 0);
    signal VN137_in3 : std_logic_vector(1 downto 0);
    signal VN137_in4 : std_logic_vector(1 downto 0);
    signal VN137_in5 : std_logic_vector(1 downto 0);
    signal VN138_in0 : std_logic_vector(1 downto 0);
    signal VN138_in1 : std_logic_vector(1 downto 0);
    signal VN138_in2 : std_logic_vector(1 downto 0);
    signal VN138_in3 : std_logic_vector(1 downto 0);
    signal VN138_in4 : std_logic_vector(1 downto 0);
    signal VN138_in5 : std_logic_vector(1 downto 0);
    signal VN139_in0 : std_logic_vector(1 downto 0);
    signal VN139_in1 : std_logic_vector(1 downto 0);
    signal VN139_in2 : std_logic_vector(1 downto 0);
    signal VN139_in3 : std_logic_vector(1 downto 0);
    signal VN139_in4 : std_logic_vector(1 downto 0);
    signal VN139_in5 : std_logic_vector(1 downto 0);
    signal VN140_in0 : std_logic_vector(1 downto 0);
    signal VN140_in1 : std_logic_vector(1 downto 0);
    signal VN140_in2 : std_logic_vector(1 downto 0);
    signal VN140_in3 : std_logic_vector(1 downto 0);
    signal VN140_in4 : std_logic_vector(1 downto 0);
    signal VN140_in5 : std_logic_vector(1 downto 0);
    signal VN141_in0 : std_logic_vector(1 downto 0);
    signal VN141_in1 : std_logic_vector(1 downto 0);
    signal VN141_in2 : std_logic_vector(1 downto 0);
    signal VN141_in3 : std_logic_vector(1 downto 0);
    signal VN141_in4 : std_logic_vector(1 downto 0);
    signal VN141_in5 : std_logic_vector(1 downto 0);
    signal VN142_in0 : std_logic_vector(1 downto 0);
    signal VN142_in1 : std_logic_vector(1 downto 0);
    signal VN142_in2 : std_logic_vector(1 downto 0);
    signal VN142_in3 : std_logic_vector(1 downto 0);
    signal VN142_in4 : std_logic_vector(1 downto 0);
    signal VN142_in5 : std_logic_vector(1 downto 0);
    signal VN143_in0 : std_logic_vector(1 downto 0);
    signal VN143_in1 : std_logic_vector(1 downto 0);
    signal VN143_in2 : std_logic_vector(1 downto 0);
    signal VN143_in3 : std_logic_vector(1 downto 0);
    signal VN143_in4 : std_logic_vector(1 downto 0);
    signal VN143_in5 : std_logic_vector(1 downto 0);
    signal VN144_in0 : std_logic_vector(1 downto 0);
    signal VN144_in1 : std_logic_vector(1 downto 0);
    signal VN144_in2 : std_logic_vector(1 downto 0);
    signal VN144_in3 : std_logic_vector(1 downto 0);
    signal VN144_in4 : std_logic_vector(1 downto 0);
    signal VN144_in5 : std_logic_vector(1 downto 0);
    signal VN145_in0 : std_logic_vector(1 downto 0);
    signal VN145_in1 : std_logic_vector(1 downto 0);
    signal VN145_in2 : std_logic_vector(1 downto 0);
    signal VN145_in3 : std_logic_vector(1 downto 0);
    signal VN145_in4 : std_logic_vector(1 downto 0);
    signal VN145_in5 : std_logic_vector(1 downto 0);
    signal VN146_in0 : std_logic_vector(1 downto 0);
    signal VN146_in1 : std_logic_vector(1 downto 0);
    signal VN146_in2 : std_logic_vector(1 downto 0);
    signal VN146_in3 : std_logic_vector(1 downto 0);
    signal VN146_in4 : std_logic_vector(1 downto 0);
    signal VN146_in5 : std_logic_vector(1 downto 0);
    signal VN147_in0 : std_logic_vector(1 downto 0);
    signal VN147_in1 : std_logic_vector(1 downto 0);
    signal VN147_in2 : std_logic_vector(1 downto 0);
    signal VN147_in3 : std_logic_vector(1 downto 0);
    signal VN147_in4 : std_logic_vector(1 downto 0);
    signal VN147_in5 : std_logic_vector(1 downto 0);
    signal VN148_in0 : std_logic_vector(1 downto 0);
    signal VN148_in1 : std_logic_vector(1 downto 0);
    signal VN148_in2 : std_logic_vector(1 downto 0);
    signal VN148_in3 : std_logic_vector(1 downto 0);
    signal VN148_in4 : std_logic_vector(1 downto 0);
    signal VN148_in5 : std_logic_vector(1 downto 0);
    signal VN149_in0 : std_logic_vector(1 downto 0);
    signal VN149_in1 : std_logic_vector(1 downto 0);
    signal VN149_in2 : std_logic_vector(1 downto 0);
    signal VN149_in3 : std_logic_vector(1 downto 0);
    signal VN149_in4 : std_logic_vector(1 downto 0);
    signal VN149_in5 : std_logic_vector(1 downto 0);
    signal VN150_in0 : std_logic_vector(1 downto 0);
    signal VN150_in1 : std_logic_vector(1 downto 0);
    signal VN150_in2 : std_logic_vector(1 downto 0);
    signal VN150_in3 : std_logic_vector(1 downto 0);
    signal VN150_in4 : std_logic_vector(1 downto 0);
    signal VN150_in5 : std_logic_vector(1 downto 0);
    signal VN151_in0 : std_logic_vector(1 downto 0);
    signal VN151_in1 : std_logic_vector(1 downto 0);
    signal VN151_in2 : std_logic_vector(1 downto 0);
    signal VN151_in3 : std_logic_vector(1 downto 0);
    signal VN151_in4 : std_logic_vector(1 downto 0);
    signal VN151_in5 : std_logic_vector(1 downto 0);
    signal VN152_in0 : std_logic_vector(1 downto 0);
    signal VN152_in1 : std_logic_vector(1 downto 0);
    signal VN152_in2 : std_logic_vector(1 downto 0);
    signal VN152_in3 : std_logic_vector(1 downto 0);
    signal VN152_in4 : std_logic_vector(1 downto 0);
    signal VN152_in5 : std_logic_vector(1 downto 0);
    signal VN153_in0 : std_logic_vector(1 downto 0);
    signal VN153_in1 : std_logic_vector(1 downto 0);
    signal VN153_in2 : std_logic_vector(1 downto 0);
    signal VN153_in3 : std_logic_vector(1 downto 0);
    signal VN153_in4 : std_logic_vector(1 downto 0);
    signal VN153_in5 : std_logic_vector(1 downto 0);
    signal VN154_in0 : std_logic_vector(1 downto 0);
    signal VN154_in1 : std_logic_vector(1 downto 0);
    signal VN154_in2 : std_logic_vector(1 downto 0);
    signal VN154_in3 : std_logic_vector(1 downto 0);
    signal VN154_in4 : std_logic_vector(1 downto 0);
    signal VN154_in5 : std_logic_vector(1 downto 0);
    signal VN155_in0 : std_logic_vector(1 downto 0);
    signal VN155_in1 : std_logic_vector(1 downto 0);
    signal VN155_in2 : std_logic_vector(1 downto 0);
    signal VN155_in3 : std_logic_vector(1 downto 0);
    signal VN155_in4 : std_logic_vector(1 downto 0);
    signal VN155_in5 : std_logic_vector(1 downto 0);
    signal VN156_in0 : std_logic_vector(1 downto 0);
    signal VN156_in1 : std_logic_vector(1 downto 0);
    signal VN156_in2 : std_logic_vector(1 downto 0);
    signal VN156_in3 : std_logic_vector(1 downto 0);
    signal VN156_in4 : std_logic_vector(1 downto 0);
    signal VN156_in5 : std_logic_vector(1 downto 0);
    signal VN157_in0 : std_logic_vector(1 downto 0);
    signal VN157_in1 : std_logic_vector(1 downto 0);
    signal VN157_in2 : std_logic_vector(1 downto 0);
    signal VN157_in3 : std_logic_vector(1 downto 0);
    signal VN157_in4 : std_logic_vector(1 downto 0);
    signal VN157_in5 : std_logic_vector(1 downto 0);
    signal VN158_in0 : std_logic_vector(1 downto 0);
    signal VN158_in1 : std_logic_vector(1 downto 0);
    signal VN158_in2 : std_logic_vector(1 downto 0);
    signal VN158_in3 : std_logic_vector(1 downto 0);
    signal VN158_in4 : std_logic_vector(1 downto 0);
    signal VN158_in5 : std_logic_vector(1 downto 0);
    signal VN159_in0 : std_logic_vector(1 downto 0);
    signal VN159_in1 : std_logic_vector(1 downto 0);
    signal VN159_in2 : std_logic_vector(1 downto 0);
    signal VN159_in3 : std_logic_vector(1 downto 0);
    signal VN159_in4 : std_logic_vector(1 downto 0);
    signal VN159_in5 : std_logic_vector(1 downto 0);
    signal VN160_in0 : std_logic_vector(1 downto 0);
    signal VN160_in1 : std_logic_vector(1 downto 0);
    signal VN160_in2 : std_logic_vector(1 downto 0);
    signal VN160_in3 : std_logic_vector(1 downto 0);
    signal VN160_in4 : std_logic_vector(1 downto 0);
    signal VN160_in5 : std_logic_vector(1 downto 0);
    signal VN161_in0 : std_logic_vector(1 downto 0);
    signal VN161_in1 : std_logic_vector(1 downto 0);
    signal VN161_in2 : std_logic_vector(1 downto 0);
    signal VN161_in3 : std_logic_vector(1 downto 0);
    signal VN161_in4 : std_logic_vector(1 downto 0);
    signal VN161_in5 : std_logic_vector(1 downto 0);
    signal VN162_in0 : std_logic_vector(1 downto 0);
    signal VN162_in1 : std_logic_vector(1 downto 0);
    signal VN162_in2 : std_logic_vector(1 downto 0);
    signal VN162_in3 : std_logic_vector(1 downto 0);
    signal VN162_in4 : std_logic_vector(1 downto 0);
    signal VN162_in5 : std_logic_vector(1 downto 0);
    signal VN163_in0 : std_logic_vector(1 downto 0);
    signal VN163_in1 : std_logic_vector(1 downto 0);
    signal VN163_in2 : std_logic_vector(1 downto 0);
    signal VN163_in3 : std_logic_vector(1 downto 0);
    signal VN163_in4 : std_logic_vector(1 downto 0);
    signal VN163_in5 : std_logic_vector(1 downto 0);
    signal VN164_in0 : std_logic_vector(1 downto 0);
    signal VN164_in1 : std_logic_vector(1 downto 0);
    signal VN164_in2 : std_logic_vector(1 downto 0);
    signal VN164_in3 : std_logic_vector(1 downto 0);
    signal VN164_in4 : std_logic_vector(1 downto 0);
    signal VN164_in5 : std_logic_vector(1 downto 0);
    signal VN165_in0 : std_logic_vector(1 downto 0);
    signal VN165_in1 : std_logic_vector(1 downto 0);
    signal VN165_in2 : std_logic_vector(1 downto 0);
    signal VN165_in3 : std_logic_vector(1 downto 0);
    signal VN165_in4 : std_logic_vector(1 downto 0);
    signal VN165_in5 : std_logic_vector(1 downto 0);
    signal VN166_in0 : std_logic_vector(1 downto 0);
    signal VN166_in1 : std_logic_vector(1 downto 0);
    signal VN166_in2 : std_logic_vector(1 downto 0);
    signal VN166_in3 : std_logic_vector(1 downto 0);
    signal VN166_in4 : std_logic_vector(1 downto 0);
    signal VN166_in5 : std_logic_vector(1 downto 0);
    signal VN167_in0 : std_logic_vector(1 downto 0);
    signal VN167_in1 : std_logic_vector(1 downto 0);
    signal VN167_in2 : std_logic_vector(1 downto 0);
    signal VN167_in3 : std_logic_vector(1 downto 0);
    signal VN167_in4 : std_logic_vector(1 downto 0);
    signal VN167_in5 : std_logic_vector(1 downto 0);
    signal VN168_in0 : std_logic_vector(1 downto 0);
    signal VN168_in1 : std_logic_vector(1 downto 0);
    signal VN168_in2 : std_logic_vector(1 downto 0);
    signal VN168_in3 : std_logic_vector(1 downto 0);
    signal VN168_in4 : std_logic_vector(1 downto 0);
    signal VN168_in5 : std_logic_vector(1 downto 0);
    signal VN169_in0 : std_logic_vector(1 downto 0);
    signal VN169_in1 : std_logic_vector(1 downto 0);
    signal VN169_in2 : std_logic_vector(1 downto 0);
    signal VN169_in3 : std_logic_vector(1 downto 0);
    signal VN169_in4 : std_logic_vector(1 downto 0);
    signal VN169_in5 : std_logic_vector(1 downto 0);
    signal VN170_in0 : std_logic_vector(1 downto 0);
    signal VN170_in1 : std_logic_vector(1 downto 0);
    signal VN170_in2 : std_logic_vector(1 downto 0);
    signal VN170_in3 : std_logic_vector(1 downto 0);
    signal VN170_in4 : std_logic_vector(1 downto 0);
    signal VN170_in5 : std_logic_vector(1 downto 0);
    signal VN171_in0 : std_logic_vector(1 downto 0);
    signal VN171_in1 : std_logic_vector(1 downto 0);
    signal VN171_in2 : std_logic_vector(1 downto 0);
    signal VN171_in3 : std_logic_vector(1 downto 0);
    signal VN171_in4 : std_logic_vector(1 downto 0);
    signal VN171_in5 : std_logic_vector(1 downto 0);
    signal VN172_in0 : std_logic_vector(1 downto 0);
    signal VN172_in1 : std_logic_vector(1 downto 0);
    signal VN172_in2 : std_logic_vector(1 downto 0);
    signal VN172_in3 : std_logic_vector(1 downto 0);
    signal VN172_in4 : std_logic_vector(1 downto 0);
    signal VN172_in5 : std_logic_vector(1 downto 0);
    signal VN173_in0 : std_logic_vector(1 downto 0);
    signal VN173_in1 : std_logic_vector(1 downto 0);
    signal VN173_in2 : std_logic_vector(1 downto 0);
    signal VN173_in3 : std_logic_vector(1 downto 0);
    signal VN173_in4 : std_logic_vector(1 downto 0);
    signal VN173_in5 : std_logic_vector(1 downto 0);
    signal VN174_in0 : std_logic_vector(1 downto 0);
    signal VN174_in1 : std_logic_vector(1 downto 0);
    signal VN174_in2 : std_logic_vector(1 downto 0);
    signal VN174_in3 : std_logic_vector(1 downto 0);
    signal VN174_in4 : std_logic_vector(1 downto 0);
    signal VN174_in5 : std_logic_vector(1 downto 0);
    signal VN175_in0 : std_logic_vector(1 downto 0);
    signal VN175_in1 : std_logic_vector(1 downto 0);
    signal VN175_in2 : std_logic_vector(1 downto 0);
    signal VN175_in3 : std_logic_vector(1 downto 0);
    signal VN175_in4 : std_logic_vector(1 downto 0);
    signal VN175_in5 : std_logic_vector(1 downto 0);
    signal VN176_in0 : std_logic_vector(1 downto 0);
    signal VN176_in1 : std_logic_vector(1 downto 0);
    signal VN176_in2 : std_logic_vector(1 downto 0);
    signal VN176_in3 : std_logic_vector(1 downto 0);
    signal VN176_in4 : std_logic_vector(1 downto 0);
    signal VN176_in5 : std_logic_vector(1 downto 0);
    signal VN177_in0 : std_logic_vector(1 downto 0);
    signal VN177_in1 : std_logic_vector(1 downto 0);
    signal VN177_in2 : std_logic_vector(1 downto 0);
    signal VN177_in3 : std_logic_vector(1 downto 0);
    signal VN177_in4 : std_logic_vector(1 downto 0);
    signal VN177_in5 : std_logic_vector(1 downto 0);
    signal VN178_in0 : std_logic_vector(1 downto 0);
    signal VN178_in1 : std_logic_vector(1 downto 0);
    signal VN178_in2 : std_logic_vector(1 downto 0);
    signal VN178_in3 : std_logic_vector(1 downto 0);
    signal VN178_in4 : std_logic_vector(1 downto 0);
    signal VN178_in5 : std_logic_vector(1 downto 0);
    signal VN179_in0 : std_logic_vector(1 downto 0);
    signal VN179_in1 : std_logic_vector(1 downto 0);
    signal VN179_in2 : std_logic_vector(1 downto 0);
    signal VN179_in3 : std_logic_vector(1 downto 0);
    signal VN179_in4 : std_logic_vector(1 downto 0);
    signal VN179_in5 : std_logic_vector(1 downto 0);
    signal VN180_in0 : std_logic_vector(1 downto 0);
    signal VN180_in1 : std_logic_vector(1 downto 0);
    signal VN180_in2 : std_logic_vector(1 downto 0);
    signal VN180_in3 : std_logic_vector(1 downto 0);
    signal VN180_in4 : std_logic_vector(1 downto 0);
    signal VN180_in5 : std_logic_vector(1 downto 0);
    signal VN181_in0 : std_logic_vector(1 downto 0);
    signal VN181_in1 : std_logic_vector(1 downto 0);
    signal VN181_in2 : std_logic_vector(1 downto 0);
    signal VN181_in3 : std_logic_vector(1 downto 0);
    signal VN181_in4 : std_logic_vector(1 downto 0);
    signal VN181_in5 : std_logic_vector(1 downto 0);
    signal VN182_in0 : std_logic_vector(1 downto 0);
    signal VN182_in1 : std_logic_vector(1 downto 0);
    signal VN182_in2 : std_logic_vector(1 downto 0);
    signal VN182_in3 : std_logic_vector(1 downto 0);
    signal VN182_in4 : std_logic_vector(1 downto 0);
    signal VN182_in5 : std_logic_vector(1 downto 0);
    signal VN183_in0 : std_logic_vector(1 downto 0);
    signal VN183_in1 : std_logic_vector(1 downto 0);
    signal VN183_in2 : std_logic_vector(1 downto 0);
    signal VN183_in3 : std_logic_vector(1 downto 0);
    signal VN183_in4 : std_logic_vector(1 downto 0);
    signal VN183_in5 : std_logic_vector(1 downto 0);
    signal VN184_in0 : std_logic_vector(1 downto 0);
    signal VN184_in1 : std_logic_vector(1 downto 0);
    signal VN184_in2 : std_logic_vector(1 downto 0);
    signal VN184_in3 : std_logic_vector(1 downto 0);
    signal VN184_in4 : std_logic_vector(1 downto 0);
    signal VN184_in5 : std_logic_vector(1 downto 0);
    signal VN185_in0 : std_logic_vector(1 downto 0);
    signal VN185_in1 : std_logic_vector(1 downto 0);
    signal VN185_in2 : std_logic_vector(1 downto 0);
    signal VN185_in3 : std_logic_vector(1 downto 0);
    signal VN185_in4 : std_logic_vector(1 downto 0);
    signal VN185_in5 : std_logic_vector(1 downto 0);
    signal VN186_in0 : std_logic_vector(1 downto 0);
    signal VN186_in1 : std_logic_vector(1 downto 0);
    signal VN186_in2 : std_logic_vector(1 downto 0);
    signal VN186_in3 : std_logic_vector(1 downto 0);
    signal VN186_in4 : std_logic_vector(1 downto 0);
    signal VN186_in5 : std_logic_vector(1 downto 0);
    signal VN187_in0 : std_logic_vector(1 downto 0);
    signal VN187_in1 : std_logic_vector(1 downto 0);
    signal VN187_in2 : std_logic_vector(1 downto 0);
    signal VN187_in3 : std_logic_vector(1 downto 0);
    signal VN187_in4 : std_logic_vector(1 downto 0);
    signal VN187_in5 : std_logic_vector(1 downto 0);
    signal VN188_in0 : std_logic_vector(1 downto 0);
    signal VN188_in1 : std_logic_vector(1 downto 0);
    signal VN188_in2 : std_logic_vector(1 downto 0);
    signal VN188_in3 : std_logic_vector(1 downto 0);
    signal VN188_in4 : std_logic_vector(1 downto 0);
    signal VN188_in5 : std_logic_vector(1 downto 0);
    signal VN189_in0 : std_logic_vector(1 downto 0);
    signal VN189_in1 : std_logic_vector(1 downto 0);
    signal VN189_in2 : std_logic_vector(1 downto 0);
    signal VN189_in3 : std_logic_vector(1 downto 0);
    signal VN189_in4 : std_logic_vector(1 downto 0);
    signal VN189_in5 : std_logic_vector(1 downto 0);
    signal VN190_in0 : std_logic_vector(1 downto 0);
    signal VN190_in1 : std_logic_vector(1 downto 0);
    signal VN190_in2 : std_logic_vector(1 downto 0);
    signal VN190_in3 : std_logic_vector(1 downto 0);
    signal VN190_in4 : std_logic_vector(1 downto 0);
    signal VN190_in5 : std_logic_vector(1 downto 0);
    signal VN191_in0 : std_logic_vector(1 downto 0);
    signal VN191_in1 : std_logic_vector(1 downto 0);
    signal VN191_in2 : std_logic_vector(1 downto 0);
    signal VN191_in3 : std_logic_vector(1 downto 0);
    signal VN191_in4 : std_logic_vector(1 downto 0);
    signal VN191_in5 : std_logic_vector(1 downto 0);
    signal VN192_in0 : std_logic_vector(1 downto 0);
    signal VN192_in1 : std_logic_vector(1 downto 0);
    signal VN192_in2 : std_logic_vector(1 downto 0);
    signal VN192_in3 : std_logic_vector(1 downto 0);
    signal VN192_in4 : std_logic_vector(1 downto 0);
    signal VN192_in5 : std_logic_vector(1 downto 0);
    signal VN193_in0 : std_logic_vector(1 downto 0);
    signal VN193_in1 : std_logic_vector(1 downto 0);
    signal VN193_in2 : std_logic_vector(1 downto 0);
    signal VN193_in3 : std_logic_vector(1 downto 0);
    signal VN193_in4 : std_logic_vector(1 downto 0);
    signal VN193_in5 : std_logic_vector(1 downto 0);
    signal VN194_in0 : std_logic_vector(1 downto 0);
    signal VN194_in1 : std_logic_vector(1 downto 0);
    signal VN194_in2 : std_logic_vector(1 downto 0);
    signal VN194_in3 : std_logic_vector(1 downto 0);
    signal VN194_in4 : std_logic_vector(1 downto 0);
    signal VN194_in5 : std_logic_vector(1 downto 0);
    signal VN195_in0 : std_logic_vector(1 downto 0);
    signal VN195_in1 : std_logic_vector(1 downto 0);
    signal VN195_in2 : std_logic_vector(1 downto 0);
    signal VN195_in3 : std_logic_vector(1 downto 0);
    signal VN195_in4 : std_logic_vector(1 downto 0);
    signal VN195_in5 : std_logic_vector(1 downto 0);
    signal VN196_in0 : std_logic_vector(1 downto 0);
    signal VN196_in1 : std_logic_vector(1 downto 0);
    signal VN196_in2 : std_logic_vector(1 downto 0);
    signal VN196_in3 : std_logic_vector(1 downto 0);
    signal VN196_in4 : std_logic_vector(1 downto 0);
    signal VN196_in5 : std_logic_vector(1 downto 0);
    signal VN197_in0 : std_logic_vector(1 downto 0);
    signal VN197_in1 : std_logic_vector(1 downto 0);
    signal VN197_in2 : std_logic_vector(1 downto 0);
    signal VN197_in3 : std_logic_vector(1 downto 0);
    signal VN197_in4 : std_logic_vector(1 downto 0);
    signal VN197_in5 : std_logic_vector(1 downto 0);
    signal VN198_in0 : std_logic_vector(1 downto 0);
    signal VN198_in1 : std_logic_vector(1 downto 0);
    signal VN198_in2 : std_logic_vector(1 downto 0);
    signal VN198_in3 : std_logic_vector(1 downto 0);
    signal VN198_in4 : std_logic_vector(1 downto 0);
    signal VN198_in5 : std_logic_vector(1 downto 0);
    signal VN199_in0 : std_logic_vector(1 downto 0);
    signal VN199_in1 : std_logic_vector(1 downto 0);
    signal VN199_in2 : std_logic_vector(1 downto 0);
    signal VN199_in3 : std_logic_vector(1 downto 0);
    signal VN199_in4 : std_logic_vector(1 downto 0);
    signal VN199_in5 : std_logic_vector(1 downto 0);
    signal VN200_in0 : std_logic_vector(1 downto 0);
    signal VN200_in1 : std_logic_vector(1 downto 0);
    signal VN200_in2 : std_logic_vector(1 downto 0);
    signal VN200_in3 : std_logic_vector(1 downto 0);
    signal VN200_in4 : std_logic_vector(1 downto 0);
    signal VN200_in5 : std_logic_vector(1 downto 0);
    signal VN201_in0 : std_logic_vector(1 downto 0);
    signal VN201_in1 : std_logic_vector(1 downto 0);
    signal VN201_in2 : std_logic_vector(1 downto 0);
    signal VN201_in3 : std_logic_vector(1 downto 0);
    signal VN201_in4 : std_logic_vector(1 downto 0);
    signal VN201_in5 : std_logic_vector(1 downto 0);
    signal VN202_in0 : std_logic_vector(1 downto 0);
    signal VN202_in1 : std_logic_vector(1 downto 0);
    signal VN202_in2 : std_logic_vector(1 downto 0);
    signal VN202_in3 : std_logic_vector(1 downto 0);
    signal VN202_in4 : std_logic_vector(1 downto 0);
    signal VN202_in5 : std_logic_vector(1 downto 0);
    signal VN203_in0 : std_logic_vector(1 downto 0);
    signal VN203_in1 : std_logic_vector(1 downto 0);
    signal VN203_in2 : std_logic_vector(1 downto 0);
    signal VN203_in3 : std_logic_vector(1 downto 0);
    signal VN203_in4 : std_logic_vector(1 downto 0);
    signal VN203_in5 : std_logic_vector(1 downto 0);
    signal VN204_in0 : std_logic_vector(1 downto 0);
    signal VN204_in1 : std_logic_vector(1 downto 0);
    signal VN204_in2 : std_logic_vector(1 downto 0);
    signal VN204_in3 : std_logic_vector(1 downto 0);
    signal VN204_in4 : std_logic_vector(1 downto 0);
    signal VN204_in5 : std_logic_vector(1 downto 0);
    signal VN205_in0 : std_logic_vector(1 downto 0);
    signal VN205_in1 : std_logic_vector(1 downto 0);
    signal VN205_in2 : std_logic_vector(1 downto 0);
    signal VN205_in3 : std_logic_vector(1 downto 0);
    signal VN205_in4 : std_logic_vector(1 downto 0);
    signal VN205_in5 : std_logic_vector(1 downto 0);
    signal VN206_in0 : std_logic_vector(1 downto 0);
    signal VN206_in1 : std_logic_vector(1 downto 0);
    signal VN206_in2 : std_logic_vector(1 downto 0);
    signal VN206_in3 : std_logic_vector(1 downto 0);
    signal VN206_in4 : std_logic_vector(1 downto 0);
    signal VN206_in5 : std_logic_vector(1 downto 0);
    signal VN207_in0 : std_logic_vector(1 downto 0);
    signal VN207_in1 : std_logic_vector(1 downto 0);
    signal VN207_in2 : std_logic_vector(1 downto 0);
    signal VN207_in3 : std_logic_vector(1 downto 0);
    signal VN207_in4 : std_logic_vector(1 downto 0);
    signal VN207_in5 : std_logic_vector(1 downto 0);
    signal VN208_in0 : std_logic_vector(1 downto 0);
    signal VN208_in1 : std_logic_vector(1 downto 0);
    signal VN208_in2 : std_logic_vector(1 downto 0);
    signal VN208_in3 : std_logic_vector(1 downto 0);
    signal VN208_in4 : std_logic_vector(1 downto 0);
    signal VN208_in5 : std_logic_vector(1 downto 0);
    signal VN209_in0 : std_logic_vector(1 downto 0);
    signal VN209_in1 : std_logic_vector(1 downto 0);
    signal VN209_in2 : std_logic_vector(1 downto 0);
    signal VN209_in3 : std_logic_vector(1 downto 0);
    signal VN209_in4 : std_logic_vector(1 downto 0);
    signal VN209_in5 : std_logic_vector(1 downto 0);
    signal VN210_in0 : std_logic_vector(1 downto 0);
    signal VN210_in1 : std_logic_vector(1 downto 0);
    signal VN210_in2 : std_logic_vector(1 downto 0);
    signal VN210_in3 : std_logic_vector(1 downto 0);
    signal VN210_in4 : std_logic_vector(1 downto 0);
    signal VN210_in5 : std_logic_vector(1 downto 0);
    signal VN211_in0 : std_logic_vector(1 downto 0);
    signal VN211_in1 : std_logic_vector(1 downto 0);
    signal VN211_in2 : std_logic_vector(1 downto 0);
    signal VN211_in3 : std_logic_vector(1 downto 0);
    signal VN211_in4 : std_logic_vector(1 downto 0);
    signal VN211_in5 : std_logic_vector(1 downto 0);
    signal VN212_in0 : std_logic_vector(1 downto 0);
    signal VN212_in1 : std_logic_vector(1 downto 0);
    signal VN212_in2 : std_logic_vector(1 downto 0);
    signal VN212_in3 : std_logic_vector(1 downto 0);
    signal VN212_in4 : std_logic_vector(1 downto 0);
    signal VN212_in5 : std_logic_vector(1 downto 0);
    signal VN213_in0 : std_logic_vector(1 downto 0);
    signal VN213_in1 : std_logic_vector(1 downto 0);
    signal VN213_in2 : std_logic_vector(1 downto 0);
    signal VN213_in3 : std_logic_vector(1 downto 0);
    signal VN213_in4 : std_logic_vector(1 downto 0);
    signal VN213_in5 : std_logic_vector(1 downto 0);
    signal VN214_in0 : std_logic_vector(1 downto 0);
    signal VN214_in1 : std_logic_vector(1 downto 0);
    signal VN214_in2 : std_logic_vector(1 downto 0);
    signal VN214_in3 : std_logic_vector(1 downto 0);
    signal VN214_in4 : std_logic_vector(1 downto 0);
    signal VN214_in5 : std_logic_vector(1 downto 0);
    signal VN215_in0 : std_logic_vector(1 downto 0);
    signal VN215_in1 : std_logic_vector(1 downto 0);
    signal VN215_in2 : std_logic_vector(1 downto 0);
    signal VN215_in3 : std_logic_vector(1 downto 0);
    signal VN215_in4 : std_logic_vector(1 downto 0);
    signal VN215_in5 : std_logic_vector(1 downto 0);
    signal VN216_in0 : std_logic_vector(1 downto 0);
    signal VN216_in1 : std_logic_vector(1 downto 0);
    signal VN216_in2 : std_logic_vector(1 downto 0);
    signal VN216_in3 : std_logic_vector(1 downto 0);
    signal VN216_in4 : std_logic_vector(1 downto 0);
    signal VN216_in5 : std_logic_vector(1 downto 0);
    signal VN217_in0 : std_logic_vector(1 downto 0);
    signal VN217_in1 : std_logic_vector(1 downto 0);
    signal VN217_in2 : std_logic_vector(1 downto 0);
    signal VN217_in3 : std_logic_vector(1 downto 0);
    signal VN217_in4 : std_logic_vector(1 downto 0);
    signal VN217_in5 : std_logic_vector(1 downto 0);
    signal VN218_in0 : std_logic_vector(1 downto 0);
    signal VN218_in1 : std_logic_vector(1 downto 0);
    signal VN218_in2 : std_logic_vector(1 downto 0);
    signal VN218_in3 : std_logic_vector(1 downto 0);
    signal VN218_in4 : std_logic_vector(1 downto 0);
    signal VN218_in5 : std_logic_vector(1 downto 0);
    signal VN219_in0 : std_logic_vector(1 downto 0);
    signal VN219_in1 : std_logic_vector(1 downto 0);
    signal VN219_in2 : std_logic_vector(1 downto 0);
    signal VN219_in3 : std_logic_vector(1 downto 0);
    signal VN219_in4 : std_logic_vector(1 downto 0);
    signal VN219_in5 : std_logic_vector(1 downto 0);
    signal VN220_in0 : std_logic_vector(1 downto 0);
    signal VN220_in1 : std_logic_vector(1 downto 0);
    signal VN220_in2 : std_logic_vector(1 downto 0);
    signal VN220_in3 : std_logic_vector(1 downto 0);
    signal VN220_in4 : std_logic_vector(1 downto 0);
    signal VN220_in5 : std_logic_vector(1 downto 0);
    signal VN221_in0 : std_logic_vector(1 downto 0);
    signal VN221_in1 : std_logic_vector(1 downto 0);
    signal VN221_in2 : std_logic_vector(1 downto 0);
    signal VN221_in3 : std_logic_vector(1 downto 0);
    signal VN221_in4 : std_logic_vector(1 downto 0);
    signal VN221_in5 : std_logic_vector(1 downto 0);
    signal VN222_in0 : std_logic_vector(1 downto 0);
    signal VN222_in1 : std_logic_vector(1 downto 0);
    signal VN222_in2 : std_logic_vector(1 downto 0);
    signal VN222_in3 : std_logic_vector(1 downto 0);
    signal VN222_in4 : std_logic_vector(1 downto 0);
    signal VN222_in5 : std_logic_vector(1 downto 0);
    signal VN223_in0 : std_logic_vector(1 downto 0);
    signal VN223_in1 : std_logic_vector(1 downto 0);
    signal VN223_in2 : std_logic_vector(1 downto 0);
    signal VN223_in3 : std_logic_vector(1 downto 0);
    signal VN223_in4 : std_logic_vector(1 downto 0);
    signal VN223_in5 : std_logic_vector(1 downto 0);
    signal VN224_in0 : std_logic_vector(1 downto 0);
    signal VN224_in1 : std_logic_vector(1 downto 0);
    signal VN224_in2 : std_logic_vector(1 downto 0);
    signal VN224_in3 : std_logic_vector(1 downto 0);
    signal VN224_in4 : std_logic_vector(1 downto 0);
    signal VN224_in5 : std_logic_vector(1 downto 0);
    signal VN225_in0 : std_logic_vector(1 downto 0);
    signal VN225_in1 : std_logic_vector(1 downto 0);
    signal VN225_in2 : std_logic_vector(1 downto 0);
    signal VN225_in3 : std_logic_vector(1 downto 0);
    signal VN225_in4 : std_logic_vector(1 downto 0);
    signal VN225_in5 : std_logic_vector(1 downto 0);
    signal VN226_in0 : std_logic_vector(1 downto 0);
    signal VN226_in1 : std_logic_vector(1 downto 0);
    signal VN226_in2 : std_logic_vector(1 downto 0);
    signal VN226_in3 : std_logic_vector(1 downto 0);
    signal VN226_in4 : std_logic_vector(1 downto 0);
    signal VN226_in5 : std_logic_vector(1 downto 0);
    signal VN227_in0 : std_logic_vector(1 downto 0);
    signal VN227_in1 : std_logic_vector(1 downto 0);
    signal VN227_in2 : std_logic_vector(1 downto 0);
    signal VN227_in3 : std_logic_vector(1 downto 0);
    signal VN227_in4 : std_logic_vector(1 downto 0);
    signal VN227_in5 : std_logic_vector(1 downto 0);
    signal VN228_in0 : std_logic_vector(1 downto 0);
    signal VN228_in1 : std_logic_vector(1 downto 0);
    signal VN228_in2 : std_logic_vector(1 downto 0);
    signal VN228_in3 : std_logic_vector(1 downto 0);
    signal VN228_in4 : std_logic_vector(1 downto 0);
    signal VN228_in5 : std_logic_vector(1 downto 0);
    signal VN229_in0 : std_logic_vector(1 downto 0);
    signal VN229_in1 : std_logic_vector(1 downto 0);
    signal VN229_in2 : std_logic_vector(1 downto 0);
    signal VN229_in3 : std_logic_vector(1 downto 0);
    signal VN229_in4 : std_logic_vector(1 downto 0);
    signal VN229_in5 : std_logic_vector(1 downto 0);
    signal VN230_in0 : std_logic_vector(1 downto 0);
    signal VN230_in1 : std_logic_vector(1 downto 0);
    signal VN230_in2 : std_logic_vector(1 downto 0);
    signal VN230_in3 : std_logic_vector(1 downto 0);
    signal VN230_in4 : std_logic_vector(1 downto 0);
    signal VN230_in5 : std_logic_vector(1 downto 0);
    signal VN231_in0 : std_logic_vector(1 downto 0);
    signal VN231_in1 : std_logic_vector(1 downto 0);
    signal VN231_in2 : std_logic_vector(1 downto 0);
    signal VN231_in3 : std_logic_vector(1 downto 0);
    signal VN231_in4 : std_logic_vector(1 downto 0);
    signal VN231_in5 : std_logic_vector(1 downto 0);
    signal VN232_in0 : std_logic_vector(1 downto 0);
    signal VN232_in1 : std_logic_vector(1 downto 0);
    signal VN232_in2 : std_logic_vector(1 downto 0);
    signal VN232_in3 : std_logic_vector(1 downto 0);
    signal VN232_in4 : std_logic_vector(1 downto 0);
    signal VN232_in5 : std_logic_vector(1 downto 0);
    signal VN233_in0 : std_logic_vector(1 downto 0);
    signal VN233_in1 : std_logic_vector(1 downto 0);
    signal VN233_in2 : std_logic_vector(1 downto 0);
    signal VN233_in3 : std_logic_vector(1 downto 0);
    signal VN233_in4 : std_logic_vector(1 downto 0);
    signal VN233_in5 : std_logic_vector(1 downto 0);
    signal VN234_in0 : std_logic_vector(1 downto 0);
    signal VN234_in1 : std_logic_vector(1 downto 0);
    signal VN234_in2 : std_logic_vector(1 downto 0);
    signal VN234_in3 : std_logic_vector(1 downto 0);
    signal VN234_in4 : std_logic_vector(1 downto 0);
    signal VN234_in5 : std_logic_vector(1 downto 0);
    signal VN235_in0 : std_logic_vector(1 downto 0);
    signal VN235_in1 : std_logic_vector(1 downto 0);
    signal VN235_in2 : std_logic_vector(1 downto 0);
    signal VN235_in3 : std_logic_vector(1 downto 0);
    signal VN235_in4 : std_logic_vector(1 downto 0);
    signal VN235_in5 : std_logic_vector(1 downto 0);
    signal VN236_in0 : std_logic_vector(1 downto 0);
    signal VN236_in1 : std_logic_vector(1 downto 0);
    signal VN236_in2 : std_logic_vector(1 downto 0);
    signal VN236_in3 : std_logic_vector(1 downto 0);
    signal VN236_in4 : std_logic_vector(1 downto 0);
    signal VN236_in5 : std_logic_vector(1 downto 0);
    signal VN237_in0 : std_logic_vector(1 downto 0);
    signal VN237_in1 : std_logic_vector(1 downto 0);
    signal VN237_in2 : std_logic_vector(1 downto 0);
    signal VN237_in3 : std_logic_vector(1 downto 0);
    signal VN237_in4 : std_logic_vector(1 downto 0);
    signal VN237_in5 : std_logic_vector(1 downto 0);
    signal VN238_in0 : std_logic_vector(1 downto 0);
    signal VN238_in1 : std_logic_vector(1 downto 0);
    signal VN238_in2 : std_logic_vector(1 downto 0);
    signal VN238_in3 : std_logic_vector(1 downto 0);
    signal VN238_in4 : std_logic_vector(1 downto 0);
    signal VN238_in5 : std_logic_vector(1 downto 0);
    signal VN239_in0 : std_logic_vector(1 downto 0);
    signal VN239_in1 : std_logic_vector(1 downto 0);
    signal VN239_in2 : std_logic_vector(1 downto 0);
    signal VN239_in3 : std_logic_vector(1 downto 0);
    signal VN239_in4 : std_logic_vector(1 downto 0);
    signal VN239_in5 : std_logic_vector(1 downto 0);
    signal VN240_in0 : std_logic_vector(1 downto 0);
    signal VN240_in1 : std_logic_vector(1 downto 0);
    signal VN240_in2 : std_logic_vector(1 downto 0);
    signal VN240_in3 : std_logic_vector(1 downto 0);
    signal VN240_in4 : std_logic_vector(1 downto 0);
    signal VN240_in5 : std_logic_vector(1 downto 0);
    signal VN241_in0 : std_logic_vector(1 downto 0);
    signal VN241_in1 : std_logic_vector(1 downto 0);
    signal VN241_in2 : std_logic_vector(1 downto 0);
    signal VN241_in3 : std_logic_vector(1 downto 0);
    signal VN241_in4 : std_logic_vector(1 downto 0);
    signal VN241_in5 : std_logic_vector(1 downto 0);
    signal VN242_in0 : std_logic_vector(1 downto 0);
    signal VN242_in1 : std_logic_vector(1 downto 0);
    signal VN242_in2 : std_logic_vector(1 downto 0);
    signal VN242_in3 : std_logic_vector(1 downto 0);
    signal VN242_in4 : std_logic_vector(1 downto 0);
    signal VN242_in5 : std_logic_vector(1 downto 0);
    signal VN243_in0 : std_logic_vector(1 downto 0);
    signal VN243_in1 : std_logic_vector(1 downto 0);
    signal VN243_in2 : std_logic_vector(1 downto 0);
    signal VN243_in3 : std_logic_vector(1 downto 0);
    signal VN243_in4 : std_logic_vector(1 downto 0);
    signal VN243_in5 : std_logic_vector(1 downto 0);
    signal VN244_in0 : std_logic_vector(1 downto 0);
    signal VN244_in1 : std_logic_vector(1 downto 0);
    signal VN244_in2 : std_logic_vector(1 downto 0);
    signal VN244_in3 : std_logic_vector(1 downto 0);
    signal VN244_in4 : std_logic_vector(1 downto 0);
    signal VN244_in5 : std_logic_vector(1 downto 0);
    signal VN245_in0 : std_logic_vector(1 downto 0);
    signal VN245_in1 : std_logic_vector(1 downto 0);
    signal VN245_in2 : std_logic_vector(1 downto 0);
    signal VN245_in3 : std_logic_vector(1 downto 0);
    signal VN245_in4 : std_logic_vector(1 downto 0);
    signal VN245_in5 : std_logic_vector(1 downto 0);
    signal VN246_in0 : std_logic_vector(1 downto 0);
    signal VN246_in1 : std_logic_vector(1 downto 0);
    signal VN246_in2 : std_logic_vector(1 downto 0);
    signal VN246_in3 : std_logic_vector(1 downto 0);
    signal VN246_in4 : std_logic_vector(1 downto 0);
    signal VN246_in5 : std_logic_vector(1 downto 0);
    signal VN247_in0 : std_logic_vector(1 downto 0);
    signal VN247_in1 : std_logic_vector(1 downto 0);
    signal VN247_in2 : std_logic_vector(1 downto 0);
    signal VN247_in3 : std_logic_vector(1 downto 0);
    signal VN247_in4 : std_logic_vector(1 downto 0);
    signal VN247_in5 : std_logic_vector(1 downto 0);
    signal VN248_in0 : std_logic_vector(1 downto 0);
    signal VN248_in1 : std_logic_vector(1 downto 0);
    signal VN248_in2 : std_logic_vector(1 downto 0);
    signal VN248_in3 : std_logic_vector(1 downto 0);
    signal VN248_in4 : std_logic_vector(1 downto 0);
    signal VN248_in5 : std_logic_vector(1 downto 0);
    signal VN249_in0 : std_logic_vector(1 downto 0);
    signal VN249_in1 : std_logic_vector(1 downto 0);
    signal VN249_in2 : std_logic_vector(1 downto 0);
    signal VN249_in3 : std_logic_vector(1 downto 0);
    signal VN249_in4 : std_logic_vector(1 downto 0);
    signal VN249_in5 : std_logic_vector(1 downto 0);
    signal VN250_in0 : std_logic_vector(1 downto 0);
    signal VN250_in1 : std_logic_vector(1 downto 0);
    signal VN250_in2 : std_logic_vector(1 downto 0);
    signal VN250_in3 : std_logic_vector(1 downto 0);
    signal VN250_in4 : std_logic_vector(1 downto 0);
    signal VN250_in5 : std_logic_vector(1 downto 0);
    signal VN251_in0 : std_logic_vector(1 downto 0);
    signal VN251_in1 : std_logic_vector(1 downto 0);
    signal VN251_in2 : std_logic_vector(1 downto 0);
    signal VN251_in3 : std_logic_vector(1 downto 0);
    signal VN251_in4 : std_logic_vector(1 downto 0);
    signal VN251_in5 : std_logic_vector(1 downto 0);
    signal VN252_in0 : std_logic_vector(1 downto 0);
    signal VN252_in1 : std_logic_vector(1 downto 0);
    signal VN252_in2 : std_logic_vector(1 downto 0);
    signal VN252_in3 : std_logic_vector(1 downto 0);
    signal VN252_in4 : std_logic_vector(1 downto 0);
    signal VN252_in5 : std_logic_vector(1 downto 0);
    signal VN253_in0 : std_logic_vector(1 downto 0);
    signal VN253_in1 : std_logic_vector(1 downto 0);
    signal VN253_in2 : std_logic_vector(1 downto 0);
    signal VN253_in3 : std_logic_vector(1 downto 0);
    signal VN253_in4 : std_logic_vector(1 downto 0);
    signal VN253_in5 : std_logic_vector(1 downto 0);
    signal VN254_in0 : std_logic_vector(1 downto 0);
    signal VN254_in1 : std_logic_vector(1 downto 0);
    signal VN254_in2 : std_logic_vector(1 downto 0);
    signal VN254_in3 : std_logic_vector(1 downto 0);
    signal VN254_in4 : std_logic_vector(1 downto 0);
    signal VN254_in5 : std_logic_vector(1 downto 0);
    signal VN255_in0 : std_logic_vector(1 downto 0);
    signal VN255_in1 : std_logic_vector(1 downto 0);
    signal VN255_in2 : std_logic_vector(1 downto 0);
    signal VN255_in3 : std_logic_vector(1 downto 0);
    signal VN255_in4 : std_logic_vector(1 downto 0);
    signal VN255_in5 : std_logic_vector(1 downto 0);
    signal VN256_in0 : std_logic_vector(1 downto 0);
    signal VN256_in1 : std_logic_vector(1 downto 0);
    signal VN256_in2 : std_logic_vector(1 downto 0);
    signal VN256_in3 : std_logic_vector(1 downto 0);
    signal VN256_in4 : std_logic_vector(1 downto 0);
    signal VN256_in5 : std_logic_vector(1 downto 0);
    signal VN257_in0 : std_logic_vector(1 downto 0);
    signal VN257_in1 : std_logic_vector(1 downto 0);
    signal VN257_in2 : std_logic_vector(1 downto 0);
    signal VN257_in3 : std_logic_vector(1 downto 0);
    signal VN257_in4 : std_logic_vector(1 downto 0);
    signal VN257_in5 : std_logic_vector(1 downto 0);
    signal VN258_in0 : std_logic_vector(1 downto 0);
    signal VN258_in1 : std_logic_vector(1 downto 0);
    signal VN258_in2 : std_logic_vector(1 downto 0);
    signal VN258_in3 : std_logic_vector(1 downto 0);
    signal VN258_in4 : std_logic_vector(1 downto 0);
    signal VN258_in5 : std_logic_vector(1 downto 0);
    signal VN259_in0 : std_logic_vector(1 downto 0);
    signal VN259_in1 : std_logic_vector(1 downto 0);
    signal VN259_in2 : std_logic_vector(1 downto 0);
    signal VN259_in3 : std_logic_vector(1 downto 0);
    signal VN259_in4 : std_logic_vector(1 downto 0);
    signal VN259_in5 : std_logic_vector(1 downto 0);
    signal VN260_in0 : std_logic_vector(1 downto 0);
    signal VN260_in1 : std_logic_vector(1 downto 0);
    signal VN260_in2 : std_logic_vector(1 downto 0);
    signal VN260_in3 : std_logic_vector(1 downto 0);
    signal VN260_in4 : std_logic_vector(1 downto 0);
    signal VN260_in5 : std_logic_vector(1 downto 0);
    signal VN261_in0 : std_logic_vector(1 downto 0);
    signal VN261_in1 : std_logic_vector(1 downto 0);
    signal VN261_in2 : std_logic_vector(1 downto 0);
    signal VN261_in3 : std_logic_vector(1 downto 0);
    signal VN261_in4 : std_logic_vector(1 downto 0);
    signal VN261_in5 : std_logic_vector(1 downto 0);
    signal VN262_in0 : std_logic_vector(1 downto 0);
    signal VN262_in1 : std_logic_vector(1 downto 0);
    signal VN262_in2 : std_logic_vector(1 downto 0);
    signal VN262_in3 : std_logic_vector(1 downto 0);
    signal VN262_in4 : std_logic_vector(1 downto 0);
    signal VN262_in5 : std_logic_vector(1 downto 0);
    signal VN263_in0 : std_logic_vector(1 downto 0);
    signal VN263_in1 : std_logic_vector(1 downto 0);
    signal VN263_in2 : std_logic_vector(1 downto 0);
    signal VN263_in3 : std_logic_vector(1 downto 0);
    signal VN263_in4 : std_logic_vector(1 downto 0);
    signal VN263_in5 : std_logic_vector(1 downto 0);
    signal VN264_in0 : std_logic_vector(1 downto 0);
    signal VN264_in1 : std_logic_vector(1 downto 0);
    signal VN264_in2 : std_logic_vector(1 downto 0);
    signal VN264_in3 : std_logic_vector(1 downto 0);
    signal VN264_in4 : std_logic_vector(1 downto 0);
    signal VN264_in5 : std_logic_vector(1 downto 0);
    signal VN265_in0 : std_logic_vector(1 downto 0);
    signal VN265_in1 : std_logic_vector(1 downto 0);
    signal VN265_in2 : std_logic_vector(1 downto 0);
    signal VN265_in3 : std_logic_vector(1 downto 0);
    signal VN265_in4 : std_logic_vector(1 downto 0);
    signal VN265_in5 : std_logic_vector(1 downto 0);
    signal VN266_in0 : std_logic_vector(1 downto 0);
    signal VN266_in1 : std_logic_vector(1 downto 0);
    signal VN266_in2 : std_logic_vector(1 downto 0);
    signal VN266_in3 : std_logic_vector(1 downto 0);
    signal VN266_in4 : std_logic_vector(1 downto 0);
    signal VN266_in5 : std_logic_vector(1 downto 0);
    signal VN267_in0 : std_logic_vector(1 downto 0);
    signal VN267_in1 : std_logic_vector(1 downto 0);
    signal VN267_in2 : std_logic_vector(1 downto 0);
    signal VN267_in3 : std_logic_vector(1 downto 0);
    signal VN267_in4 : std_logic_vector(1 downto 0);
    signal VN267_in5 : std_logic_vector(1 downto 0);
    signal VN268_in0 : std_logic_vector(1 downto 0);
    signal VN268_in1 : std_logic_vector(1 downto 0);
    signal VN268_in2 : std_logic_vector(1 downto 0);
    signal VN268_in3 : std_logic_vector(1 downto 0);
    signal VN268_in4 : std_logic_vector(1 downto 0);
    signal VN268_in5 : std_logic_vector(1 downto 0);
    signal VN269_in0 : std_logic_vector(1 downto 0);
    signal VN269_in1 : std_logic_vector(1 downto 0);
    signal VN269_in2 : std_logic_vector(1 downto 0);
    signal VN269_in3 : std_logic_vector(1 downto 0);
    signal VN269_in4 : std_logic_vector(1 downto 0);
    signal VN269_in5 : std_logic_vector(1 downto 0);
    signal VN270_in0 : std_logic_vector(1 downto 0);
    signal VN270_in1 : std_logic_vector(1 downto 0);
    signal VN270_in2 : std_logic_vector(1 downto 0);
    signal VN270_in3 : std_logic_vector(1 downto 0);
    signal VN270_in4 : std_logic_vector(1 downto 0);
    signal VN270_in5 : std_logic_vector(1 downto 0);
    signal VN271_in0 : std_logic_vector(1 downto 0);
    signal VN271_in1 : std_logic_vector(1 downto 0);
    signal VN271_in2 : std_logic_vector(1 downto 0);
    signal VN271_in3 : std_logic_vector(1 downto 0);
    signal VN271_in4 : std_logic_vector(1 downto 0);
    signal VN271_in5 : std_logic_vector(1 downto 0);
    signal VN272_in0 : std_logic_vector(1 downto 0);
    signal VN272_in1 : std_logic_vector(1 downto 0);
    signal VN272_in2 : std_logic_vector(1 downto 0);
    signal VN272_in3 : std_logic_vector(1 downto 0);
    signal VN272_in4 : std_logic_vector(1 downto 0);
    signal VN272_in5 : std_logic_vector(1 downto 0);
    signal VN273_in0 : std_logic_vector(1 downto 0);
    signal VN273_in1 : std_logic_vector(1 downto 0);
    signal VN273_in2 : std_logic_vector(1 downto 0);
    signal VN273_in3 : std_logic_vector(1 downto 0);
    signal VN273_in4 : std_logic_vector(1 downto 0);
    signal VN273_in5 : std_logic_vector(1 downto 0);
    signal VN274_in0 : std_logic_vector(1 downto 0);
    signal VN274_in1 : std_logic_vector(1 downto 0);
    signal VN274_in2 : std_logic_vector(1 downto 0);
    signal VN274_in3 : std_logic_vector(1 downto 0);
    signal VN274_in4 : std_logic_vector(1 downto 0);
    signal VN274_in5 : std_logic_vector(1 downto 0);
    signal VN275_in0 : std_logic_vector(1 downto 0);
    signal VN275_in1 : std_logic_vector(1 downto 0);
    signal VN275_in2 : std_logic_vector(1 downto 0);
    signal VN275_in3 : std_logic_vector(1 downto 0);
    signal VN275_in4 : std_logic_vector(1 downto 0);
    signal VN275_in5 : std_logic_vector(1 downto 0);
    signal VN276_in0 : std_logic_vector(1 downto 0);
    signal VN276_in1 : std_logic_vector(1 downto 0);
    signal VN276_in2 : std_logic_vector(1 downto 0);
    signal VN276_in3 : std_logic_vector(1 downto 0);
    signal VN276_in4 : std_logic_vector(1 downto 0);
    signal VN276_in5 : std_logic_vector(1 downto 0);
    signal VN277_in0 : std_logic_vector(1 downto 0);
    signal VN277_in1 : std_logic_vector(1 downto 0);
    signal VN277_in2 : std_logic_vector(1 downto 0);
    signal VN277_in3 : std_logic_vector(1 downto 0);
    signal VN277_in4 : std_logic_vector(1 downto 0);
    signal VN277_in5 : std_logic_vector(1 downto 0);
    signal VN278_in0 : std_logic_vector(1 downto 0);
    signal VN278_in1 : std_logic_vector(1 downto 0);
    signal VN278_in2 : std_logic_vector(1 downto 0);
    signal VN278_in3 : std_logic_vector(1 downto 0);
    signal VN278_in4 : std_logic_vector(1 downto 0);
    signal VN278_in5 : std_logic_vector(1 downto 0);
    signal VN279_in0 : std_logic_vector(1 downto 0);
    signal VN279_in1 : std_logic_vector(1 downto 0);
    signal VN279_in2 : std_logic_vector(1 downto 0);
    signal VN279_in3 : std_logic_vector(1 downto 0);
    signal VN279_in4 : std_logic_vector(1 downto 0);
    signal VN279_in5 : std_logic_vector(1 downto 0);
    signal VN280_in0 : std_logic_vector(1 downto 0);
    signal VN280_in1 : std_logic_vector(1 downto 0);
    signal VN280_in2 : std_logic_vector(1 downto 0);
    signal VN280_in3 : std_logic_vector(1 downto 0);
    signal VN280_in4 : std_logic_vector(1 downto 0);
    signal VN280_in5 : std_logic_vector(1 downto 0);
    signal VN281_in0 : std_logic_vector(1 downto 0);
    signal VN281_in1 : std_logic_vector(1 downto 0);
    signal VN281_in2 : std_logic_vector(1 downto 0);
    signal VN281_in3 : std_logic_vector(1 downto 0);
    signal VN281_in4 : std_logic_vector(1 downto 0);
    signal VN281_in5 : std_logic_vector(1 downto 0);
    signal VN282_in0 : std_logic_vector(1 downto 0);
    signal VN282_in1 : std_logic_vector(1 downto 0);
    signal VN282_in2 : std_logic_vector(1 downto 0);
    signal VN282_in3 : std_logic_vector(1 downto 0);
    signal VN282_in4 : std_logic_vector(1 downto 0);
    signal VN282_in5 : std_logic_vector(1 downto 0);
    signal VN283_in0 : std_logic_vector(1 downto 0);
    signal VN283_in1 : std_logic_vector(1 downto 0);
    signal VN283_in2 : std_logic_vector(1 downto 0);
    signal VN283_in3 : std_logic_vector(1 downto 0);
    signal VN283_in4 : std_logic_vector(1 downto 0);
    signal VN283_in5 : std_logic_vector(1 downto 0);
    signal VN284_in0 : std_logic_vector(1 downto 0);
    signal VN284_in1 : std_logic_vector(1 downto 0);
    signal VN284_in2 : std_logic_vector(1 downto 0);
    signal VN284_in3 : std_logic_vector(1 downto 0);
    signal VN284_in4 : std_logic_vector(1 downto 0);
    signal VN284_in5 : std_logic_vector(1 downto 0);
    signal VN285_in0 : std_logic_vector(1 downto 0);
    signal VN285_in1 : std_logic_vector(1 downto 0);
    signal VN285_in2 : std_logic_vector(1 downto 0);
    signal VN285_in3 : std_logic_vector(1 downto 0);
    signal VN285_in4 : std_logic_vector(1 downto 0);
    signal VN285_in5 : std_logic_vector(1 downto 0);
    signal VN286_in0 : std_logic_vector(1 downto 0);
    signal VN286_in1 : std_logic_vector(1 downto 0);
    signal VN286_in2 : std_logic_vector(1 downto 0);
    signal VN286_in3 : std_logic_vector(1 downto 0);
    signal VN286_in4 : std_logic_vector(1 downto 0);
    signal VN286_in5 : std_logic_vector(1 downto 0);
    signal VN287_in0 : std_logic_vector(1 downto 0);
    signal VN287_in1 : std_logic_vector(1 downto 0);
    signal VN287_in2 : std_logic_vector(1 downto 0);
    signal VN287_in3 : std_logic_vector(1 downto 0);
    signal VN287_in4 : std_logic_vector(1 downto 0);
    signal VN287_in5 : std_logic_vector(1 downto 0);
    signal VN288_in0 : std_logic_vector(1 downto 0);
    signal VN288_in1 : std_logic_vector(1 downto 0);
    signal VN288_in2 : std_logic_vector(1 downto 0);
    signal VN288_in3 : std_logic_vector(1 downto 0);
    signal VN288_in4 : std_logic_vector(1 downto 0);
    signal VN288_in5 : std_logic_vector(1 downto 0);
    signal VN289_in0 : std_logic_vector(1 downto 0);
    signal VN289_in1 : std_logic_vector(1 downto 0);
    signal VN289_in2 : std_logic_vector(1 downto 0);
    signal VN289_in3 : std_logic_vector(1 downto 0);
    signal VN289_in4 : std_logic_vector(1 downto 0);
    signal VN289_in5 : std_logic_vector(1 downto 0);
    signal VN290_in0 : std_logic_vector(1 downto 0);
    signal VN290_in1 : std_logic_vector(1 downto 0);
    signal VN290_in2 : std_logic_vector(1 downto 0);
    signal VN290_in3 : std_logic_vector(1 downto 0);
    signal VN290_in4 : std_logic_vector(1 downto 0);
    signal VN290_in5 : std_logic_vector(1 downto 0);
    signal VN291_in0 : std_logic_vector(1 downto 0);
    signal VN291_in1 : std_logic_vector(1 downto 0);
    signal VN291_in2 : std_logic_vector(1 downto 0);
    signal VN291_in3 : std_logic_vector(1 downto 0);
    signal VN291_in4 : std_logic_vector(1 downto 0);
    signal VN291_in5 : std_logic_vector(1 downto 0);
    signal VN292_in0 : std_logic_vector(1 downto 0);
    signal VN292_in1 : std_logic_vector(1 downto 0);
    signal VN292_in2 : std_logic_vector(1 downto 0);
    signal VN292_in3 : std_logic_vector(1 downto 0);
    signal VN292_in4 : std_logic_vector(1 downto 0);
    signal VN292_in5 : std_logic_vector(1 downto 0);
    signal VN293_in0 : std_logic_vector(1 downto 0);
    signal VN293_in1 : std_logic_vector(1 downto 0);
    signal VN293_in2 : std_logic_vector(1 downto 0);
    signal VN293_in3 : std_logic_vector(1 downto 0);
    signal VN293_in4 : std_logic_vector(1 downto 0);
    signal VN293_in5 : std_logic_vector(1 downto 0);
    signal VN294_in0 : std_logic_vector(1 downto 0);
    signal VN294_in1 : std_logic_vector(1 downto 0);
    signal VN294_in2 : std_logic_vector(1 downto 0);
    signal VN294_in3 : std_logic_vector(1 downto 0);
    signal VN294_in4 : std_logic_vector(1 downto 0);
    signal VN294_in5 : std_logic_vector(1 downto 0);
    signal VN295_in0 : std_logic_vector(1 downto 0);
    signal VN295_in1 : std_logic_vector(1 downto 0);
    signal VN295_in2 : std_logic_vector(1 downto 0);
    signal VN295_in3 : std_logic_vector(1 downto 0);
    signal VN295_in4 : std_logic_vector(1 downto 0);
    signal VN295_in5 : std_logic_vector(1 downto 0);
    signal VN296_in0 : std_logic_vector(1 downto 0);
    signal VN296_in1 : std_logic_vector(1 downto 0);
    signal VN296_in2 : std_logic_vector(1 downto 0);
    signal VN296_in3 : std_logic_vector(1 downto 0);
    signal VN296_in4 : std_logic_vector(1 downto 0);
    signal VN296_in5 : std_logic_vector(1 downto 0);
    signal VN297_in0 : std_logic_vector(1 downto 0);
    signal VN297_in1 : std_logic_vector(1 downto 0);
    signal VN297_in2 : std_logic_vector(1 downto 0);
    signal VN297_in3 : std_logic_vector(1 downto 0);
    signal VN297_in4 : std_logic_vector(1 downto 0);
    signal VN297_in5 : std_logic_vector(1 downto 0);
    signal VN298_in0 : std_logic_vector(1 downto 0);
    signal VN298_in1 : std_logic_vector(1 downto 0);
    signal VN298_in2 : std_logic_vector(1 downto 0);
    signal VN298_in3 : std_logic_vector(1 downto 0);
    signal VN298_in4 : std_logic_vector(1 downto 0);
    signal VN298_in5 : std_logic_vector(1 downto 0);
    signal VN299_in0 : std_logic_vector(1 downto 0);
    signal VN299_in1 : std_logic_vector(1 downto 0);
    signal VN299_in2 : std_logic_vector(1 downto 0);
    signal VN299_in3 : std_logic_vector(1 downto 0);
    signal VN299_in4 : std_logic_vector(1 downto 0);
    signal VN299_in5 : std_logic_vector(1 downto 0);
    signal VN300_in0 : std_logic_vector(1 downto 0);
    signal VN300_in1 : std_logic_vector(1 downto 0);
    signal VN300_in2 : std_logic_vector(1 downto 0);
    signal VN300_in3 : std_logic_vector(1 downto 0);
    signal VN300_in4 : std_logic_vector(1 downto 0);
    signal VN300_in5 : std_logic_vector(1 downto 0);
    signal VN301_in0 : std_logic_vector(1 downto 0);
    signal VN301_in1 : std_logic_vector(1 downto 0);
    signal VN301_in2 : std_logic_vector(1 downto 0);
    signal VN301_in3 : std_logic_vector(1 downto 0);
    signal VN301_in4 : std_logic_vector(1 downto 0);
    signal VN301_in5 : std_logic_vector(1 downto 0);
    signal VN302_in0 : std_logic_vector(1 downto 0);
    signal VN302_in1 : std_logic_vector(1 downto 0);
    signal VN302_in2 : std_logic_vector(1 downto 0);
    signal VN302_in3 : std_logic_vector(1 downto 0);
    signal VN302_in4 : std_logic_vector(1 downto 0);
    signal VN302_in5 : std_logic_vector(1 downto 0);
    signal VN303_in0 : std_logic_vector(1 downto 0);
    signal VN303_in1 : std_logic_vector(1 downto 0);
    signal VN303_in2 : std_logic_vector(1 downto 0);
    signal VN303_in3 : std_logic_vector(1 downto 0);
    signal VN303_in4 : std_logic_vector(1 downto 0);
    signal VN303_in5 : std_logic_vector(1 downto 0);
    signal VN304_in0 : std_logic_vector(1 downto 0);
    signal VN304_in1 : std_logic_vector(1 downto 0);
    signal VN304_in2 : std_logic_vector(1 downto 0);
    signal VN304_in3 : std_logic_vector(1 downto 0);
    signal VN304_in4 : std_logic_vector(1 downto 0);
    signal VN304_in5 : std_logic_vector(1 downto 0);
    signal VN305_in0 : std_logic_vector(1 downto 0);
    signal VN305_in1 : std_logic_vector(1 downto 0);
    signal VN305_in2 : std_logic_vector(1 downto 0);
    signal VN305_in3 : std_logic_vector(1 downto 0);
    signal VN305_in4 : std_logic_vector(1 downto 0);
    signal VN305_in5 : std_logic_vector(1 downto 0);
    signal VN306_in0 : std_logic_vector(1 downto 0);
    signal VN306_in1 : std_logic_vector(1 downto 0);
    signal VN306_in2 : std_logic_vector(1 downto 0);
    signal VN306_in3 : std_logic_vector(1 downto 0);
    signal VN306_in4 : std_logic_vector(1 downto 0);
    signal VN306_in5 : std_logic_vector(1 downto 0);
    signal VN307_in0 : std_logic_vector(1 downto 0);
    signal VN307_in1 : std_logic_vector(1 downto 0);
    signal VN307_in2 : std_logic_vector(1 downto 0);
    signal VN307_in3 : std_logic_vector(1 downto 0);
    signal VN307_in4 : std_logic_vector(1 downto 0);
    signal VN307_in5 : std_logic_vector(1 downto 0);
    signal VN308_in0 : std_logic_vector(1 downto 0);
    signal VN308_in1 : std_logic_vector(1 downto 0);
    signal VN308_in2 : std_logic_vector(1 downto 0);
    signal VN308_in3 : std_logic_vector(1 downto 0);
    signal VN308_in4 : std_logic_vector(1 downto 0);
    signal VN308_in5 : std_logic_vector(1 downto 0);
    signal VN309_in0 : std_logic_vector(1 downto 0);
    signal VN309_in1 : std_logic_vector(1 downto 0);
    signal VN309_in2 : std_logic_vector(1 downto 0);
    signal VN309_in3 : std_logic_vector(1 downto 0);
    signal VN309_in4 : std_logic_vector(1 downto 0);
    signal VN309_in5 : std_logic_vector(1 downto 0);
    signal VN310_in0 : std_logic_vector(1 downto 0);
    signal VN310_in1 : std_logic_vector(1 downto 0);
    signal VN310_in2 : std_logic_vector(1 downto 0);
    signal VN310_in3 : std_logic_vector(1 downto 0);
    signal VN310_in4 : std_logic_vector(1 downto 0);
    signal VN310_in5 : std_logic_vector(1 downto 0);
    signal VN311_in0 : std_logic_vector(1 downto 0);
    signal VN311_in1 : std_logic_vector(1 downto 0);
    signal VN311_in2 : std_logic_vector(1 downto 0);
    signal VN311_in3 : std_logic_vector(1 downto 0);
    signal VN311_in4 : std_logic_vector(1 downto 0);
    signal VN311_in5 : std_logic_vector(1 downto 0);
    signal VN312_in0 : std_logic_vector(1 downto 0);
    signal VN312_in1 : std_logic_vector(1 downto 0);
    signal VN312_in2 : std_logic_vector(1 downto 0);
    signal VN312_in3 : std_logic_vector(1 downto 0);
    signal VN312_in4 : std_logic_vector(1 downto 0);
    signal VN312_in5 : std_logic_vector(1 downto 0);
    signal VN313_in0 : std_logic_vector(1 downto 0);
    signal VN313_in1 : std_logic_vector(1 downto 0);
    signal VN313_in2 : std_logic_vector(1 downto 0);
    signal VN313_in3 : std_logic_vector(1 downto 0);
    signal VN313_in4 : std_logic_vector(1 downto 0);
    signal VN313_in5 : std_logic_vector(1 downto 0);
    signal VN314_in0 : std_logic_vector(1 downto 0);
    signal VN314_in1 : std_logic_vector(1 downto 0);
    signal VN314_in2 : std_logic_vector(1 downto 0);
    signal VN314_in3 : std_logic_vector(1 downto 0);
    signal VN314_in4 : std_logic_vector(1 downto 0);
    signal VN314_in5 : std_logic_vector(1 downto 0);
    signal VN315_in0 : std_logic_vector(1 downto 0);
    signal VN315_in1 : std_logic_vector(1 downto 0);
    signal VN315_in2 : std_logic_vector(1 downto 0);
    signal VN315_in3 : std_logic_vector(1 downto 0);
    signal VN315_in4 : std_logic_vector(1 downto 0);
    signal VN315_in5 : std_logic_vector(1 downto 0);
    signal VN316_in0 : std_logic_vector(1 downto 0);
    signal VN316_in1 : std_logic_vector(1 downto 0);
    signal VN316_in2 : std_logic_vector(1 downto 0);
    signal VN316_in3 : std_logic_vector(1 downto 0);
    signal VN316_in4 : std_logic_vector(1 downto 0);
    signal VN316_in5 : std_logic_vector(1 downto 0);
    signal VN317_in0 : std_logic_vector(1 downto 0);
    signal VN317_in1 : std_logic_vector(1 downto 0);
    signal VN317_in2 : std_logic_vector(1 downto 0);
    signal VN317_in3 : std_logic_vector(1 downto 0);
    signal VN317_in4 : std_logic_vector(1 downto 0);
    signal VN317_in5 : std_logic_vector(1 downto 0);
    signal VN318_in0 : std_logic_vector(1 downto 0);
    signal VN318_in1 : std_logic_vector(1 downto 0);
    signal VN318_in2 : std_logic_vector(1 downto 0);
    signal VN318_in3 : std_logic_vector(1 downto 0);
    signal VN318_in4 : std_logic_vector(1 downto 0);
    signal VN318_in5 : std_logic_vector(1 downto 0);
    signal VN319_in0 : std_logic_vector(1 downto 0);
    signal VN319_in1 : std_logic_vector(1 downto 0);
    signal VN319_in2 : std_logic_vector(1 downto 0);
    signal VN319_in3 : std_logic_vector(1 downto 0);
    signal VN319_in4 : std_logic_vector(1 downto 0);
    signal VN319_in5 : std_logic_vector(1 downto 0);
    signal VN320_in0 : std_logic_vector(1 downto 0);
    signal VN320_in1 : std_logic_vector(1 downto 0);
    signal VN320_in2 : std_logic_vector(1 downto 0);
    signal VN320_in3 : std_logic_vector(1 downto 0);
    signal VN320_in4 : std_logic_vector(1 downto 0);
    signal VN320_in5 : std_logic_vector(1 downto 0);
    signal VN321_in0 : std_logic_vector(1 downto 0);
    signal VN321_in1 : std_logic_vector(1 downto 0);
    signal VN321_in2 : std_logic_vector(1 downto 0);
    signal VN321_in3 : std_logic_vector(1 downto 0);
    signal VN321_in4 : std_logic_vector(1 downto 0);
    signal VN321_in5 : std_logic_vector(1 downto 0);
    signal VN322_in0 : std_logic_vector(1 downto 0);
    signal VN322_in1 : std_logic_vector(1 downto 0);
    signal VN322_in2 : std_logic_vector(1 downto 0);
    signal VN322_in3 : std_logic_vector(1 downto 0);
    signal VN322_in4 : std_logic_vector(1 downto 0);
    signal VN322_in5 : std_logic_vector(1 downto 0);
    signal VN323_in0 : std_logic_vector(1 downto 0);
    signal VN323_in1 : std_logic_vector(1 downto 0);
    signal VN323_in2 : std_logic_vector(1 downto 0);
    signal VN323_in3 : std_logic_vector(1 downto 0);
    signal VN323_in4 : std_logic_vector(1 downto 0);
    signal VN323_in5 : std_logic_vector(1 downto 0);
    signal VN324_in0 : std_logic_vector(1 downto 0);
    signal VN324_in1 : std_logic_vector(1 downto 0);
    signal VN324_in2 : std_logic_vector(1 downto 0);
    signal VN324_in3 : std_logic_vector(1 downto 0);
    signal VN324_in4 : std_logic_vector(1 downto 0);
    signal VN324_in5 : std_logic_vector(1 downto 0);
    signal VN325_in0 : std_logic_vector(1 downto 0);
    signal VN325_in1 : std_logic_vector(1 downto 0);
    signal VN325_in2 : std_logic_vector(1 downto 0);
    signal VN325_in3 : std_logic_vector(1 downto 0);
    signal VN325_in4 : std_logic_vector(1 downto 0);
    signal VN325_in5 : std_logic_vector(1 downto 0);
    signal VN326_in0 : std_logic_vector(1 downto 0);
    signal VN326_in1 : std_logic_vector(1 downto 0);
    signal VN326_in2 : std_logic_vector(1 downto 0);
    signal VN326_in3 : std_logic_vector(1 downto 0);
    signal VN326_in4 : std_logic_vector(1 downto 0);
    signal VN326_in5 : std_logic_vector(1 downto 0);
    signal VN327_in0 : std_logic_vector(1 downto 0);
    signal VN327_in1 : std_logic_vector(1 downto 0);
    signal VN327_in2 : std_logic_vector(1 downto 0);
    signal VN327_in3 : std_logic_vector(1 downto 0);
    signal VN327_in4 : std_logic_vector(1 downto 0);
    signal VN327_in5 : std_logic_vector(1 downto 0);
    signal VN328_in0 : std_logic_vector(1 downto 0);
    signal VN328_in1 : std_logic_vector(1 downto 0);
    signal VN328_in2 : std_logic_vector(1 downto 0);
    signal VN328_in3 : std_logic_vector(1 downto 0);
    signal VN328_in4 : std_logic_vector(1 downto 0);
    signal VN328_in5 : std_logic_vector(1 downto 0);
    signal VN329_in0 : std_logic_vector(1 downto 0);
    signal VN329_in1 : std_logic_vector(1 downto 0);
    signal VN329_in2 : std_logic_vector(1 downto 0);
    signal VN329_in3 : std_logic_vector(1 downto 0);
    signal VN329_in4 : std_logic_vector(1 downto 0);
    signal VN329_in5 : std_logic_vector(1 downto 0);
    signal VN330_in0 : std_logic_vector(1 downto 0);
    signal VN330_in1 : std_logic_vector(1 downto 0);
    signal VN330_in2 : std_logic_vector(1 downto 0);
    signal VN330_in3 : std_logic_vector(1 downto 0);
    signal VN330_in4 : std_logic_vector(1 downto 0);
    signal VN330_in5 : std_logic_vector(1 downto 0);
    signal VN331_in0 : std_logic_vector(1 downto 0);
    signal VN331_in1 : std_logic_vector(1 downto 0);
    signal VN331_in2 : std_logic_vector(1 downto 0);
    signal VN331_in3 : std_logic_vector(1 downto 0);
    signal VN331_in4 : std_logic_vector(1 downto 0);
    signal VN331_in5 : std_logic_vector(1 downto 0);
    signal VN332_in0 : std_logic_vector(1 downto 0);
    signal VN332_in1 : std_logic_vector(1 downto 0);
    signal VN332_in2 : std_logic_vector(1 downto 0);
    signal VN332_in3 : std_logic_vector(1 downto 0);
    signal VN332_in4 : std_logic_vector(1 downto 0);
    signal VN332_in5 : std_logic_vector(1 downto 0);
    signal VN333_in0 : std_logic_vector(1 downto 0);
    signal VN333_in1 : std_logic_vector(1 downto 0);
    signal VN333_in2 : std_logic_vector(1 downto 0);
    signal VN333_in3 : std_logic_vector(1 downto 0);
    signal VN333_in4 : std_logic_vector(1 downto 0);
    signal VN333_in5 : std_logic_vector(1 downto 0);
    signal VN334_in0 : std_logic_vector(1 downto 0);
    signal VN334_in1 : std_logic_vector(1 downto 0);
    signal VN334_in2 : std_logic_vector(1 downto 0);
    signal VN334_in3 : std_logic_vector(1 downto 0);
    signal VN334_in4 : std_logic_vector(1 downto 0);
    signal VN334_in5 : std_logic_vector(1 downto 0);
    signal VN335_in0 : std_logic_vector(1 downto 0);
    signal VN335_in1 : std_logic_vector(1 downto 0);
    signal VN335_in2 : std_logic_vector(1 downto 0);
    signal VN335_in3 : std_logic_vector(1 downto 0);
    signal VN335_in4 : std_logic_vector(1 downto 0);
    signal VN335_in5 : std_logic_vector(1 downto 0);
    signal VN336_in0 : std_logic_vector(1 downto 0);
    signal VN336_in1 : std_logic_vector(1 downto 0);
    signal VN336_in2 : std_logic_vector(1 downto 0);
    signal VN336_in3 : std_logic_vector(1 downto 0);
    signal VN336_in4 : std_logic_vector(1 downto 0);
    signal VN336_in5 : std_logic_vector(1 downto 0);
    signal VN337_in0 : std_logic_vector(1 downto 0);
    signal VN337_in1 : std_logic_vector(1 downto 0);
    signal VN337_in2 : std_logic_vector(1 downto 0);
    signal VN337_in3 : std_logic_vector(1 downto 0);
    signal VN337_in4 : std_logic_vector(1 downto 0);
    signal VN337_in5 : std_logic_vector(1 downto 0);
    signal VN338_in0 : std_logic_vector(1 downto 0);
    signal VN338_in1 : std_logic_vector(1 downto 0);
    signal VN338_in2 : std_logic_vector(1 downto 0);
    signal VN338_in3 : std_logic_vector(1 downto 0);
    signal VN338_in4 : std_logic_vector(1 downto 0);
    signal VN338_in5 : std_logic_vector(1 downto 0);
    signal VN339_in0 : std_logic_vector(1 downto 0);
    signal VN339_in1 : std_logic_vector(1 downto 0);
    signal VN339_in2 : std_logic_vector(1 downto 0);
    signal VN339_in3 : std_logic_vector(1 downto 0);
    signal VN339_in4 : std_logic_vector(1 downto 0);
    signal VN339_in5 : std_logic_vector(1 downto 0);
    signal VN340_in0 : std_logic_vector(1 downto 0);
    signal VN340_in1 : std_logic_vector(1 downto 0);
    signal VN340_in2 : std_logic_vector(1 downto 0);
    signal VN340_in3 : std_logic_vector(1 downto 0);
    signal VN340_in4 : std_logic_vector(1 downto 0);
    signal VN340_in5 : std_logic_vector(1 downto 0);
    signal VN341_in0 : std_logic_vector(1 downto 0);
    signal VN341_in1 : std_logic_vector(1 downto 0);
    signal VN341_in2 : std_logic_vector(1 downto 0);
    signal VN341_in3 : std_logic_vector(1 downto 0);
    signal VN341_in4 : std_logic_vector(1 downto 0);
    signal VN341_in5 : std_logic_vector(1 downto 0);
    signal VN342_in0 : std_logic_vector(1 downto 0);
    signal VN342_in1 : std_logic_vector(1 downto 0);
    signal VN342_in2 : std_logic_vector(1 downto 0);
    signal VN342_in3 : std_logic_vector(1 downto 0);
    signal VN342_in4 : std_logic_vector(1 downto 0);
    signal VN342_in5 : std_logic_vector(1 downto 0);
    signal VN343_in0 : std_logic_vector(1 downto 0);
    signal VN343_in1 : std_logic_vector(1 downto 0);
    signal VN343_in2 : std_logic_vector(1 downto 0);
    signal VN343_in3 : std_logic_vector(1 downto 0);
    signal VN343_in4 : std_logic_vector(1 downto 0);
    signal VN343_in5 : std_logic_vector(1 downto 0);
    signal VN344_in0 : std_logic_vector(1 downto 0);
    signal VN344_in1 : std_logic_vector(1 downto 0);
    signal VN344_in2 : std_logic_vector(1 downto 0);
    signal VN344_in3 : std_logic_vector(1 downto 0);
    signal VN344_in4 : std_logic_vector(1 downto 0);
    signal VN344_in5 : std_logic_vector(1 downto 0);
    signal VN345_in0 : std_logic_vector(1 downto 0);
    signal VN345_in1 : std_logic_vector(1 downto 0);
    signal VN345_in2 : std_logic_vector(1 downto 0);
    signal VN345_in3 : std_logic_vector(1 downto 0);
    signal VN345_in4 : std_logic_vector(1 downto 0);
    signal VN345_in5 : std_logic_vector(1 downto 0);
    signal VN346_in0 : std_logic_vector(1 downto 0);
    signal VN346_in1 : std_logic_vector(1 downto 0);
    signal VN346_in2 : std_logic_vector(1 downto 0);
    signal VN346_in3 : std_logic_vector(1 downto 0);
    signal VN346_in4 : std_logic_vector(1 downto 0);
    signal VN346_in5 : std_logic_vector(1 downto 0);
    signal VN347_in0 : std_logic_vector(1 downto 0);
    signal VN347_in1 : std_logic_vector(1 downto 0);
    signal VN347_in2 : std_logic_vector(1 downto 0);
    signal VN347_in3 : std_logic_vector(1 downto 0);
    signal VN347_in4 : std_logic_vector(1 downto 0);
    signal VN347_in5 : std_logic_vector(1 downto 0);
    signal VN348_in0 : std_logic_vector(1 downto 0);
    signal VN348_in1 : std_logic_vector(1 downto 0);
    signal VN348_in2 : std_logic_vector(1 downto 0);
    signal VN348_in3 : std_logic_vector(1 downto 0);
    signal VN348_in4 : std_logic_vector(1 downto 0);
    signal VN348_in5 : std_logic_vector(1 downto 0);
    signal VN349_in0 : std_logic_vector(1 downto 0);
    signal VN349_in1 : std_logic_vector(1 downto 0);
    signal VN349_in2 : std_logic_vector(1 downto 0);
    signal VN349_in3 : std_logic_vector(1 downto 0);
    signal VN349_in4 : std_logic_vector(1 downto 0);
    signal VN349_in5 : std_logic_vector(1 downto 0);
    signal VN350_in0 : std_logic_vector(1 downto 0);
    signal VN350_in1 : std_logic_vector(1 downto 0);
    signal VN350_in2 : std_logic_vector(1 downto 0);
    signal VN350_in3 : std_logic_vector(1 downto 0);
    signal VN350_in4 : std_logic_vector(1 downto 0);
    signal VN350_in5 : std_logic_vector(1 downto 0);
    signal VN351_in0 : std_logic_vector(1 downto 0);
    signal VN351_in1 : std_logic_vector(1 downto 0);
    signal VN351_in2 : std_logic_vector(1 downto 0);
    signal VN351_in3 : std_logic_vector(1 downto 0);
    signal VN351_in4 : std_logic_vector(1 downto 0);
    signal VN351_in5 : std_logic_vector(1 downto 0);
    signal VN352_in0 : std_logic_vector(1 downto 0);
    signal VN352_in1 : std_logic_vector(1 downto 0);
    signal VN352_in2 : std_logic_vector(1 downto 0);
    signal VN352_in3 : std_logic_vector(1 downto 0);
    signal VN352_in4 : std_logic_vector(1 downto 0);
    signal VN352_in5 : std_logic_vector(1 downto 0);
    signal VN353_in0 : std_logic_vector(1 downto 0);
    signal VN353_in1 : std_logic_vector(1 downto 0);
    signal VN353_in2 : std_logic_vector(1 downto 0);
    signal VN353_in3 : std_logic_vector(1 downto 0);
    signal VN353_in4 : std_logic_vector(1 downto 0);
    signal VN353_in5 : std_logic_vector(1 downto 0);
    signal VN354_in0 : std_logic_vector(1 downto 0);
    signal VN354_in1 : std_logic_vector(1 downto 0);
    signal VN354_in2 : std_logic_vector(1 downto 0);
    signal VN354_in3 : std_logic_vector(1 downto 0);
    signal VN354_in4 : std_logic_vector(1 downto 0);
    signal VN354_in5 : std_logic_vector(1 downto 0);
    signal VN355_in0 : std_logic_vector(1 downto 0);
    signal VN355_in1 : std_logic_vector(1 downto 0);
    signal VN355_in2 : std_logic_vector(1 downto 0);
    signal VN355_in3 : std_logic_vector(1 downto 0);
    signal VN355_in4 : std_logic_vector(1 downto 0);
    signal VN355_in5 : std_logic_vector(1 downto 0);
    signal VN356_in0 : std_logic_vector(1 downto 0);
    signal VN356_in1 : std_logic_vector(1 downto 0);
    signal VN356_in2 : std_logic_vector(1 downto 0);
    signal VN356_in3 : std_logic_vector(1 downto 0);
    signal VN356_in4 : std_logic_vector(1 downto 0);
    signal VN356_in5 : std_logic_vector(1 downto 0);
    signal VN357_in0 : std_logic_vector(1 downto 0);
    signal VN357_in1 : std_logic_vector(1 downto 0);
    signal VN357_in2 : std_logic_vector(1 downto 0);
    signal VN357_in3 : std_logic_vector(1 downto 0);
    signal VN357_in4 : std_logic_vector(1 downto 0);
    signal VN357_in5 : std_logic_vector(1 downto 0);
    signal VN358_in0 : std_logic_vector(1 downto 0);
    signal VN358_in1 : std_logic_vector(1 downto 0);
    signal VN358_in2 : std_logic_vector(1 downto 0);
    signal VN358_in3 : std_logic_vector(1 downto 0);
    signal VN358_in4 : std_logic_vector(1 downto 0);
    signal VN358_in5 : std_logic_vector(1 downto 0);
    signal VN359_in0 : std_logic_vector(1 downto 0);
    signal VN359_in1 : std_logic_vector(1 downto 0);
    signal VN359_in2 : std_logic_vector(1 downto 0);
    signal VN359_in3 : std_logic_vector(1 downto 0);
    signal VN359_in4 : std_logic_vector(1 downto 0);
    signal VN359_in5 : std_logic_vector(1 downto 0);
    signal VN360_in0 : std_logic_vector(1 downto 0);
    signal VN360_in1 : std_logic_vector(1 downto 0);
    signal VN360_in2 : std_logic_vector(1 downto 0);
    signal VN360_in3 : std_logic_vector(1 downto 0);
    signal VN360_in4 : std_logic_vector(1 downto 0);
    signal VN360_in5 : std_logic_vector(1 downto 0);
    signal VN361_in0 : std_logic_vector(1 downto 0);
    signal VN361_in1 : std_logic_vector(1 downto 0);
    signal VN361_in2 : std_logic_vector(1 downto 0);
    signal VN361_in3 : std_logic_vector(1 downto 0);
    signal VN361_in4 : std_logic_vector(1 downto 0);
    signal VN361_in5 : std_logic_vector(1 downto 0);
    signal VN362_in0 : std_logic_vector(1 downto 0);
    signal VN362_in1 : std_logic_vector(1 downto 0);
    signal VN362_in2 : std_logic_vector(1 downto 0);
    signal VN362_in3 : std_logic_vector(1 downto 0);
    signal VN362_in4 : std_logic_vector(1 downto 0);
    signal VN362_in5 : std_logic_vector(1 downto 0);
    signal VN363_in0 : std_logic_vector(1 downto 0);
    signal VN363_in1 : std_logic_vector(1 downto 0);
    signal VN363_in2 : std_logic_vector(1 downto 0);
    signal VN363_in3 : std_logic_vector(1 downto 0);
    signal VN363_in4 : std_logic_vector(1 downto 0);
    signal VN363_in5 : std_logic_vector(1 downto 0);
    signal VN364_in0 : std_logic_vector(1 downto 0);
    signal VN364_in1 : std_logic_vector(1 downto 0);
    signal VN364_in2 : std_logic_vector(1 downto 0);
    signal VN364_in3 : std_logic_vector(1 downto 0);
    signal VN364_in4 : std_logic_vector(1 downto 0);
    signal VN364_in5 : std_logic_vector(1 downto 0);
    signal VN365_in0 : std_logic_vector(1 downto 0);
    signal VN365_in1 : std_logic_vector(1 downto 0);
    signal VN365_in2 : std_logic_vector(1 downto 0);
    signal VN365_in3 : std_logic_vector(1 downto 0);
    signal VN365_in4 : std_logic_vector(1 downto 0);
    signal VN365_in5 : std_logic_vector(1 downto 0);
    signal VN366_in0 : std_logic_vector(1 downto 0);
    signal VN366_in1 : std_logic_vector(1 downto 0);
    signal VN366_in2 : std_logic_vector(1 downto 0);
    signal VN366_in3 : std_logic_vector(1 downto 0);
    signal VN366_in4 : std_logic_vector(1 downto 0);
    signal VN366_in5 : std_logic_vector(1 downto 0);
    signal VN367_in0 : std_logic_vector(1 downto 0);
    signal VN367_in1 : std_logic_vector(1 downto 0);
    signal VN367_in2 : std_logic_vector(1 downto 0);
    signal VN367_in3 : std_logic_vector(1 downto 0);
    signal VN367_in4 : std_logic_vector(1 downto 0);
    signal VN367_in5 : std_logic_vector(1 downto 0);
    signal VN368_in0 : std_logic_vector(1 downto 0);
    signal VN368_in1 : std_logic_vector(1 downto 0);
    signal VN368_in2 : std_logic_vector(1 downto 0);
    signal VN368_in3 : std_logic_vector(1 downto 0);
    signal VN368_in4 : std_logic_vector(1 downto 0);
    signal VN368_in5 : std_logic_vector(1 downto 0);
    signal VN369_in0 : std_logic_vector(1 downto 0);
    signal VN369_in1 : std_logic_vector(1 downto 0);
    signal VN369_in2 : std_logic_vector(1 downto 0);
    signal VN369_in3 : std_logic_vector(1 downto 0);
    signal VN369_in4 : std_logic_vector(1 downto 0);
    signal VN369_in5 : std_logic_vector(1 downto 0);
    signal VN370_in0 : std_logic_vector(1 downto 0);
    signal VN370_in1 : std_logic_vector(1 downto 0);
    signal VN370_in2 : std_logic_vector(1 downto 0);
    signal VN370_in3 : std_logic_vector(1 downto 0);
    signal VN370_in4 : std_logic_vector(1 downto 0);
    signal VN370_in5 : std_logic_vector(1 downto 0);
    signal VN371_in0 : std_logic_vector(1 downto 0);
    signal VN371_in1 : std_logic_vector(1 downto 0);
    signal VN371_in2 : std_logic_vector(1 downto 0);
    signal VN371_in3 : std_logic_vector(1 downto 0);
    signal VN371_in4 : std_logic_vector(1 downto 0);
    signal VN371_in5 : std_logic_vector(1 downto 0);
    signal VN372_in0 : std_logic_vector(1 downto 0);
    signal VN372_in1 : std_logic_vector(1 downto 0);
    signal VN372_in2 : std_logic_vector(1 downto 0);
    signal VN372_in3 : std_logic_vector(1 downto 0);
    signal VN372_in4 : std_logic_vector(1 downto 0);
    signal VN372_in5 : std_logic_vector(1 downto 0);
    signal VN373_in0 : std_logic_vector(1 downto 0);
    signal VN373_in1 : std_logic_vector(1 downto 0);
    signal VN373_in2 : std_logic_vector(1 downto 0);
    signal VN373_in3 : std_logic_vector(1 downto 0);
    signal VN373_in4 : std_logic_vector(1 downto 0);
    signal VN373_in5 : std_logic_vector(1 downto 0);
    signal VN374_in0 : std_logic_vector(1 downto 0);
    signal VN374_in1 : std_logic_vector(1 downto 0);
    signal VN374_in2 : std_logic_vector(1 downto 0);
    signal VN374_in3 : std_logic_vector(1 downto 0);
    signal VN374_in4 : std_logic_vector(1 downto 0);
    signal VN374_in5 : std_logic_vector(1 downto 0);
    signal VN375_in0 : std_logic_vector(1 downto 0);
    signal VN375_in1 : std_logic_vector(1 downto 0);
    signal VN375_in2 : std_logic_vector(1 downto 0);
    signal VN375_in3 : std_logic_vector(1 downto 0);
    signal VN375_in4 : std_logic_vector(1 downto 0);
    signal VN375_in5 : std_logic_vector(1 downto 0);
    signal VN376_in0 : std_logic_vector(1 downto 0);
    signal VN376_in1 : std_logic_vector(1 downto 0);
    signal VN376_in2 : std_logic_vector(1 downto 0);
    signal VN376_in3 : std_logic_vector(1 downto 0);
    signal VN376_in4 : std_logic_vector(1 downto 0);
    signal VN376_in5 : std_logic_vector(1 downto 0);
    signal VN377_in0 : std_logic_vector(1 downto 0);
    signal VN377_in1 : std_logic_vector(1 downto 0);
    signal VN377_in2 : std_logic_vector(1 downto 0);
    signal VN377_in3 : std_logic_vector(1 downto 0);
    signal VN377_in4 : std_logic_vector(1 downto 0);
    signal VN377_in5 : std_logic_vector(1 downto 0);
    signal VN378_in0 : std_logic_vector(1 downto 0);
    signal VN378_in1 : std_logic_vector(1 downto 0);
    signal VN378_in2 : std_logic_vector(1 downto 0);
    signal VN378_in3 : std_logic_vector(1 downto 0);
    signal VN378_in4 : std_logic_vector(1 downto 0);
    signal VN378_in5 : std_logic_vector(1 downto 0);
    signal VN379_in0 : std_logic_vector(1 downto 0);
    signal VN379_in1 : std_logic_vector(1 downto 0);
    signal VN379_in2 : std_logic_vector(1 downto 0);
    signal VN379_in3 : std_logic_vector(1 downto 0);
    signal VN379_in4 : std_logic_vector(1 downto 0);
    signal VN379_in5 : std_logic_vector(1 downto 0);
    signal VN380_in0 : std_logic_vector(1 downto 0);
    signal VN380_in1 : std_logic_vector(1 downto 0);
    signal VN380_in2 : std_logic_vector(1 downto 0);
    signal VN380_in3 : std_logic_vector(1 downto 0);
    signal VN380_in4 : std_logic_vector(1 downto 0);
    signal VN380_in5 : std_logic_vector(1 downto 0);
    signal VN381_in0 : std_logic_vector(1 downto 0);
    signal VN381_in1 : std_logic_vector(1 downto 0);
    signal VN381_in2 : std_logic_vector(1 downto 0);
    signal VN381_in3 : std_logic_vector(1 downto 0);
    signal VN381_in4 : std_logic_vector(1 downto 0);
    signal VN381_in5 : std_logic_vector(1 downto 0);
    signal VN382_in0 : std_logic_vector(1 downto 0);
    signal VN382_in1 : std_logic_vector(1 downto 0);
    signal VN382_in2 : std_logic_vector(1 downto 0);
    signal VN382_in3 : std_logic_vector(1 downto 0);
    signal VN382_in4 : std_logic_vector(1 downto 0);
    signal VN382_in5 : std_logic_vector(1 downto 0);
    signal VN383_in0 : std_logic_vector(1 downto 0);
    signal VN383_in1 : std_logic_vector(1 downto 0);
    signal VN383_in2 : std_logic_vector(1 downto 0);
    signal VN383_in3 : std_logic_vector(1 downto 0);
    signal VN383_in4 : std_logic_vector(1 downto 0);
    signal VN383_in5 : std_logic_vector(1 downto 0);
    signal VN384_in0 : std_logic_vector(1 downto 0);
    signal VN384_in1 : std_logic_vector(1 downto 0);
    signal VN384_in2 : std_logic_vector(1 downto 0);
    signal VN384_in3 : std_logic_vector(1 downto 0);
    signal VN384_in4 : std_logic_vector(1 downto 0);
    signal VN384_in5 : std_logic_vector(1 downto 0);
    signal VN385_in0 : std_logic_vector(1 downto 0);
    signal VN385_in1 : std_logic_vector(1 downto 0);
    signal VN385_in2 : std_logic_vector(1 downto 0);
    signal VN385_in3 : std_logic_vector(1 downto 0);
    signal VN385_in4 : std_logic_vector(1 downto 0);
    signal VN385_in5 : std_logic_vector(1 downto 0);
    signal VN386_in0 : std_logic_vector(1 downto 0);
    signal VN386_in1 : std_logic_vector(1 downto 0);
    signal VN386_in2 : std_logic_vector(1 downto 0);
    signal VN386_in3 : std_logic_vector(1 downto 0);
    signal VN386_in4 : std_logic_vector(1 downto 0);
    signal VN386_in5 : std_logic_vector(1 downto 0);
    signal VN387_in0 : std_logic_vector(1 downto 0);
    signal VN387_in1 : std_logic_vector(1 downto 0);
    signal VN387_in2 : std_logic_vector(1 downto 0);
    signal VN387_in3 : std_logic_vector(1 downto 0);
    signal VN387_in4 : std_logic_vector(1 downto 0);
    signal VN387_in5 : std_logic_vector(1 downto 0);
    signal VN388_in0 : std_logic_vector(1 downto 0);
    signal VN388_in1 : std_logic_vector(1 downto 0);
    signal VN388_in2 : std_logic_vector(1 downto 0);
    signal VN388_in3 : std_logic_vector(1 downto 0);
    signal VN388_in4 : std_logic_vector(1 downto 0);
    signal VN388_in5 : std_logic_vector(1 downto 0);
    signal VN389_in0 : std_logic_vector(1 downto 0);
    signal VN389_in1 : std_logic_vector(1 downto 0);
    signal VN389_in2 : std_logic_vector(1 downto 0);
    signal VN389_in3 : std_logic_vector(1 downto 0);
    signal VN389_in4 : std_logic_vector(1 downto 0);
    signal VN389_in5 : std_logic_vector(1 downto 0);
    signal VN390_in0 : std_logic_vector(1 downto 0);
    signal VN390_in1 : std_logic_vector(1 downto 0);
    signal VN390_in2 : std_logic_vector(1 downto 0);
    signal VN390_in3 : std_logic_vector(1 downto 0);
    signal VN390_in4 : std_logic_vector(1 downto 0);
    signal VN390_in5 : std_logic_vector(1 downto 0);
    signal VN391_in0 : std_logic_vector(1 downto 0);
    signal VN391_in1 : std_logic_vector(1 downto 0);
    signal VN391_in2 : std_logic_vector(1 downto 0);
    signal VN391_in3 : std_logic_vector(1 downto 0);
    signal VN391_in4 : std_logic_vector(1 downto 0);
    signal VN391_in5 : std_logic_vector(1 downto 0);
    signal VN392_in0 : std_logic_vector(1 downto 0);
    signal VN392_in1 : std_logic_vector(1 downto 0);
    signal VN392_in2 : std_logic_vector(1 downto 0);
    signal VN392_in3 : std_logic_vector(1 downto 0);
    signal VN392_in4 : std_logic_vector(1 downto 0);
    signal VN392_in5 : std_logic_vector(1 downto 0);
    signal VN393_in0 : std_logic_vector(1 downto 0);
    signal VN393_in1 : std_logic_vector(1 downto 0);
    signal VN393_in2 : std_logic_vector(1 downto 0);
    signal VN393_in3 : std_logic_vector(1 downto 0);
    signal VN393_in4 : std_logic_vector(1 downto 0);
    signal VN393_in5 : std_logic_vector(1 downto 0);
    signal VN394_in0 : std_logic_vector(1 downto 0);
    signal VN394_in1 : std_logic_vector(1 downto 0);
    signal VN394_in2 : std_logic_vector(1 downto 0);
    signal VN394_in3 : std_logic_vector(1 downto 0);
    signal VN394_in4 : std_logic_vector(1 downto 0);
    signal VN394_in5 : std_logic_vector(1 downto 0);
    signal VN395_in0 : std_logic_vector(1 downto 0);
    signal VN395_in1 : std_logic_vector(1 downto 0);
    signal VN395_in2 : std_logic_vector(1 downto 0);
    signal VN395_in3 : std_logic_vector(1 downto 0);
    signal VN395_in4 : std_logic_vector(1 downto 0);
    signal VN395_in5 : std_logic_vector(1 downto 0);
    signal VN396_in0 : std_logic_vector(1 downto 0);
    signal VN396_in1 : std_logic_vector(1 downto 0);
    signal VN396_in2 : std_logic_vector(1 downto 0);
    signal VN396_in3 : std_logic_vector(1 downto 0);
    signal VN396_in4 : std_logic_vector(1 downto 0);
    signal VN396_in5 : std_logic_vector(1 downto 0);
    signal VN397_in0 : std_logic_vector(1 downto 0);
    signal VN397_in1 : std_logic_vector(1 downto 0);
    signal VN397_in2 : std_logic_vector(1 downto 0);
    signal VN397_in3 : std_logic_vector(1 downto 0);
    signal VN397_in4 : std_logic_vector(1 downto 0);
    signal VN397_in5 : std_logic_vector(1 downto 0);
    signal VN398_in0 : std_logic_vector(1 downto 0);
    signal VN398_in1 : std_logic_vector(1 downto 0);
    signal VN398_in2 : std_logic_vector(1 downto 0);
    signal VN398_in3 : std_logic_vector(1 downto 0);
    signal VN398_in4 : std_logic_vector(1 downto 0);
    signal VN398_in5 : std_logic_vector(1 downto 0);
    signal VN399_in0 : std_logic_vector(1 downto 0);
    signal VN399_in1 : std_logic_vector(1 downto 0);
    signal VN399_in2 : std_logic_vector(1 downto 0);
    signal VN399_in3 : std_logic_vector(1 downto 0);
    signal VN399_in4 : std_logic_vector(1 downto 0);
    signal VN399_in5 : std_logic_vector(1 downto 0);
    signal VN400_in0 : std_logic_vector(1 downto 0);
    signal VN400_in1 : std_logic_vector(1 downto 0);
    signal VN400_in2 : std_logic_vector(1 downto 0);
    signal VN400_in3 : std_logic_vector(1 downto 0);
    signal VN400_in4 : std_logic_vector(1 downto 0);
    signal VN400_in5 : std_logic_vector(1 downto 0);
    signal VN401_in0 : std_logic_vector(1 downto 0);
    signal VN401_in1 : std_logic_vector(1 downto 0);
    signal VN401_in2 : std_logic_vector(1 downto 0);
    signal VN401_in3 : std_logic_vector(1 downto 0);
    signal VN401_in4 : std_logic_vector(1 downto 0);
    signal VN401_in5 : std_logic_vector(1 downto 0);
    signal VN402_in0 : std_logic_vector(1 downto 0);
    signal VN402_in1 : std_logic_vector(1 downto 0);
    signal VN402_in2 : std_logic_vector(1 downto 0);
    signal VN402_in3 : std_logic_vector(1 downto 0);
    signal VN402_in4 : std_logic_vector(1 downto 0);
    signal VN402_in5 : std_logic_vector(1 downto 0);
    signal VN403_in0 : std_logic_vector(1 downto 0);
    signal VN403_in1 : std_logic_vector(1 downto 0);
    signal VN403_in2 : std_logic_vector(1 downto 0);
    signal VN403_in3 : std_logic_vector(1 downto 0);
    signal VN403_in4 : std_logic_vector(1 downto 0);
    signal VN403_in5 : std_logic_vector(1 downto 0);
    signal VN404_in0 : std_logic_vector(1 downto 0);
    signal VN404_in1 : std_logic_vector(1 downto 0);
    signal VN404_in2 : std_logic_vector(1 downto 0);
    signal VN404_in3 : std_logic_vector(1 downto 0);
    signal VN404_in4 : std_logic_vector(1 downto 0);
    signal VN404_in5 : std_logic_vector(1 downto 0);
    signal VN405_in0 : std_logic_vector(1 downto 0);
    signal VN405_in1 : std_logic_vector(1 downto 0);
    signal VN405_in2 : std_logic_vector(1 downto 0);
    signal VN405_in3 : std_logic_vector(1 downto 0);
    signal VN405_in4 : std_logic_vector(1 downto 0);
    signal VN405_in5 : std_logic_vector(1 downto 0);
    signal VN406_in0 : std_logic_vector(1 downto 0);
    signal VN406_in1 : std_logic_vector(1 downto 0);
    signal VN406_in2 : std_logic_vector(1 downto 0);
    signal VN406_in3 : std_logic_vector(1 downto 0);
    signal VN406_in4 : std_logic_vector(1 downto 0);
    signal VN406_in5 : std_logic_vector(1 downto 0);
    signal VN407_in0 : std_logic_vector(1 downto 0);
    signal VN407_in1 : std_logic_vector(1 downto 0);
    signal VN407_in2 : std_logic_vector(1 downto 0);
    signal VN407_in3 : std_logic_vector(1 downto 0);
    signal VN407_in4 : std_logic_vector(1 downto 0);
    signal VN407_in5 : std_logic_vector(1 downto 0);
    signal VN408_in0 : std_logic_vector(1 downto 0);
    signal VN408_in1 : std_logic_vector(1 downto 0);
    signal VN408_in2 : std_logic_vector(1 downto 0);
    signal VN408_in3 : std_logic_vector(1 downto 0);
    signal VN408_in4 : std_logic_vector(1 downto 0);
    signal VN408_in5 : std_logic_vector(1 downto 0);
    signal VN409_in0 : std_logic_vector(1 downto 0);
    signal VN409_in1 : std_logic_vector(1 downto 0);
    signal VN409_in2 : std_logic_vector(1 downto 0);
    signal VN409_in3 : std_logic_vector(1 downto 0);
    signal VN409_in4 : std_logic_vector(1 downto 0);
    signal VN409_in5 : std_logic_vector(1 downto 0);
    signal VN410_in0 : std_logic_vector(1 downto 0);
    signal VN410_in1 : std_logic_vector(1 downto 0);
    signal VN410_in2 : std_logic_vector(1 downto 0);
    signal VN410_in3 : std_logic_vector(1 downto 0);
    signal VN410_in4 : std_logic_vector(1 downto 0);
    signal VN410_in5 : std_logic_vector(1 downto 0);
    signal VN411_in0 : std_logic_vector(1 downto 0);
    signal VN411_in1 : std_logic_vector(1 downto 0);
    signal VN411_in2 : std_logic_vector(1 downto 0);
    signal VN411_in3 : std_logic_vector(1 downto 0);
    signal VN411_in4 : std_logic_vector(1 downto 0);
    signal VN411_in5 : std_logic_vector(1 downto 0);
    signal VN412_in0 : std_logic_vector(1 downto 0);
    signal VN412_in1 : std_logic_vector(1 downto 0);
    signal VN412_in2 : std_logic_vector(1 downto 0);
    signal VN412_in3 : std_logic_vector(1 downto 0);
    signal VN412_in4 : std_logic_vector(1 downto 0);
    signal VN412_in5 : std_logic_vector(1 downto 0);
    signal VN413_in0 : std_logic_vector(1 downto 0);
    signal VN413_in1 : std_logic_vector(1 downto 0);
    signal VN413_in2 : std_logic_vector(1 downto 0);
    signal VN413_in3 : std_logic_vector(1 downto 0);
    signal VN413_in4 : std_logic_vector(1 downto 0);
    signal VN413_in5 : std_logic_vector(1 downto 0);
    signal VN414_in0 : std_logic_vector(1 downto 0);
    signal VN414_in1 : std_logic_vector(1 downto 0);
    signal VN414_in2 : std_logic_vector(1 downto 0);
    signal VN414_in3 : std_logic_vector(1 downto 0);
    signal VN414_in4 : std_logic_vector(1 downto 0);
    signal VN414_in5 : std_logic_vector(1 downto 0);
    signal VN415_in0 : std_logic_vector(1 downto 0);
    signal VN415_in1 : std_logic_vector(1 downto 0);
    signal VN415_in2 : std_logic_vector(1 downto 0);
    signal VN415_in3 : std_logic_vector(1 downto 0);
    signal VN415_in4 : std_logic_vector(1 downto 0);
    signal VN415_in5 : std_logic_vector(1 downto 0);
    signal VN416_in0 : std_logic_vector(1 downto 0);
    signal VN416_in1 : std_logic_vector(1 downto 0);
    signal VN416_in2 : std_logic_vector(1 downto 0);
    signal VN416_in3 : std_logic_vector(1 downto 0);
    signal VN416_in4 : std_logic_vector(1 downto 0);
    signal VN416_in5 : std_logic_vector(1 downto 0);
    signal VN417_in0 : std_logic_vector(1 downto 0);
    signal VN417_in1 : std_logic_vector(1 downto 0);
    signal VN417_in2 : std_logic_vector(1 downto 0);
    signal VN417_in3 : std_logic_vector(1 downto 0);
    signal VN417_in4 : std_logic_vector(1 downto 0);
    signal VN417_in5 : std_logic_vector(1 downto 0);
    signal VN418_in0 : std_logic_vector(1 downto 0);
    signal VN418_in1 : std_logic_vector(1 downto 0);
    signal VN418_in2 : std_logic_vector(1 downto 0);
    signal VN418_in3 : std_logic_vector(1 downto 0);
    signal VN418_in4 : std_logic_vector(1 downto 0);
    signal VN418_in5 : std_logic_vector(1 downto 0);
    signal VN419_in0 : std_logic_vector(1 downto 0);
    signal VN419_in1 : std_logic_vector(1 downto 0);
    signal VN419_in2 : std_logic_vector(1 downto 0);
    signal VN419_in3 : std_logic_vector(1 downto 0);
    signal VN419_in4 : std_logic_vector(1 downto 0);
    signal VN419_in5 : std_logic_vector(1 downto 0);
    signal VN420_in0 : std_logic_vector(1 downto 0);
    signal VN420_in1 : std_logic_vector(1 downto 0);
    signal VN420_in2 : std_logic_vector(1 downto 0);
    signal VN420_in3 : std_logic_vector(1 downto 0);
    signal VN420_in4 : std_logic_vector(1 downto 0);
    signal VN420_in5 : std_logic_vector(1 downto 0);
    signal VN421_in0 : std_logic_vector(1 downto 0);
    signal VN421_in1 : std_logic_vector(1 downto 0);
    signal VN421_in2 : std_logic_vector(1 downto 0);
    signal VN421_in3 : std_logic_vector(1 downto 0);
    signal VN421_in4 : std_logic_vector(1 downto 0);
    signal VN421_in5 : std_logic_vector(1 downto 0);
    signal VN422_in0 : std_logic_vector(1 downto 0);
    signal VN422_in1 : std_logic_vector(1 downto 0);
    signal VN422_in2 : std_logic_vector(1 downto 0);
    signal VN422_in3 : std_logic_vector(1 downto 0);
    signal VN422_in4 : std_logic_vector(1 downto 0);
    signal VN422_in5 : std_logic_vector(1 downto 0);
    signal VN423_in0 : std_logic_vector(1 downto 0);
    signal VN423_in1 : std_logic_vector(1 downto 0);
    signal VN423_in2 : std_logic_vector(1 downto 0);
    signal VN423_in3 : std_logic_vector(1 downto 0);
    signal VN423_in4 : std_logic_vector(1 downto 0);
    signal VN423_in5 : std_logic_vector(1 downto 0);
    signal VN424_in0 : std_logic_vector(1 downto 0);
    signal VN424_in1 : std_logic_vector(1 downto 0);
    signal VN424_in2 : std_logic_vector(1 downto 0);
    signal VN424_in3 : std_logic_vector(1 downto 0);
    signal VN424_in4 : std_logic_vector(1 downto 0);
    signal VN424_in5 : std_logic_vector(1 downto 0);
    signal VN425_in0 : std_logic_vector(1 downto 0);
    signal VN425_in1 : std_logic_vector(1 downto 0);
    signal VN425_in2 : std_logic_vector(1 downto 0);
    signal VN425_in3 : std_logic_vector(1 downto 0);
    signal VN425_in4 : std_logic_vector(1 downto 0);
    signal VN425_in5 : std_logic_vector(1 downto 0);
    signal VN426_in0 : std_logic_vector(1 downto 0);
    signal VN426_in1 : std_logic_vector(1 downto 0);
    signal VN426_in2 : std_logic_vector(1 downto 0);
    signal VN426_in3 : std_logic_vector(1 downto 0);
    signal VN426_in4 : std_logic_vector(1 downto 0);
    signal VN426_in5 : std_logic_vector(1 downto 0);
    signal VN427_in0 : std_logic_vector(1 downto 0);
    signal VN427_in1 : std_logic_vector(1 downto 0);
    signal VN427_in2 : std_logic_vector(1 downto 0);
    signal VN427_in3 : std_logic_vector(1 downto 0);
    signal VN427_in4 : std_logic_vector(1 downto 0);
    signal VN427_in5 : std_logic_vector(1 downto 0);
    signal VN428_in0 : std_logic_vector(1 downto 0);
    signal VN428_in1 : std_logic_vector(1 downto 0);
    signal VN428_in2 : std_logic_vector(1 downto 0);
    signal VN428_in3 : std_logic_vector(1 downto 0);
    signal VN428_in4 : std_logic_vector(1 downto 0);
    signal VN428_in5 : std_logic_vector(1 downto 0);
    signal VN429_in0 : std_logic_vector(1 downto 0);
    signal VN429_in1 : std_logic_vector(1 downto 0);
    signal VN429_in2 : std_logic_vector(1 downto 0);
    signal VN429_in3 : std_logic_vector(1 downto 0);
    signal VN429_in4 : std_logic_vector(1 downto 0);
    signal VN429_in5 : std_logic_vector(1 downto 0);
    signal VN430_in0 : std_logic_vector(1 downto 0);
    signal VN430_in1 : std_logic_vector(1 downto 0);
    signal VN430_in2 : std_logic_vector(1 downto 0);
    signal VN430_in3 : std_logic_vector(1 downto 0);
    signal VN430_in4 : std_logic_vector(1 downto 0);
    signal VN430_in5 : std_logic_vector(1 downto 0);
    signal VN431_in0 : std_logic_vector(1 downto 0);
    signal VN431_in1 : std_logic_vector(1 downto 0);
    signal VN431_in2 : std_logic_vector(1 downto 0);
    signal VN431_in3 : std_logic_vector(1 downto 0);
    signal VN431_in4 : std_logic_vector(1 downto 0);
    signal VN431_in5 : std_logic_vector(1 downto 0);
    signal VN432_in0 : std_logic_vector(1 downto 0);
    signal VN432_in1 : std_logic_vector(1 downto 0);
    signal VN432_in2 : std_logic_vector(1 downto 0);
    signal VN432_in3 : std_logic_vector(1 downto 0);
    signal VN432_in4 : std_logic_vector(1 downto 0);
    signal VN432_in5 : std_logic_vector(1 downto 0);
    signal VN433_in0 : std_logic_vector(1 downto 0);
    signal VN433_in1 : std_logic_vector(1 downto 0);
    signal VN433_in2 : std_logic_vector(1 downto 0);
    signal VN433_in3 : std_logic_vector(1 downto 0);
    signal VN433_in4 : std_logic_vector(1 downto 0);
    signal VN433_in5 : std_logic_vector(1 downto 0);
    signal VN434_in0 : std_logic_vector(1 downto 0);
    signal VN434_in1 : std_logic_vector(1 downto 0);
    signal VN434_in2 : std_logic_vector(1 downto 0);
    signal VN434_in3 : std_logic_vector(1 downto 0);
    signal VN434_in4 : std_logic_vector(1 downto 0);
    signal VN434_in5 : std_logic_vector(1 downto 0);
    signal VN435_in0 : std_logic_vector(1 downto 0);
    signal VN435_in1 : std_logic_vector(1 downto 0);
    signal VN435_in2 : std_logic_vector(1 downto 0);
    signal VN435_in3 : std_logic_vector(1 downto 0);
    signal VN435_in4 : std_logic_vector(1 downto 0);
    signal VN435_in5 : std_logic_vector(1 downto 0);
    signal VN436_in0 : std_logic_vector(1 downto 0);
    signal VN436_in1 : std_logic_vector(1 downto 0);
    signal VN436_in2 : std_logic_vector(1 downto 0);
    signal VN436_in3 : std_logic_vector(1 downto 0);
    signal VN436_in4 : std_logic_vector(1 downto 0);
    signal VN436_in5 : std_logic_vector(1 downto 0);
    signal VN437_in0 : std_logic_vector(1 downto 0);
    signal VN437_in1 : std_logic_vector(1 downto 0);
    signal VN437_in2 : std_logic_vector(1 downto 0);
    signal VN437_in3 : std_logic_vector(1 downto 0);
    signal VN437_in4 : std_logic_vector(1 downto 0);
    signal VN437_in5 : std_logic_vector(1 downto 0);
    signal VN438_in0 : std_logic_vector(1 downto 0);
    signal VN438_in1 : std_logic_vector(1 downto 0);
    signal VN438_in2 : std_logic_vector(1 downto 0);
    signal VN438_in3 : std_logic_vector(1 downto 0);
    signal VN438_in4 : std_logic_vector(1 downto 0);
    signal VN438_in5 : std_logic_vector(1 downto 0);
    signal VN439_in0 : std_logic_vector(1 downto 0);
    signal VN439_in1 : std_logic_vector(1 downto 0);
    signal VN439_in2 : std_logic_vector(1 downto 0);
    signal VN439_in3 : std_logic_vector(1 downto 0);
    signal VN439_in4 : std_logic_vector(1 downto 0);
    signal VN439_in5 : std_logic_vector(1 downto 0);
    signal VN440_in0 : std_logic_vector(1 downto 0);
    signal VN440_in1 : std_logic_vector(1 downto 0);
    signal VN440_in2 : std_logic_vector(1 downto 0);
    signal VN440_in3 : std_logic_vector(1 downto 0);
    signal VN440_in4 : std_logic_vector(1 downto 0);
    signal VN440_in5 : std_logic_vector(1 downto 0);
    signal VN441_in0 : std_logic_vector(1 downto 0);
    signal VN441_in1 : std_logic_vector(1 downto 0);
    signal VN441_in2 : std_logic_vector(1 downto 0);
    signal VN441_in3 : std_logic_vector(1 downto 0);
    signal VN441_in4 : std_logic_vector(1 downto 0);
    signal VN441_in5 : std_logic_vector(1 downto 0);
    signal VN442_in0 : std_logic_vector(1 downto 0);
    signal VN442_in1 : std_logic_vector(1 downto 0);
    signal VN442_in2 : std_logic_vector(1 downto 0);
    signal VN442_in3 : std_logic_vector(1 downto 0);
    signal VN442_in4 : std_logic_vector(1 downto 0);
    signal VN442_in5 : std_logic_vector(1 downto 0);
    signal VN443_in0 : std_logic_vector(1 downto 0);
    signal VN443_in1 : std_logic_vector(1 downto 0);
    signal VN443_in2 : std_logic_vector(1 downto 0);
    signal VN443_in3 : std_logic_vector(1 downto 0);
    signal VN443_in4 : std_logic_vector(1 downto 0);
    signal VN443_in5 : std_logic_vector(1 downto 0);
    signal VN444_in0 : std_logic_vector(1 downto 0);
    signal VN444_in1 : std_logic_vector(1 downto 0);
    signal VN444_in2 : std_logic_vector(1 downto 0);
    signal VN444_in3 : std_logic_vector(1 downto 0);
    signal VN444_in4 : std_logic_vector(1 downto 0);
    signal VN444_in5 : std_logic_vector(1 downto 0);
    signal VN445_in0 : std_logic_vector(1 downto 0);
    signal VN445_in1 : std_logic_vector(1 downto 0);
    signal VN445_in2 : std_logic_vector(1 downto 0);
    signal VN445_in3 : std_logic_vector(1 downto 0);
    signal VN445_in4 : std_logic_vector(1 downto 0);
    signal VN445_in5 : std_logic_vector(1 downto 0);
    signal VN446_in0 : std_logic_vector(1 downto 0);
    signal VN446_in1 : std_logic_vector(1 downto 0);
    signal VN446_in2 : std_logic_vector(1 downto 0);
    signal VN446_in3 : std_logic_vector(1 downto 0);
    signal VN446_in4 : std_logic_vector(1 downto 0);
    signal VN446_in5 : std_logic_vector(1 downto 0);
    signal VN447_in0 : std_logic_vector(1 downto 0);
    signal VN447_in1 : std_logic_vector(1 downto 0);
    signal VN447_in2 : std_logic_vector(1 downto 0);
    signal VN447_in3 : std_logic_vector(1 downto 0);
    signal VN447_in4 : std_logic_vector(1 downto 0);
    signal VN447_in5 : std_logic_vector(1 downto 0);
    signal VN448_in0 : std_logic_vector(1 downto 0);
    signal VN448_in1 : std_logic_vector(1 downto 0);
    signal VN448_in2 : std_logic_vector(1 downto 0);
    signal VN448_in3 : std_logic_vector(1 downto 0);
    signal VN448_in4 : std_logic_vector(1 downto 0);
    signal VN448_in5 : std_logic_vector(1 downto 0);
    signal VN449_in0 : std_logic_vector(1 downto 0);
    signal VN449_in1 : std_logic_vector(1 downto 0);
    signal VN449_in2 : std_logic_vector(1 downto 0);
    signal VN449_in3 : std_logic_vector(1 downto 0);
    signal VN449_in4 : std_logic_vector(1 downto 0);
    signal VN449_in5 : std_logic_vector(1 downto 0);
    signal VN450_in0 : std_logic_vector(1 downto 0);
    signal VN450_in1 : std_logic_vector(1 downto 0);
    signal VN450_in2 : std_logic_vector(1 downto 0);
    signal VN450_in3 : std_logic_vector(1 downto 0);
    signal VN450_in4 : std_logic_vector(1 downto 0);
    signal VN450_in5 : std_logic_vector(1 downto 0);
    signal VN451_in0 : std_logic_vector(1 downto 0);
    signal VN451_in1 : std_logic_vector(1 downto 0);
    signal VN451_in2 : std_logic_vector(1 downto 0);
    signal VN451_in3 : std_logic_vector(1 downto 0);
    signal VN451_in4 : std_logic_vector(1 downto 0);
    signal VN451_in5 : std_logic_vector(1 downto 0);
    signal VN452_in0 : std_logic_vector(1 downto 0);
    signal VN452_in1 : std_logic_vector(1 downto 0);
    signal VN452_in2 : std_logic_vector(1 downto 0);
    signal VN452_in3 : std_logic_vector(1 downto 0);
    signal VN452_in4 : std_logic_vector(1 downto 0);
    signal VN452_in5 : std_logic_vector(1 downto 0);
    signal VN453_in0 : std_logic_vector(1 downto 0);
    signal VN453_in1 : std_logic_vector(1 downto 0);
    signal VN453_in2 : std_logic_vector(1 downto 0);
    signal VN453_in3 : std_logic_vector(1 downto 0);
    signal VN453_in4 : std_logic_vector(1 downto 0);
    signal VN453_in5 : std_logic_vector(1 downto 0);
    signal VN454_in0 : std_logic_vector(1 downto 0);
    signal VN454_in1 : std_logic_vector(1 downto 0);
    signal VN454_in2 : std_logic_vector(1 downto 0);
    signal VN454_in3 : std_logic_vector(1 downto 0);
    signal VN454_in4 : std_logic_vector(1 downto 0);
    signal VN454_in5 : std_logic_vector(1 downto 0);
    signal VN455_in0 : std_logic_vector(1 downto 0);
    signal VN455_in1 : std_logic_vector(1 downto 0);
    signal VN455_in2 : std_logic_vector(1 downto 0);
    signal VN455_in3 : std_logic_vector(1 downto 0);
    signal VN455_in4 : std_logic_vector(1 downto 0);
    signal VN455_in5 : std_logic_vector(1 downto 0);
    signal VN456_in0 : std_logic_vector(1 downto 0);
    signal VN456_in1 : std_logic_vector(1 downto 0);
    signal VN456_in2 : std_logic_vector(1 downto 0);
    signal VN456_in3 : std_logic_vector(1 downto 0);
    signal VN456_in4 : std_logic_vector(1 downto 0);
    signal VN456_in5 : std_logic_vector(1 downto 0);
    signal VN457_in0 : std_logic_vector(1 downto 0);
    signal VN457_in1 : std_logic_vector(1 downto 0);
    signal VN457_in2 : std_logic_vector(1 downto 0);
    signal VN457_in3 : std_logic_vector(1 downto 0);
    signal VN457_in4 : std_logic_vector(1 downto 0);
    signal VN457_in5 : std_logic_vector(1 downto 0);
    signal VN458_in0 : std_logic_vector(1 downto 0);
    signal VN458_in1 : std_logic_vector(1 downto 0);
    signal VN458_in2 : std_logic_vector(1 downto 0);
    signal VN458_in3 : std_logic_vector(1 downto 0);
    signal VN458_in4 : std_logic_vector(1 downto 0);
    signal VN458_in5 : std_logic_vector(1 downto 0);
    signal VN459_in0 : std_logic_vector(1 downto 0);
    signal VN459_in1 : std_logic_vector(1 downto 0);
    signal VN459_in2 : std_logic_vector(1 downto 0);
    signal VN459_in3 : std_logic_vector(1 downto 0);
    signal VN459_in4 : std_logic_vector(1 downto 0);
    signal VN459_in5 : std_logic_vector(1 downto 0);
    signal VN460_in0 : std_logic_vector(1 downto 0);
    signal VN460_in1 : std_logic_vector(1 downto 0);
    signal VN460_in2 : std_logic_vector(1 downto 0);
    signal VN460_in3 : std_logic_vector(1 downto 0);
    signal VN460_in4 : std_logic_vector(1 downto 0);
    signal VN460_in5 : std_logic_vector(1 downto 0);
    signal VN461_in0 : std_logic_vector(1 downto 0);
    signal VN461_in1 : std_logic_vector(1 downto 0);
    signal VN461_in2 : std_logic_vector(1 downto 0);
    signal VN461_in3 : std_logic_vector(1 downto 0);
    signal VN461_in4 : std_logic_vector(1 downto 0);
    signal VN461_in5 : std_logic_vector(1 downto 0);
    signal VN462_in0 : std_logic_vector(1 downto 0);
    signal VN462_in1 : std_logic_vector(1 downto 0);
    signal VN462_in2 : std_logic_vector(1 downto 0);
    signal VN462_in3 : std_logic_vector(1 downto 0);
    signal VN462_in4 : std_logic_vector(1 downto 0);
    signal VN462_in5 : std_logic_vector(1 downto 0);
    signal VN463_in0 : std_logic_vector(1 downto 0);
    signal VN463_in1 : std_logic_vector(1 downto 0);
    signal VN463_in2 : std_logic_vector(1 downto 0);
    signal VN463_in3 : std_logic_vector(1 downto 0);
    signal VN463_in4 : std_logic_vector(1 downto 0);
    signal VN463_in5 : std_logic_vector(1 downto 0);
    signal VN464_in0 : std_logic_vector(1 downto 0);
    signal VN464_in1 : std_logic_vector(1 downto 0);
    signal VN464_in2 : std_logic_vector(1 downto 0);
    signal VN464_in3 : std_logic_vector(1 downto 0);
    signal VN464_in4 : std_logic_vector(1 downto 0);
    signal VN464_in5 : std_logic_vector(1 downto 0);
    signal VN465_in0 : std_logic_vector(1 downto 0);
    signal VN465_in1 : std_logic_vector(1 downto 0);
    signal VN465_in2 : std_logic_vector(1 downto 0);
    signal VN465_in3 : std_logic_vector(1 downto 0);
    signal VN465_in4 : std_logic_vector(1 downto 0);
    signal VN465_in5 : std_logic_vector(1 downto 0);
    signal VN466_in0 : std_logic_vector(1 downto 0);
    signal VN466_in1 : std_logic_vector(1 downto 0);
    signal VN466_in2 : std_logic_vector(1 downto 0);
    signal VN466_in3 : std_logic_vector(1 downto 0);
    signal VN466_in4 : std_logic_vector(1 downto 0);
    signal VN466_in5 : std_logic_vector(1 downto 0);
    signal VN467_in0 : std_logic_vector(1 downto 0);
    signal VN467_in1 : std_logic_vector(1 downto 0);
    signal VN467_in2 : std_logic_vector(1 downto 0);
    signal VN467_in3 : std_logic_vector(1 downto 0);
    signal VN467_in4 : std_logic_vector(1 downto 0);
    signal VN467_in5 : std_logic_vector(1 downto 0);
    signal VN468_in0 : std_logic_vector(1 downto 0);
    signal VN468_in1 : std_logic_vector(1 downto 0);
    signal VN468_in2 : std_logic_vector(1 downto 0);
    signal VN468_in3 : std_logic_vector(1 downto 0);
    signal VN468_in4 : std_logic_vector(1 downto 0);
    signal VN468_in5 : std_logic_vector(1 downto 0);
    signal VN469_in0 : std_logic_vector(1 downto 0);
    signal VN469_in1 : std_logic_vector(1 downto 0);
    signal VN469_in2 : std_logic_vector(1 downto 0);
    signal VN469_in3 : std_logic_vector(1 downto 0);
    signal VN469_in4 : std_logic_vector(1 downto 0);
    signal VN469_in5 : std_logic_vector(1 downto 0);
    signal VN470_in0 : std_logic_vector(1 downto 0);
    signal VN470_in1 : std_logic_vector(1 downto 0);
    signal VN470_in2 : std_logic_vector(1 downto 0);
    signal VN470_in3 : std_logic_vector(1 downto 0);
    signal VN470_in4 : std_logic_vector(1 downto 0);
    signal VN470_in5 : std_logic_vector(1 downto 0);
    signal VN471_in0 : std_logic_vector(1 downto 0);
    signal VN471_in1 : std_logic_vector(1 downto 0);
    signal VN471_in2 : std_logic_vector(1 downto 0);
    signal VN471_in3 : std_logic_vector(1 downto 0);
    signal VN471_in4 : std_logic_vector(1 downto 0);
    signal VN471_in5 : std_logic_vector(1 downto 0);
    signal VN472_in0 : std_logic_vector(1 downto 0);
    signal VN472_in1 : std_logic_vector(1 downto 0);
    signal VN472_in2 : std_logic_vector(1 downto 0);
    signal VN472_in3 : std_logic_vector(1 downto 0);
    signal VN472_in4 : std_logic_vector(1 downto 0);
    signal VN472_in5 : std_logic_vector(1 downto 0);
    signal VN473_in0 : std_logic_vector(1 downto 0);
    signal VN473_in1 : std_logic_vector(1 downto 0);
    signal VN473_in2 : std_logic_vector(1 downto 0);
    signal VN473_in3 : std_logic_vector(1 downto 0);
    signal VN473_in4 : std_logic_vector(1 downto 0);
    signal VN473_in5 : std_logic_vector(1 downto 0);
    signal VN474_in0 : std_logic_vector(1 downto 0);
    signal VN474_in1 : std_logic_vector(1 downto 0);
    signal VN474_in2 : std_logic_vector(1 downto 0);
    signal VN474_in3 : std_logic_vector(1 downto 0);
    signal VN474_in4 : std_logic_vector(1 downto 0);
    signal VN474_in5 : std_logic_vector(1 downto 0);
    signal VN475_in0 : std_logic_vector(1 downto 0);
    signal VN475_in1 : std_logic_vector(1 downto 0);
    signal VN475_in2 : std_logic_vector(1 downto 0);
    signal VN475_in3 : std_logic_vector(1 downto 0);
    signal VN475_in4 : std_logic_vector(1 downto 0);
    signal VN475_in5 : std_logic_vector(1 downto 0);
    signal VN476_in0 : std_logic_vector(1 downto 0);
    signal VN476_in1 : std_logic_vector(1 downto 0);
    signal VN476_in2 : std_logic_vector(1 downto 0);
    signal VN476_in3 : std_logic_vector(1 downto 0);
    signal VN476_in4 : std_logic_vector(1 downto 0);
    signal VN476_in5 : std_logic_vector(1 downto 0);
    signal VN477_in0 : std_logic_vector(1 downto 0);
    signal VN477_in1 : std_logic_vector(1 downto 0);
    signal VN477_in2 : std_logic_vector(1 downto 0);
    signal VN477_in3 : std_logic_vector(1 downto 0);
    signal VN477_in4 : std_logic_vector(1 downto 0);
    signal VN477_in5 : std_logic_vector(1 downto 0);
    signal VN478_in0 : std_logic_vector(1 downto 0);
    signal VN478_in1 : std_logic_vector(1 downto 0);
    signal VN478_in2 : std_logic_vector(1 downto 0);
    signal VN478_in3 : std_logic_vector(1 downto 0);
    signal VN478_in4 : std_logic_vector(1 downto 0);
    signal VN478_in5 : std_logic_vector(1 downto 0);
    signal VN479_in0 : std_logic_vector(1 downto 0);
    signal VN479_in1 : std_logic_vector(1 downto 0);
    signal VN479_in2 : std_logic_vector(1 downto 0);
    signal VN479_in3 : std_logic_vector(1 downto 0);
    signal VN479_in4 : std_logic_vector(1 downto 0);
    signal VN479_in5 : std_logic_vector(1 downto 0);
    signal VN480_in0 : std_logic_vector(1 downto 0);
    signal VN480_in1 : std_logic_vector(1 downto 0);
    signal VN480_in2 : std_logic_vector(1 downto 0);
    signal VN480_in3 : std_logic_vector(1 downto 0);
    signal VN480_in4 : std_logic_vector(1 downto 0);
    signal VN480_in5 : std_logic_vector(1 downto 0);
    signal VN481_in0 : std_logic_vector(1 downto 0);
    signal VN481_in1 : std_logic_vector(1 downto 0);
    signal VN481_in2 : std_logic_vector(1 downto 0);
    signal VN481_in3 : std_logic_vector(1 downto 0);
    signal VN481_in4 : std_logic_vector(1 downto 0);
    signal VN481_in5 : std_logic_vector(1 downto 0);
    signal VN482_in0 : std_logic_vector(1 downto 0);
    signal VN482_in1 : std_logic_vector(1 downto 0);
    signal VN482_in2 : std_logic_vector(1 downto 0);
    signal VN482_in3 : std_logic_vector(1 downto 0);
    signal VN482_in4 : std_logic_vector(1 downto 0);
    signal VN482_in5 : std_logic_vector(1 downto 0);
    signal VN483_in0 : std_logic_vector(1 downto 0);
    signal VN483_in1 : std_logic_vector(1 downto 0);
    signal VN483_in2 : std_logic_vector(1 downto 0);
    signal VN483_in3 : std_logic_vector(1 downto 0);
    signal VN483_in4 : std_logic_vector(1 downto 0);
    signal VN483_in5 : std_logic_vector(1 downto 0);
    signal VN484_in0 : std_logic_vector(1 downto 0);
    signal VN484_in1 : std_logic_vector(1 downto 0);
    signal VN484_in2 : std_logic_vector(1 downto 0);
    signal VN484_in3 : std_logic_vector(1 downto 0);
    signal VN484_in4 : std_logic_vector(1 downto 0);
    signal VN484_in5 : std_logic_vector(1 downto 0);
    signal VN485_in0 : std_logic_vector(1 downto 0);
    signal VN485_in1 : std_logic_vector(1 downto 0);
    signal VN485_in2 : std_logic_vector(1 downto 0);
    signal VN485_in3 : std_logic_vector(1 downto 0);
    signal VN485_in4 : std_logic_vector(1 downto 0);
    signal VN485_in5 : std_logic_vector(1 downto 0);
    signal VN486_in0 : std_logic_vector(1 downto 0);
    signal VN486_in1 : std_logic_vector(1 downto 0);
    signal VN486_in2 : std_logic_vector(1 downto 0);
    signal VN486_in3 : std_logic_vector(1 downto 0);
    signal VN486_in4 : std_logic_vector(1 downto 0);
    signal VN486_in5 : std_logic_vector(1 downto 0);
    signal VN487_in0 : std_logic_vector(1 downto 0);
    signal VN487_in1 : std_logic_vector(1 downto 0);
    signal VN487_in2 : std_logic_vector(1 downto 0);
    signal VN487_in3 : std_logic_vector(1 downto 0);
    signal VN487_in4 : std_logic_vector(1 downto 0);
    signal VN487_in5 : std_logic_vector(1 downto 0);
    signal VN488_in0 : std_logic_vector(1 downto 0);
    signal VN488_in1 : std_logic_vector(1 downto 0);
    signal VN488_in2 : std_logic_vector(1 downto 0);
    signal VN488_in3 : std_logic_vector(1 downto 0);
    signal VN488_in4 : std_logic_vector(1 downto 0);
    signal VN488_in5 : std_logic_vector(1 downto 0);
    signal VN489_in0 : std_logic_vector(1 downto 0);
    signal VN489_in1 : std_logic_vector(1 downto 0);
    signal VN489_in2 : std_logic_vector(1 downto 0);
    signal VN489_in3 : std_logic_vector(1 downto 0);
    signal VN489_in4 : std_logic_vector(1 downto 0);
    signal VN489_in5 : std_logic_vector(1 downto 0);
    signal VN490_in0 : std_logic_vector(1 downto 0);
    signal VN490_in1 : std_logic_vector(1 downto 0);
    signal VN490_in2 : std_logic_vector(1 downto 0);
    signal VN490_in3 : std_logic_vector(1 downto 0);
    signal VN490_in4 : std_logic_vector(1 downto 0);
    signal VN490_in5 : std_logic_vector(1 downto 0);
    signal VN491_in0 : std_logic_vector(1 downto 0);
    signal VN491_in1 : std_logic_vector(1 downto 0);
    signal VN491_in2 : std_logic_vector(1 downto 0);
    signal VN491_in3 : std_logic_vector(1 downto 0);
    signal VN491_in4 : std_logic_vector(1 downto 0);
    signal VN491_in5 : std_logic_vector(1 downto 0);
    signal VN492_in0 : std_logic_vector(1 downto 0);
    signal VN492_in1 : std_logic_vector(1 downto 0);
    signal VN492_in2 : std_logic_vector(1 downto 0);
    signal VN492_in3 : std_logic_vector(1 downto 0);
    signal VN492_in4 : std_logic_vector(1 downto 0);
    signal VN492_in5 : std_logic_vector(1 downto 0);
    signal VN493_in0 : std_logic_vector(1 downto 0);
    signal VN493_in1 : std_logic_vector(1 downto 0);
    signal VN493_in2 : std_logic_vector(1 downto 0);
    signal VN493_in3 : std_logic_vector(1 downto 0);
    signal VN493_in4 : std_logic_vector(1 downto 0);
    signal VN493_in5 : std_logic_vector(1 downto 0);
    signal VN494_in0 : std_logic_vector(1 downto 0);
    signal VN494_in1 : std_logic_vector(1 downto 0);
    signal VN494_in2 : std_logic_vector(1 downto 0);
    signal VN494_in3 : std_logic_vector(1 downto 0);
    signal VN494_in4 : std_logic_vector(1 downto 0);
    signal VN494_in5 : std_logic_vector(1 downto 0);
    signal VN495_in0 : std_logic_vector(1 downto 0);
    signal VN495_in1 : std_logic_vector(1 downto 0);
    signal VN495_in2 : std_logic_vector(1 downto 0);
    signal VN495_in3 : std_logic_vector(1 downto 0);
    signal VN495_in4 : std_logic_vector(1 downto 0);
    signal VN495_in5 : std_logic_vector(1 downto 0);
    signal VN496_in0 : std_logic_vector(1 downto 0);
    signal VN496_in1 : std_logic_vector(1 downto 0);
    signal VN496_in2 : std_logic_vector(1 downto 0);
    signal VN496_in3 : std_logic_vector(1 downto 0);
    signal VN496_in4 : std_logic_vector(1 downto 0);
    signal VN496_in5 : std_logic_vector(1 downto 0);
    signal VN497_in0 : std_logic_vector(1 downto 0);
    signal VN497_in1 : std_logic_vector(1 downto 0);
    signal VN497_in2 : std_logic_vector(1 downto 0);
    signal VN497_in3 : std_logic_vector(1 downto 0);
    signal VN497_in4 : std_logic_vector(1 downto 0);
    signal VN497_in5 : std_logic_vector(1 downto 0);
    signal VN498_in0 : std_logic_vector(1 downto 0);
    signal VN498_in1 : std_logic_vector(1 downto 0);
    signal VN498_in2 : std_logic_vector(1 downto 0);
    signal VN498_in3 : std_logic_vector(1 downto 0);
    signal VN498_in4 : std_logic_vector(1 downto 0);
    signal VN498_in5 : std_logic_vector(1 downto 0);
    signal VN499_in0 : std_logic_vector(1 downto 0);
    signal VN499_in1 : std_logic_vector(1 downto 0);
    signal VN499_in2 : std_logic_vector(1 downto 0);
    signal VN499_in3 : std_logic_vector(1 downto 0);
    signal VN499_in4 : std_logic_vector(1 downto 0);
    signal VN499_in5 : std_logic_vector(1 downto 0);
    signal VN500_in0 : std_logic_vector(1 downto 0);
    signal VN500_in1 : std_logic_vector(1 downto 0);
    signal VN500_in2 : std_logic_vector(1 downto 0);
    signal VN500_in3 : std_logic_vector(1 downto 0);
    signal VN500_in4 : std_logic_vector(1 downto 0);
    signal VN500_in5 : std_logic_vector(1 downto 0);
    signal VN501_in0 : std_logic_vector(1 downto 0);
    signal VN501_in1 : std_logic_vector(1 downto 0);
    signal VN501_in2 : std_logic_vector(1 downto 0);
    signal VN501_in3 : std_logic_vector(1 downto 0);
    signal VN501_in4 : std_logic_vector(1 downto 0);
    signal VN501_in5 : std_logic_vector(1 downto 0);
    signal VN502_in0 : std_logic_vector(1 downto 0);
    signal VN502_in1 : std_logic_vector(1 downto 0);
    signal VN502_in2 : std_logic_vector(1 downto 0);
    signal VN502_in3 : std_logic_vector(1 downto 0);
    signal VN502_in4 : std_logic_vector(1 downto 0);
    signal VN502_in5 : std_logic_vector(1 downto 0);
    signal VN503_in0 : std_logic_vector(1 downto 0);
    signal VN503_in1 : std_logic_vector(1 downto 0);
    signal VN503_in2 : std_logic_vector(1 downto 0);
    signal VN503_in3 : std_logic_vector(1 downto 0);
    signal VN503_in4 : std_logic_vector(1 downto 0);
    signal VN503_in5 : std_logic_vector(1 downto 0);
    signal VN504_in0 : std_logic_vector(1 downto 0);
    signal VN504_in1 : std_logic_vector(1 downto 0);
    signal VN504_in2 : std_logic_vector(1 downto 0);
    signal VN504_in3 : std_logic_vector(1 downto 0);
    signal VN504_in4 : std_logic_vector(1 downto 0);
    signal VN504_in5 : std_logic_vector(1 downto 0);
    signal VN505_in0 : std_logic_vector(1 downto 0);
    signal VN505_in1 : std_logic_vector(1 downto 0);
    signal VN505_in2 : std_logic_vector(1 downto 0);
    signal VN505_in3 : std_logic_vector(1 downto 0);
    signal VN505_in4 : std_logic_vector(1 downto 0);
    signal VN505_in5 : std_logic_vector(1 downto 0);
    signal VN506_in0 : std_logic_vector(1 downto 0);
    signal VN506_in1 : std_logic_vector(1 downto 0);
    signal VN506_in2 : std_logic_vector(1 downto 0);
    signal VN506_in3 : std_logic_vector(1 downto 0);
    signal VN506_in4 : std_logic_vector(1 downto 0);
    signal VN506_in5 : std_logic_vector(1 downto 0);
    signal VN507_in0 : std_logic_vector(1 downto 0);
    signal VN507_in1 : std_logic_vector(1 downto 0);
    signal VN507_in2 : std_logic_vector(1 downto 0);
    signal VN507_in3 : std_logic_vector(1 downto 0);
    signal VN507_in4 : std_logic_vector(1 downto 0);
    signal VN507_in5 : std_logic_vector(1 downto 0);
    signal VN508_in0 : std_logic_vector(1 downto 0);
    signal VN508_in1 : std_logic_vector(1 downto 0);
    signal VN508_in2 : std_logic_vector(1 downto 0);
    signal VN508_in3 : std_logic_vector(1 downto 0);
    signal VN508_in4 : std_logic_vector(1 downto 0);
    signal VN508_in5 : std_logic_vector(1 downto 0);
    signal VN509_in0 : std_logic_vector(1 downto 0);
    signal VN509_in1 : std_logic_vector(1 downto 0);
    signal VN509_in2 : std_logic_vector(1 downto 0);
    signal VN509_in3 : std_logic_vector(1 downto 0);
    signal VN509_in4 : std_logic_vector(1 downto 0);
    signal VN509_in5 : std_logic_vector(1 downto 0);
    signal VN510_in0 : std_logic_vector(1 downto 0);
    signal VN510_in1 : std_logic_vector(1 downto 0);
    signal VN510_in2 : std_logic_vector(1 downto 0);
    signal VN510_in3 : std_logic_vector(1 downto 0);
    signal VN510_in4 : std_logic_vector(1 downto 0);
    signal VN510_in5 : std_logic_vector(1 downto 0);
    signal VN511_in0 : std_logic_vector(1 downto 0);
    signal VN511_in1 : std_logic_vector(1 downto 0);
    signal VN511_in2 : std_logic_vector(1 downto 0);
    signal VN511_in3 : std_logic_vector(1 downto 0);
    signal VN511_in4 : std_logic_vector(1 downto 0);
    signal VN511_in5 : std_logic_vector(1 downto 0);
    signal VN512_in0 : std_logic_vector(1 downto 0);
    signal VN512_in1 : std_logic_vector(1 downto 0);
    signal VN512_in2 : std_logic_vector(1 downto 0);
    signal VN512_in3 : std_logic_vector(1 downto 0);
    signal VN512_in4 : std_logic_vector(1 downto 0);
    signal VN512_in5 : std_logic_vector(1 downto 0);
    signal VN513_in0 : std_logic_vector(1 downto 0);
    signal VN513_in1 : std_logic_vector(1 downto 0);
    signal VN513_in2 : std_logic_vector(1 downto 0);
    signal VN513_in3 : std_logic_vector(1 downto 0);
    signal VN513_in4 : std_logic_vector(1 downto 0);
    signal VN513_in5 : std_logic_vector(1 downto 0);
    signal VN514_in0 : std_logic_vector(1 downto 0);
    signal VN514_in1 : std_logic_vector(1 downto 0);
    signal VN514_in2 : std_logic_vector(1 downto 0);
    signal VN514_in3 : std_logic_vector(1 downto 0);
    signal VN514_in4 : std_logic_vector(1 downto 0);
    signal VN514_in5 : std_logic_vector(1 downto 0);
    signal VN515_in0 : std_logic_vector(1 downto 0);
    signal VN515_in1 : std_logic_vector(1 downto 0);
    signal VN515_in2 : std_logic_vector(1 downto 0);
    signal VN515_in3 : std_logic_vector(1 downto 0);
    signal VN515_in4 : std_logic_vector(1 downto 0);
    signal VN515_in5 : std_logic_vector(1 downto 0);
    signal VN516_in0 : std_logic_vector(1 downto 0);
    signal VN516_in1 : std_logic_vector(1 downto 0);
    signal VN516_in2 : std_logic_vector(1 downto 0);
    signal VN516_in3 : std_logic_vector(1 downto 0);
    signal VN516_in4 : std_logic_vector(1 downto 0);
    signal VN516_in5 : std_logic_vector(1 downto 0);
    signal VN517_in0 : std_logic_vector(1 downto 0);
    signal VN517_in1 : std_logic_vector(1 downto 0);
    signal VN517_in2 : std_logic_vector(1 downto 0);
    signal VN517_in3 : std_logic_vector(1 downto 0);
    signal VN517_in4 : std_logic_vector(1 downto 0);
    signal VN517_in5 : std_logic_vector(1 downto 0);
    signal VN518_in0 : std_logic_vector(1 downto 0);
    signal VN518_in1 : std_logic_vector(1 downto 0);
    signal VN518_in2 : std_logic_vector(1 downto 0);
    signal VN518_in3 : std_logic_vector(1 downto 0);
    signal VN518_in4 : std_logic_vector(1 downto 0);
    signal VN518_in5 : std_logic_vector(1 downto 0);
    signal VN519_in0 : std_logic_vector(1 downto 0);
    signal VN519_in1 : std_logic_vector(1 downto 0);
    signal VN519_in2 : std_logic_vector(1 downto 0);
    signal VN519_in3 : std_logic_vector(1 downto 0);
    signal VN519_in4 : std_logic_vector(1 downto 0);
    signal VN519_in5 : std_logic_vector(1 downto 0);
    signal VN520_in0 : std_logic_vector(1 downto 0);
    signal VN520_in1 : std_logic_vector(1 downto 0);
    signal VN520_in2 : std_logic_vector(1 downto 0);
    signal VN520_in3 : std_logic_vector(1 downto 0);
    signal VN520_in4 : std_logic_vector(1 downto 0);
    signal VN520_in5 : std_logic_vector(1 downto 0);
    signal VN521_in0 : std_logic_vector(1 downto 0);
    signal VN521_in1 : std_logic_vector(1 downto 0);
    signal VN521_in2 : std_logic_vector(1 downto 0);
    signal VN521_in3 : std_logic_vector(1 downto 0);
    signal VN521_in4 : std_logic_vector(1 downto 0);
    signal VN521_in5 : std_logic_vector(1 downto 0);
    signal VN522_in0 : std_logic_vector(1 downto 0);
    signal VN522_in1 : std_logic_vector(1 downto 0);
    signal VN522_in2 : std_logic_vector(1 downto 0);
    signal VN522_in3 : std_logic_vector(1 downto 0);
    signal VN522_in4 : std_logic_vector(1 downto 0);
    signal VN522_in5 : std_logic_vector(1 downto 0);
    signal VN523_in0 : std_logic_vector(1 downto 0);
    signal VN523_in1 : std_logic_vector(1 downto 0);
    signal VN523_in2 : std_logic_vector(1 downto 0);
    signal VN523_in3 : std_logic_vector(1 downto 0);
    signal VN523_in4 : std_logic_vector(1 downto 0);
    signal VN523_in5 : std_logic_vector(1 downto 0);
    signal VN524_in0 : std_logic_vector(1 downto 0);
    signal VN524_in1 : std_logic_vector(1 downto 0);
    signal VN524_in2 : std_logic_vector(1 downto 0);
    signal VN524_in3 : std_logic_vector(1 downto 0);
    signal VN524_in4 : std_logic_vector(1 downto 0);
    signal VN524_in5 : std_logic_vector(1 downto 0);
    signal VN525_in0 : std_logic_vector(1 downto 0);
    signal VN525_in1 : std_logic_vector(1 downto 0);
    signal VN525_in2 : std_logic_vector(1 downto 0);
    signal VN525_in3 : std_logic_vector(1 downto 0);
    signal VN525_in4 : std_logic_vector(1 downto 0);
    signal VN525_in5 : std_logic_vector(1 downto 0);
    signal VN526_in0 : std_logic_vector(1 downto 0);
    signal VN526_in1 : std_logic_vector(1 downto 0);
    signal VN526_in2 : std_logic_vector(1 downto 0);
    signal VN526_in3 : std_logic_vector(1 downto 0);
    signal VN526_in4 : std_logic_vector(1 downto 0);
    signal VN526_in5 : std_logic_vector(1 downto 0);
    signal VN527_in0 : std_logic_vector(1 downto 0);
    signal VN527_in1 : std_logic_vector(1 downto 0);
    signal VN527_in2 : std_logic_vector(1 downto 0);
    signal VN527_in3 : std_logic_vector(1 downto 0);
    signal VN527_in4 : std_logic_vector(1 downto 0);
    signal VN527_in5 : std_logic_vector(1 downto 0);
    signal VN528_in0 : std_logic_vector(1 downto 0);
    signal VN528_in1 : std_logic_vector(1 downto 0);
    signal VN528_in2 : std_logic_vector(1 downto 0);
    signal VN528_in3 : std_logic_vector(1 downto 0);
    signal VN528_in4 : std_logic_vector(1 downto 0);
    signal VN528_in5 : std_logic_vector(1 downto 0);
    signal VN529_in0 : std_logic_vector(1 downto 0);
    signal VN529_in1 : std_logic_vector(1 downto 0);
    signal VN529_in2 : std_logic_vector(1 downto 0);
    signal VN529_in3 : std_logic_vector(1 downto 0);
    signal VN529_in4 : std_logic_vector(1 downto 0);
    signal VN529_in5 : std_logic_vector(1 downto 0);
    signal VN530_in0 : std_logic_vector(1 downto 0);
    signal VN530_in1 : std_logic_vector(1 downto 0);
    signal VN530_in2 : std_logic_vector(1 downto 0);
    signal VN530_in3 : std_logic_vector(1 downto 0);
    signal VN530_in4 : std_logic_vector(1 downto 0);
    signal VN530_in5 : std_logic_vector(1 downto 0);
    signal VN531_in0 : std_logic_vector(1 downto 0);
    signal VN531_in1 : std_logic_vector(1 downto 0);
    signal VN531_in2 : std_logic_vector(1 downto 0);
    signal VN531_in3 : std_logic_vector(1 downto 0);
    signal VN531_in4 : std_logic_vector(1 downto 0);
    signal VN531_in5 : std_logic_vector(1 downto 0);
    signal VN532_in0 : std_logic_vector(1 downto 0);
    signal VN532_in1 : std_logic_vector(1 downto 0);
    signal VN532_in2 : std_logic_vector(1 downto 0);
    signal VN532_in3 : std_logic_vector(1 downto 0);
    signal VN532_in4 : std_logic_vector(1 downto 0);
    signal VN532_in5 : std_logic_vector(1 downto 0);
    signal VN533_in0 : std_logic_vector(1 downto 0);
    signal VN533_in1 : std_logic_vector(1 downto 0);
    signal VN533_in2 : std_logic_vector(1 downto 0);
    signal VN533_in3 : std_logic_vector(1 downto 0);
    signal VN533_in4 : std_logic_vector(1 downto 0);
    signal VN533_in5 : std_logic_vector(1 downto 0);
    signal VN534_in0 : std_logic_vector(1 downto 0);
    signal VN534_in1 : std_logic_vector(1 downto 0);
    signal VN534_in2 : std_logic_vector(1 downto 0);
    signal VN534_in3 : std_logic_vector(1 downto 0);
    signal VN534_in4 : std_logic_vector(1 downto 0);
    signal VN534_in5 : std_logic_vector(1 downto 0);
    signal VN535_in0 : std_logic_vector(1 downto 0);
    signal VN535_in1 : std_logic_vector(1 downto 0);
    signal VN535_in2 : std_logic_vector(1 downto 0);
    signal VN535_in3 : std_logic_vector(1 downto 0);
    signal VN535_in4 : std_logic_vector(1 downto 0);
    signal VN535_in5 : std_logic_vector(1 downto 0);
    signal VN536_in0 : std_logic_vector(1 downto 0);
    signal VN536_in1 : std_logic_vector(1 downto 0);
    signal VN536_in2 : std_logic_vector(1 downto 0);
    signal VN536_in3 : std_logic_vector(1 downto 0);
    signal VN536_in4 : std_logic_vector(1 downto 0);
    signal VN536_in5 : std_logic_vector(1 downto 0);
    signal VN537_in0 : std_logic_vector(1 downto 0);
    signal VN537_in1 : std_logic_vector(1 downto 0);
    signal VN537_in2 : std_logic_vector(1 downto 0);
    signal VN537_in3 : std_logic_vector(1 downto 0);
    signal VN537_in4 : std_logic_vector(1 downto 0);
    signal VN537_in5 : std_logic_vector(1 downto 0);
    signal VN538_in0 : std_logic_vector(1 downto 0);
    signal VN538_in1 : std_logic_vector(1 downto 0);
    signal VN538_in2 : std_logic_vector(1 downto 0);
    signal VN538_in3 : std_logic_vector(1 downto 0);
    signal VN538_in4 : std_logic_vector(1 downto 0);
    signal VN538_in5 : std_logic_vector(1 downto 0);
    signal VN539_in0 : std_logic_vector(1 downto 0);
    signal VN539_in1 : std_logic_vector(1 downto 0);
    signal VN539_in2 : std_logic_vector(1 downto 0);
    signal VN539_in3 : std_logic_vector(1 downto 0);
    signal VN539_in4 : std_logic_vector(1 downto 0);
    signal VN539_in5 : std_logic_vector(1 downto 0);
    signal VN540_in0 : std_logic_vector(1 downto 0);
    signal VN540_in1 : std_logic_vector(1 downto 0);
    signal VN540_in2 : std_logic_vector(1 downto 0);
    signal VN540_in3 : std_logic_vector(1 downto 0);
    signal VN540_in4 : std_logic_vector(1 downto 0);
    signal VN540_in5 : std_logic_vector(1 downto 0);
    signal VN541_in0 : std_logic_vector(1 downto 0);
    signal VN541_in1 : std_logic_vector(1 downto 0);
    signal VN541_in2 : std_logic_vector(1 downto 0);
    signal VN541_in3 : std_logic_vector(1 downto 0);
    signal VN541_in4 : std_logic_vector(1 downto 0);
    signal VN541_in5 : std_logic_vector(1 downto 0);
    signal VN542_in0 : std_logic_vector(1 downto 0);
    signal VN542_in1 : std_logic_vector(1 downto 0);
    signal VN542_in2 : std_logic_vector(1 downto 0);
    signal VN542_in3 : std_logic_vector(1 downto 0);
    signal VN542_in4 : std_logic_vector(1 downto 0);
    signal VN542_in5 : std_logic_vector(1 downto 0);
    signal VN543_in0 : std_logic_vector(1 downto 0);
    signal VN543_in1 : std_logic_vector(1 downto 0);
    signal VN543_in2 : std_logic_vector(1 downto 0);
    signal VN543_in3 : std_logic_vector(1 downto 0);
    signal VN543_in4 : std_logic_vector(1 downto 0);
    signal VN543_in5 : std_logic_vector(1 downto 0);
    signal VN544_in0 : std_logic_vector(1 downto 0);
    signal VN544_in1 : std_logic_vector(1 downto 0);
    signal VN544_in2 : std_logic_vector(1 downto 0);
    signal VN544_in3 : std_logic_vector(1 downto 0);
    signal VN544_in4 : std_logic_vector(1 downto 0);
    signal VN544_in5 : std_logic_vector(1 downto 0);
    signal VN545_in0 : std_logic_vector(1 downto 0);
    signal VN545_in1 : std_logic_vector(1 downto 0);
    signal VN545_in2 : std_logic_vector(1 downto 0);
    signal VN545_in3 : std_logic_vector(1 downto 0);
    signal VN545_in4 : std_logic_vector(1 downto 0);
    signal VN545_in5 : std_logic_vector(1 downto 0);
    signal VN546_in0 : std_logic_vector(1 downto 0);
    signal VN546_in1 : std_logic_vector(1 downto 0);
    signal VN546_in2 : std_logic_vector(1 downto 0);
    signal VN546_in3 : std_logic_vector(1 downto 0);
    signal VN546_in4 : std_logic_vector(1 downto 0);
    signal VN546_in5 : std_logic_vector(1 downto 0);
    signal VN547_in0 : std_logic_vector(1 downto 0);
    signal VN547_in1 : std_logic_vector(1 downto 0);
    signal VN547_in2 : std_logic_vector(1 downto 0);
    signal VN547_in3 : std_logic_vector(1 downto 0);
    signal VN547_in4 : std_logic_vector(1 downto 0);
    signal VN547_in5 : std_logic_vector(1 downto 0);
    signal VN548_in0 : std_logic_vector(1 downto 0);
    signal VN548_in1 : std_logic_vector(1 downto 0);
    signal VN548_in2 : std_logic_vector(1 downto 0);
    signal VN548_in3 : std_logic_vector(1 downto 0);
    signal VN548_in4 : std_logic_vector(1 downto 0);
    signal VN548_in5 : std_logic_vector(1 downto 0);
    signal VN549_in0 : std_logic_vector(1 downto 0);
    signal VN549_in1 : std_logic_vector(1 downto 0);
    signal VN549_in2 : std_logic_vector(1 downto 0);
    signal VN549_in3 : std_logic_vector(1 downto 0);
    signal VN549_in4 : std_logic_vector(1 downto 0);
    signal VN549_in5 : std_logic_vector(1 downto 0);
    signal VN550_in0 : std_logic_vector(1 downto 0);
    signal VN550_in1 : std_logic_vector(1 downto 0);
    signal VN550_in2 : std_logic_vector(1 downto 0);
    signal VN550_in3 : std_logic_vector(1 downto 0);
    signal VN550_in4 : std_logic_vector(1 downto 0);
    signal VN550_in5 : std_logic_vector(1 downto 0);
    signal VN551_in0 : std_logic_vector(1 downto 0);
    signal VN551_in1 : std_logic_vector(1 downto 0);
    signal VN551_in2 : std_logic_vector(1 downto 0);
    signal VN551_in3 : std_logic_vector(1 downto 0);
    signal VN551_in4 : std_logic_vector(1 downto 0);
    signal VN551_in5 : std_logic_vector(1 downto 0);
    signal VN552_in0 : std_logic_vector(1 downto 0);
    signal VN552_in1 : std_logic_vector(1 downto 0);
    signal VN552_in2 : std_logic_vector(1 downto 0);
    signal VN552_in3 : std_logic_vector(1 downto 0);
    signal VN552_in4 : std_logic_vector(1 downto 0);
    signal VN552_in5 : std_logic_vector(1 downto 0);
    signal VN553_in0 : std_logic_vector(1 downto 0);
    signal VN553_in1 : std_logic_vector(1 downto 0);
    signal VN553_in2 : std_logic_vector(1 downto 0);
    signal VN553_in3 : std_logic_vector(1 downto 0);
    signal VN553_in4 : std_logic_vector(1 downto 0);
    signal VN553_in5 : std_logic_vector(1 downto 0);
    signal VN554_in0 : std_logic_vector(1 downto 0);
    signal VN554_in1 : std_logic_vector(1 downto 0);
    signal VN554_in2 : std_logic_vector(1 downto 0);
    signal VN554_in3 : std_logic_vector(1 downto 0);
    signal VN554_in4 : std_logic_vector(1 downto 0);
    signal VN554_in5 : std_logic_vector(1 downto 0);
    signal VN555_in0 : std_logic_vector(1 downto 0);
    signal VN555_in1 : std_logic_vector(1 downto 0);
    signal VN555_in2 : std_logic_vector(1 downto 0);
    signal VN555_in3 : std_logic_vector(1 downto 0);
    signal VN555_in4 : std_logic_vector(1 downto 0);
    signal VN555_in5 : std_logic_vector(1 downto 0);
    signal VN556_in0 : std_logic_vector(1 downto 0);
    signal VN556_in1 : std_logic_vector(1 downto 0);
    signal VN556_in2 : std_logic_vector(1 downto 0);
    signal VN556_in3 : std_logic_vector(1 downto 0);
    signal VN556_in4 : std_logic_vector(1 downto 0);
    signal VN556_in5 : std_logic_vector(1 downto 0);
    signal VN557_in0 : std_logic_vector(1 downto 0);
    signal VN557_in1 : std_logic_vector(1 downto 0);
    signal VN557_in2 : std_logic_vector(1 downto 0);
    signal VN557_in3 : std_logic_vector(1 downto 0);
    signal VN557_in4 : std_logic_vector(1 downto 0);
    signal VN557_in5 : std_logic_vector(1 downto 0);
    signal VN558_in0 : std_logic_vector(1 downto 0);
    signal VN558_in1 : std_logic_vector(1 downto 0);
    signal VN558_in2 : std_logic_vector(1 downto 0);
    signal VN558_in3 : std_logic_vector(1 downto 0);
    signal VN558_in4 : std_logic_vector(1 downto 0);
    signal VN558_in5 : std_logic_vector(1 downto 0);
    signal VN559_in0 : std_logic_vector(1 downto 0);
    signal VN559_in1 : std_logic_vector(1 downto 0);
    signal VN559_in2 : std_logic_vector(1 downto 0);
    signal VN559_in3 : std_logic_vector(1 downto 0);
    signal VN559_in4 : std_logic_vector(1 downto 0);
    signal VN559_in5 : std_logic_vector(1 downto 0);
    signal VN560_in0 : std_logic_vector(1 downto 0);
    signal VN560_in1 : std_logic_vector(1 downto 0);
    signal VN560_in2 : std_logic_vector(1 downto 0);
    signal VN560_in3 : std_logic_vector(1 downto 0);
    signal VN560_in4 : std_logic_vector(1 downto 0);
    signal VN560_in5 : std_logic_vector(1 downto 0);
    signal VN561_in0 : std_logic_vector(1 downto 0);
    signal VN561_in1 : std_logic_vector(1 downto 0);
    signal VN561_in2 : std_logic_vector(1 downto 0);
    signal VN561_in3 : std_logic_vector(1 downto 0);
    signal VN561_in4 : std_logic_vector(1 downto 0);
    signal VN561_in5 : std_logic_vector(1 downto 0);
    signal VN562_in0 : std_logic_vector(1 downto 0);
    signal VN562_in1 : std_logic_vector(1 downto 0);
    signal VN562_in2 : std_logic_vector(1 downto 0);
    signal VN562_in3 : std_logic_vector(1 downto 0);
    signal VN562_in4 : std_logic_vector(1 downto 0);
    signal VN562_in5 : std_logic_vector(1 downto 0);
    signal VN563_in0 : std_logic_vector(1 downto 0);
    signal VN563_in1 : std_logic_vector(1 downto 0);
    signal VN563_in2 : std_logic_vector(1 downto 0);
    signal VN563_in3 : std_logic_vector(1 downto 0);
    signal VN563_in4 : std_logic_vector(1 downto 0);
    signal VN563_in5 : std_logic_vector(1 downto 0);
    signal VN564_in0 : std_logic_vector(1 downto 0);
    signal VN564_in1 : std_logic_vector(1 downto 0);
    signal VN564_in2 : std_logic_vector(1 downto 0);
    signal VN564_in3 : std_logic_vector(1 downto 0);
    signal VN564_in4 : std_logic_vector(1 downto 0);
    signal VN564_in5 : std_logic_vector(1 downto 0);
    signal VN565_in0 : std_logic_vector(1 downto 0);
    signal VN565_in1 : std_logic_vector(1 downto 0);
    signal VN565_in2 : std_logic_vector(1 downto 0);
    signal VN565_in3 : std_logic_vector(1 downto 0);
    signal VN565_in4 : std_logic_vector(1 downto 0);
    signal VN565_in5 : std_logic_vector(1 downto 0);
    signal VN566_in0 : std_logic_vector(1 downto 0);
    signal VN566_in1 : std_logic_vector(1 downto 0);
    signal VN566_in2 : std_logic_vector(1 downto 0);
    signal VN566_in3 : std_logic_vector(1 downto 0);
    signal VN566_in4 : std_logic_vector(1 downto 0);
    signal VN566_in5 : std_logic_vector(1 downto 0);
    signal VN567_in0 : std_logic_vector(1 downto 0);
    signal VN567_in1 : std_logic_vector(1 downto 0);
    signal VN567_in2 : std_logic_vector(1 downto 0);
    signal VN567_in3 : std_logic_vector(1 downto 0);
    signal VN567_in4 : std_logic_vector(1 downto 0);
    signal VN567_in5 : std_logic_vector(1 downto 0);
    signal VN568_in0 : std_logic_vector(1 downto 0);
    signal VN568_in1 : std_logic_vector(1 downto 0);
    signal VN568_in2 : std_logic_vector(1 downto 0);
    signal VN568_in3 : std_logic_vector(1 downto 0);
    signal VN568_in4 : std_logic_vector(1 downto 0);
    signal VN568_in5 : std_logic_vector(1 downto 0);
    signal VN569_in0 : std_logic_vector(1 downto 0);
    signal VN569_in1 : std_logic_vector(1 downto 0);
    signal VN569_in2 : std_logic_vector(1 downto 0);
    signal VN569_in3 : std_logic_vector(1 downto 0);
    signal VN569_in4 : std_logic_vector(1 downto 0);
    signal VN569_in5 : std_logic_vector(1 downto 0);
    signal VN570_in0 : std_logic_vector(1 downto 0);
    signal VN570_in1 : std_logic_vector(1 downto 0);
    signal VN570_in2 : std_logic_vector(1 downto 0);
    signal VN570_in3 : std_logic_vector(1 downto 0);
    signal VN570_in4 : std_logic_vector(1 downto 0);
    signal VN570_in5 : std_logic_vector(1 downto 0);
    signal VN571_in0 : std_logic_vector(1 downto 0);
    signal VN571_in1 : std_logic_vector(1 downto 0);
    signal VN571_in2 : std_logic_vector(1 downto 0);
    signal VN571_in3 : std_logic_vector(1 downto 0);
    signal VN571_in4 : std_logic_vector(1 downto 0);
    signal VN571_in5 : std_logic_vector(1 downto 0);
    signal VN572_in0 : std_logic_vector(1 downto 0);
    signal VN572_in1 : std_logic_vector(1 downto 0);
    signal VN572_in2 : std_logic_vector(1 downto 0);
    signal VN572_in3 : std_logic_vector(1 downto 0);
    signal VN572_in4 : std_logic_vector(1 downto 0);
    signal VN572_in5 : std_logic_vector(1 downto 0);
    signal VN573_in0 : std_logic_vector(1 downto 0);
    signal VN573_in1 : std_logic_vector(1 downto 0);
    signal VN573_in2 : std_logic_vector(1 downto 0);
    signal VN573_in3 : std_logic_vector(1 downto 0);
    signal VN573_in4 : std_logic_vector(1 downto 0);
    signal VN573_in5 : std_logic_vector(1 downto 0);
    signal VN574_in0 : std_logic_vector(1 downto 0);
    signal VN574_in1 : std_logic_vector(1 downto 0);
    signal VN574_in2 : std_logic_vector(1 downto 0);
    signal VN574_in3 : std_logic_vector(1 downto 0);
    signal VN574_in4 : std_logic_vector(1 downto 0);
    signal VN574_in5 : std_logic_vector(1 downto 0);
    signal VN575_in0 : std_logic_vector(1 downto 0);
    signal VN575_in1 : std_logic_vector(1 downto 0);
    signal VN575_in2 : std_logic_vector(1 downto 0);
    signal VN575_in3 : std_logic_vector(1 downto 0);
    signal VN575_in4 : std_logic_vector(1 downto 0);
    signal VN575_in5 : std_logic_vector(1 downto 0);
    signal VN576_in0 : std_logic_vector(1 downto 0);
    signal VN576_in1 : std_logic_vector(1 downto 0);
    signal VN576_in2 : std_logic_vector(1 downto 0);
    signal VN576_in3 : std_logic_vector(1 downto 0);
    signal VN576_in4 : std_logic_vector(1 downto 0);
    signal VN576_in5 : std_logic_vector(1 downto 0);
    signal VN577_in0 : std_logic_vector(1 downto 0);
    signal VN577_in1 : std_logic_vector(1 downto 0);
    signal VN577_in2 : std_logic_vector(1 downto 0);
    signal VN577_in3 : std_logic_vector(1 downto 0);
    signal VN577_in4 : std_logic_vector(1 downto 0);
    signal VN577_in5 : std_logic_vector(1 downto 0);
    signal VN578_in0 : std_logic_vector(1 downto 0);
    signal VN578_in1 : std_logic_vector(1 downto 0);
    signal VN578_in2 : std_logic_vector(1 downto 0);
    signal VN578_in3 : std_logic_vector(1 downto 0);
    signal VN578_in4 : std_logic_vector(1 downto 0);
    signal VN578_in5 : std_logic_vector(1 downto 0);
    signal VN579_in0 : std_logic_vector(1 downto 0);
    signal VN579_in1 : std_logic_vector(1 downto 0);
    signal VN579_in2 : std_logic_vector(1 downto 0);
    signal VN579_in3 : std_logic_vector(1 downto 0);
    signal VN579_in4 : std_logic_vector(1 downto 0);
    signal VN579_in5 : std_logic_vector(1 downto 0);
    signal VN580_in0 : std_logic_vector(1 downto 0);
    signal VN580_in1 : std_logic_vector(1 downto 0);
    signal VN580_in2 : std_logic_vector(1 downto 0);
    signal VN580_in3 : std_logic_vector(1 downto 0);
    signal VN580_in4 : std_logic_vector(1 downto 0);
    signal VN580_in5 : std_logic_vector(1 downto 0);
    signal VN581_in0 : std_logic_vector(1 downto 0);
    signal VN581_in1 : std_logic_vector(1 downto 0);
    signal VN581_in2 : std_logic_vector(1 downto 0);
    signal VN581_in3 : std_logic_vector(1 downto 0);
    signal VN581_in4 : std_logic_vector(1 downto 0);
    signal VN581_in5 : std_logic_vector(1 downto 0);
    signal VN582_in0 : std_logic_vector(1 downto 0);
    signal VN582_in1 : std_logic_vector(1 downto 0);
    signal VN582_in2 : std_logic_vector(1 downto 0);
    signal VN582_in3 : std_logic_vector(1 downto 0);
    signal VN582_in4 : std_logic_vector(1 downto 0);
    signal VN582_in5 : std_logic_vector(1 downto 0);
    signal VN583_in0 : std_logic_vector(1 downto 0);
    signal VN583_in1 : std_logic_vector(1 downto 0);
    signal VN583_in2 : std_logic_vector(1 downto 0);
    signal VN583_in3 : std_logic_vector(1 downto 0);
    signal VN583_in4 : std_logic_vector(1 downto 0);
    signal VN583_in5 : std_logic_vector(1 downto 0);
    signal VN584_in0 : std_logic_vector(1 downto 0);
    signal VN584_in1 : std_logic_vector(1 downto 0);
    signal VN584_in2 : std_logic_vector(1 downto 0);
    signal VN584_in3 : std_logic_vector(1 downto 0);
    signal VN584_in4 : std_logic_vector(1 downto 0);
    signal VN584_in5 : std_logic_vector(1 downto 0);
    signal VN585_in0 : std_logic_vector(1 downto 0);
    signal VN585_in1 : std_logic_vector(1 downto 0);
    signal VN585_in2 : std_logic_vector(1 downto 0);
    signal VN585_in3 : std_logic_vector(1 downto 0);
    signal VN585_in4 : std_logic_vector(1 downto 0);
    signal VN585_in5 : std_logic_vector(1 downto 0);
    signal VN586_in0 : std_logic_vector(1 downto 0);
    signal VN586_in1 : std_logic_vector(1 downto 0);
    signal VN586_in2 : std_logic_vector(1 downto 0);
    signal VN586_in3 : std_logic_vector(1 downto 0);
    signal VN586_in4 : std_logic_vector(1 downto 0);
    signal VN586_in5 : std_logic_vector(1 downto 0);
    signal VN587_in0 : std_logic_vector(1 downto 0);
    signal VN587_in1 : std_logic_vector(1 downto 0);
    signal VN587_in2 : std_logic_vector(1 downto 0);
    signal VN587_in3 : std_logic_vector(1 downto 0);
    signal VN587_in4 : std_logic_vector(1 downto 0);
    signal VN587_in5 : std_logic_vector(1 downto 0);
    signal VN588_in0 : std_logic_vector(1 downto 0);
    signal VN588_in1 : std_logic_vector(1 downto 0);
    signal VN588_in2 : std_logic_vector(1 downto 0);
    signal VN588_in3 : std_logic_vector(1 downto 0);
    signal VN588_in4 : std_logic_vector(1 downto 0);
    signal VN588_in5 : std_logic_vector(1 downto 0);
    signal VN589_in0 : std_logic_vector(1 downto 0);
    signal VN589_in1 : std_logic_vector(1 downto 0);
    signal VN589_in2 : std_logic_vector(1 downto 0);
    signal VN589_in3 : std_logic_vector(1 downto 0);
    signal VN589_in4 : std_logic_vector(1 downto 0);
    signal VN589_in5 : std_logic_vector(1 downto 0);
    signal VN590_in0 : std_logic_vector(1 downto 0);
    signal VN590_in1 : std_logic_vector(1 downto 0);
    signal VN590_in2 : std_logic_vector(1 downto 0);
    signal VN590_in3 : std_logic_vector(1 downto 0);
    signal VN590_in4 : std_logic_vector(1 downto 0);
    signal VN590_in5 : std_logic_vector(1 downto 0);
    signal VN591_in0 : std_logic_vector(1 downto 0);
    signal VN591_in1 : std_logic_vector(1 downto 0);
    signal VN591_in2 : std_logic_vector(1 downto 0);
    signal VN591_in3 : std_logic_vector(1 downto 0);
    signal VN591_in4 : std_logic_vector(1 downto 0);
    signal VN591_in5 : std_logic_vector(1 downto 0);
    signal VN592_in0 : std_logic_vector(1 downto 0);
    signal VN592_in1 : std_logic_vector(1 downto 0);
    signal VN592_in2 : std_logic_vector(1 downto 0);
    signal VN592_in3 : std_logic_vector(1 downto 0);
    signal VN592_in4 : std_logic_vector(1 downto 0);
    signal VN592_in5 : std_logic_vector(1 downto 0);
    signal VN593_in0 : std_logic_vector(1 downto 0);
    signal VN593_in1 : std_logic_vector(1 downto 0);
    signal VN593_in2 : std_logic_vector(1 downto 0);
    signal VN593_in3 : std_logic_vector(1 downto 0);
    signal VN593_in4 : std_logic_vector(1 downto 0);
    signal VN593_in5 : std_logic_vector(1 downto 0);
    signal VN594_in0 : std_logic_vector(1 downto 0);
    signal VN594_in1 : std_logic_vector(1 downto 0);
    signal VN594_in2 : std_logic_vector(1 downto 0);
    signal VN594_in3 : std_logic_vector(1 downto 0);
    signal VN594_in4 : std_logic_vector(1 downto 0);
    signal VN594_in5 : std_logic_vector(1 downto 0);
    signal VN595_in0 : std_logic_vector(1 downto 0);
    signal VN595_in1 : std_logic_vector(1 downto 0);
    signal VN595_in2 : std_logic_vector(1 downto 0);
    signal VN595_in3 : std_logic_vector(1 downto 0);
    signal VN595_in4 : std_logic_vector(1 downto 0);
    signal VN595_in5 : std_logic_vector(1 downto 0);
    signal VN596_in0 : std_logic_vector(1 downto 0);
    signal VN596_in1 : std_logic_vector(1 downto 0);
    signal VN596_in2 : std_logic_vector(1 downto 0);
    signal VN596_in3 : std_logic_vector(1 downto 0);
    signal VN596_in4 : std_logic_vector(1 downto 0);
    signal VN596_in5 : std_logic_vector(1 downto 0);
    signal VN597_in0 : std_logic_vector(1 downto 0);
    signal VN597_in1 : std_logic_vector(1 downto 0);
    signal VN597_in2 : std_logic_vector(1 downto 0);
    signal VN597_in3 : std_logic_vector(1 downto 0);
    signal VN597_in4 : std_logic_vector(1 downto 0);
    signal VN597_in5 : std_logic_vector(1 downto 0);
    signal VN598_in0 : std_logic_vector(1 downto 0);
    signal VN598_in1 : std_logic_vector(1 downto 0);
    signal VN598_in2 : std_logic_vector(1 downto 0);
    signal VN598_in3 : std_logic_vector(1 downto 0);
    signal VN598_in4 : std_logic_vector(1 downto 0);
    signal VN598_in5 : std_logic_vector(1 downto 0);
    signal VN599_in0 : std_logic_vector(1 downto 0);
    signal VN599_in1 : std_logic_vector(1 downto 0);
    signal VN599_in2 : std_logic_vector(1 downto 0);
    signal VN599_in3 : std_logic_vector(1 downto 0);
    signal VN599_in4 : std_logic_vector(1 downto 0);
    signal VN599_in5 : std_logic_vector(1 downto 0);
    signal VN600_in0 : std_logic_vector(1 downto 0);
    signal VN600_in1 : std_logic_vector(1 downto 0);
    signal VN600_in2 : std_logic_vector(1 downto 0);
    signal VN600_in3 : std_logic_vector(1 downto 0);
    signal VN600_in4 : std_logic_vector(1 downto 0);
    signal VN600_in5 : std_logic_vector(1 downto 0);
    signal VN601_in0 : std_logic_vector(1 downto 0);
    signal VN601_in1 : std_logic_vector(1 downto 0);
    signal VN601_in2 : std_logic_vector(1 downto 0);
    signal VN601_in3 : std_logic_vector(1 downto 0);
    signal VN601_in4 : std_logic_vector(1 downto 0);
    signal VN601_in5 : std_logic_vector(1 downto 0);
    signal VN602_in0 : std_logic_vector(1 downto 0);
    signal VN602_in1 : std_logic_vector(1 downto 0);
    signal VN602_in2 : std_logic_vector(1 downto 0);
    signal VN602_in3 : std_logic_vector(1 downto 0);
    signal VN602_in4 : std_logic_vector(1 downto 0);
    signal VN602_in5 : std_logic_vector(1 downto 0);
    signal VN603_in0 : std_logic_vector(1 downto 0);
    signal VN603_in1 : std_logic_vector(1 downto 0);
    signal VN603_in2 : std_logic_vector(1 downto 0);
    signal VN603_in3 : std_logic_vector(1 downto 0);
    signal VN603_in4 : std_logic_vector(1 downto 0);
    signal VN603_in5 : std_logic_vector(1 downto 0);
    signal VN604_in0 : std_logic_vector(1 downto 0);
    signal VN604_in1 : std_logic_vector(1 downto 0);
    signal VN604_in2 : std_logic_vector(1 downto 0);
    signal VN604_in3 : std_logic_vector(1 downto 0);
    signal VN604_in4 : std_logic_vector(1 downto 0);
    signal VN604_in5 : std_logic_vector(1 downto 0);
    signal VN605_in0 : std_logic_vector(1 downto 0);
    signal VN605_in1 : std_logic_vector(1 downto 0);
    signal VN605_in2 : std_logic_vector(1 downto 0);
    signal VN605_in3 : std_logic_vector(1 downto 0);
    signal VN605_in4 : std_logic_vector(1 downto 0);
    signal VN605_in5 : std_logic_vector(1 downto 0);
    signal VN606_in0 : std_logic_vector(1 downto 0);
    signal VN606_in1 : std_logic_vector(1 downto 0);
    signal VN606_in2 : std_logic_vector(1 downto 0);
    signal VN606_in3 : std_logic_vector(1 downto 0);
    signal VN606_in4 : std_logic_vector(1 downto 0);
    signal VN606_in5 : std_logic_vector(1 downto 0);
    signal VN607_in0 : std_logic_vector(1 downto 0);
    signal VN607_in1 : std_logic_vector(1 downto 0);
    signal VN607_in2 : std_logic_vector(1 downto 0);
    signal VN607_in3 : std_logic_vector(1 downto 0);
    signal VN607_in4 : std_logic_vector(1 downto 0);
    signal VN607_in5 : std_logic_vector(1 downto 0);
    signal VN608_in0 : std_logic_vector(1 downto 0);
    signal VN608_in1 : std_logic_vector(1 downto 0);
    signal VN608_in2 : std_logic_vector(1 downto 0);
    signal VN608_in3 : std_logic_vector(1 downto 0);
    signal VN608_in4 : std_logic_vector(1 downto 0);
    signal VN608_in5 : std_logic_vector(1 downto 0);
    signal VN609_in0 : std_logic_vector(1 downto 0);
    signal VN609_in1 : std_logic_vector(1 downto 0);
    signal VN609_in2 : std_logic_vector(1 downto 0);
    signal VN609_in3 : std_logic_vector(1 downto 0);
    signal VN609_in4 : std_logic_vector(1 downto 0);
    signal VN609_in5 : std_logic_vector(1 downto 0);
    signal VN610_in0 : std_logic_vector(1 downto 0);
    signal VN610_in1 : std_logic_vector(1 downto 0);
    signal VN610_in2 : std_logic_vector(1 downto 0);
    signal VN610_in3 : std_logic_vector(1 downto 0);
    signal VN610_in4 : std_logic_vector(1 downto 0);
    signal VN610_in5 : std_logic_vector(1 downto 0);
    signal VN611_in0 : std_logic_vector(1 downto 0);
    signal VN611_in1 : std_logic_vector(1 downto 0);
    signal VN611_in2 : std_logic_vector(1 downto 0);
    signal VN611_in3 : std_logic_vector(1 downto 0);
    signal VN611_in4 : std_logic_vector(1 downto 0);
    signal VN611_in5 : std_logic_vector(1 downto 0);
    signal VN612_in0 : std_logic_vector(1 downto 0);
    signal VN612_in1 : std_logic_vector(1 downto 0);
    signal VN612_in2 : std_logic_vector(1 downto 0);
    signal VN612_in3 : std_logic_vector(1 downto 0);
    signal VN612_in4 : std_logic_vector(1 downto 0);
    signal VN612_in5 : std_logic_vector(1 downto 0);
    signal VN613_in0 : std_logic_vector(1 downto 0);
    signal VN613_in1 : std_logic_vector(1 downto 0);
    signal VN613_in2 : std_logic_vector(1 downto 0);
    signal VN613_in3 : std_logic_vector(1 downto 0);
    signal VN613_in4 : std_logic_vector(1 downto 0);
    signal VN613_in5 : std_logic_vector(1 downto 0);
    signal VN614_in0 : std_logic_vector(1 downto 0);
    signal VN614_in1 : std_logic_vector(1 downto 0);
    signal VN614_in2 : std_logic_vector(1 downto 0);
    signal VN614_in3 : std_logic_vector(1 downto 0);
    signal VN614_in4 : std_logic_vector(1 downto 0);
    signal VN614_in5 : std_logic_vector(1 downto 0);
    signal VN615_in0 : std_logic_vector(1 downto 0);
    signal VN615_in1 : std_logic_vector(1 downto 0);
    signal VN615_in2 : std_logic_vector(1 downto 0);
    signal VN615_in3 : std_logic_vector(1 downto 0);
    signal VN615_in4 : std_logic_vector(1 downto 0);
    signal VN615_in5 : std_logic_vector(1 downto 0);
    signal VN616_in0 : std_logic_vector(1 downto 0);
    signal VN616_in1 : std_logic_vector(1 downto 0);
    signal VN616_in2 : std_logic_vector(1 downto 0);
    signal VN616_in3 : std_logic_vector(1 downto 0);
    signal VN616_in4 : std_logic_vector(1 downto 0);
    signal VN616_in5 : std_logic_vector(1 downto 0);
    signal VN617_in0 : std_logic_vector(1 downto 0);
    signal VN617_in1 : std_logic_vector(1 downto 0);
    signal VN617_in2 : std_logic_vector(1 downto 0);
    signal VN617_in3 : std_logic_vector(1 downto 0);
    signal VN617_in4 : std_logic_vector(1 downto 0);
    signal VN617_in5 : std_logic_vector(1 downto 0);
    signal VN618_in0 : std_logic_vector(1 downto 0);
    signal VN618_in1 : std_logic_vector(1 downto 0);
    signal VN618_in2 : std_logic_vector(1 downto 0);
    signal VN618_in3 : std_logic_vector(1 downto 0);
    signal VN618_in4 : std_logic_vector(1 downto 0);
    signal VN618_in5 : std_logic_vector(1 downto 0);
    signal VN619_in0 : std_logic_vector(1 downto 0);
    signal VN619_in1 : std_logic_vector(1 downto 0);
    signal VN619_in2 : std_logic_vector(1 downto 0);
    signal VN619_in3 : std_logic_vector(1 downto 0);
    signal VN619_in4 : std_logic_vector(1 downto 0);
    signal VN619_in5 : std_logic_vector(1 downto 0);
    signal VN620_in0 : std_logic_vector(1 downto 0);
    signal VN620_in1 : std_logic_vector(1 downto 0);
    signal VN620_in2 : std_logic_vector(1 downto 0);
    signal VN620_in3 : std_logic_vector(1 downto 0);
    signal VN620_in4 : std_logic_vector(1 downto 0);
    signal VN620_in5 : std_logic_vector(1 downto 0);
    signal VN621_in0 : std_logic_vector(1 downto 0);
    signal VN621_in1 : std_logic_vector(1 downto 0);
    signal VN621_in2 : std_logic_vector(1 downto 0);
    signal VN621_in3 : std_logic_vector(1 downto 0);
    signal VN621_in4 : std_logic_vector(1 downto 0);
    signal VN621_in5 : std_logic_vector(1 downto 0);
    signal VN622_in0 : std_logic_vector(1 downto 0);
    signal VN622_in1 : std_logic_vector(1 downto 0);
    signal VN622_in2 : std_logic_vector(1 downto 0);
    signal VN622_in3 : std_logic_vector(1 downto 0);
    signal VN622_in4 : std_logic_vector(1 downto 0);
    signal VN622_in5 : std_logic_vector(1 downto 0);
    signal VN623_in0 : std_logic_vector(1 downto 0);
    signal VN623_in1 : std_logic_vector(1 downto 0);
    signal VN623_in2 : std_logic_vector(1 downto 0);
    signal VN623_in3 : std_logic_vector(1 downto 0);
    signal VN623_in4 : std_logic_vector(1 downto 0);
    signal VN623_in5 : std_logic_vector(1 downto 0);
    signal VN624_in0 : std_logic_vector(1 downto 0);
    signal VN624_in1 : std_logic_vector(1 downto 0);
    signal VN624_in2 : std_logic_vector(1 downto 0);
    signal VN624_in3 : std_logic_vector(1 downto 0);
    signal VN624_in4 : std_logic_vector(1 downto 0);
    signal VN624_in5 : std_logic_vector(1 downto 0);
    signal VN625_in0 : std_logic_vector(1 downto 0);
    signal VN625_in1 : std_logic_vector(1 downto 0);
    signal VN625_in2 : std_logic_vector(1 downto 0);
    signal VN625_in3 : std_logic_vector(1 downto 0);
    signal VN625_in4 : std_logic_vector(1 downto 0);
    signal VN625_in5 : std_logic_vector(1 downto 0);
    signal VN626_in0 : std_logic_vector(1 downto 0);
    signal VN626_in1 : std_logic_vector(1 downto 0);
    signal VN626_in2 : std_logic_vector(1 downto 0);
    signal VN626_in3 : std_logic_vector(1 downto 0);
    signal VN626_in4 : std_logic_vector(1 downto 0);
    signal VN626_in5 : std_logic_vector(1 downto 0);
    signal VN627_in0 : std_logic_vector(1 downto 0);
    signal VN627_in1 : std_logic_vector(1 downto 0);
    signal VN627_in2 : std_logic_vector(1 downto 0);
    signal VN627_in3 : std_logic_vector(1 downto 0);
    signal VN627_in4 : std_logic_vector(1 downto 0);
    signal VN627_in5 : std_logic_vector(1 downto 0);
    signal VN628_in0 : std_logic_vector(1 downto 0);
    signal VN628_in1 : std_logic_vector(1 downto 0);
    signal VN628_in2 : std_logic_vector(1 downto 0);
    signal VN628_in3 : std_logic_vector(1 downto 0);
    signal VN628_in4 : std_logic_vector(1 downto 0);
    signal VN628_in5 : std_logic_vector(1 downto 0);
    signal VN629_in0 : std_logic_vector(1 downto 0);
    signal VN629_in1 : std_logic_vector(1 downto 0);
    signal VN629_in2 : std_logic_vector(1 downto 0);
    signal VN629_in3 : std_logic_vector(1 downto 0);
    signal VN629_in4 : std_logic_vector(1 downto 0);
    signal VN629_in5 : std_logic_vector(1 downto 0);
    signal VN630_in0 : std_logic_vector(1 downto 0);
    signal VN630_in1 : std_logic_vector(1 downto 0);
    signal VN630_in2 : std_logic_vector(1 downto 0);
    signal VN630_in3 : std_logic_vector(1 downto 0);
    signal VN630_in4 : std_logic_vector(1 downto 0);
    signal VN630_in5 : std_logic_vector(1 downto 0);
    signal VN631_in0 : std_logic_vector(1 downto 0);
    signal VN631_in1 : std_logic_vector(1 downto 0);
    signal VN631_in2 : std_logic_vector(1 downto 0);
    signal VN631_in3 : std_logic_vector(1 downto 0);
    signal VN631_in4 : std_logic_vector(1 downto 0);
    signal VN631_in5 : std_logic_vector(1 downto 0);
    signal VN632_in0 : std_logic_vector(1 downto 0);
    signal VN632_in1 : std_logic_vector(1 downto 0);
    signal VN632_in2 : std_logic_vector(1 downto 0);
    signal VN632_in3 : std_logic_vector(1 downto 0);
    signal VN632_in4 : std_logic_vector(1 downto 0);
    signal VN632_in5 : std_logic_vector(1 downto 0);
    signal VN633_in0 : std_logic_vector(1 downto 0);
    signal VN633_in1 : std_logic_vector(1 downto 0);
    signal VN633_in2 : std_logic_vector(1 downto 0);
    signal VN633_in3 : std_logic_vector(1 downto 0);
    signal VN633_in4 : std_logic_vector(1 downto 0);
    signal VN633_in5 : std_logic_vector(1 downto 0);
    signal VN634_in0 : std_logic_vector(1 downto 0);
    signal VN634_in1 : std_logic_vector(1 downto 0);
    signal VN634_in2 : std_logic_vector(1 downto 0);
    signal VN634_in3 : std_logic_vector(1 downto 0);
    signal VN634_in4 : std_logic_vector(1 downto 0);
    signal VN634_in5 : std_logic_vector(1 downto 0);
    signal VN635_in0 : std_logic_vector(1 downto 0);
    signal VN635_in1 : std_logic_vector(1 downto 0);
    signal VN635_in2 : std_logic_vector(1 downto 0);
    signal VN635_in3 : std_logic_vector(1 downto 0);
    signal VN635_in4 : std_logic_vector(1 downto 0);
    signal VN635_in5 : std_logic_vector(1 downto 0);
    signal VN636_in0 : std_logic_vector(1 downto 0);
    signal VN636_in1 : std_logic_vector(1 downto 0);
    signal VN636_in2 : std_logic_vector(1 downto 0);
    signal VN636_in3 : std_logic_vector(1 downto 0);
    signal VN636_in4 : std_logic_vector(1 downto 0);
    signal VN636_in5 : std_logic_vector(1 downto 0);
    signal VN637_in0 : std_logic_vector(1 downto 0);
    signal VN637_in1 : std_logic_vector(1 downto 0);
    signal VN637_in2 : std_logic_vector(1 downto 0);
    signal VN637_in3 : std_logic_vector(1 downto 0);
    signal VN637_in4 : std_logic_vector(1 downto 0);
    signal VN637_in5 : std_logic_vector(1 downto 0);
    signal VN638_in0 : std_logic_vector(1 downto 0);
    signal VN638_in1 : std_logic_vector(1 downto 0);
    signal VN638_in2 : std_logic_vector(1 downto 0);
    signal VN638_in3 : std_logic_vector(1 downto 0);
    signal VN638_in4 : std_logic_vector(1 downto 0);
    signal VN638_in5 : std_logic_vector(1 downto 0);
    signal VN639_in0 : std_logic_vector(1 downto 0);
    signal VN639_in1 : std_logic_vector(1 downto 0);
    signal VN639_in2 : std_logic_vector(1 downto 0);
    signal VN639_in3 : std_logic_vector(1 downto 0);
    signal VN639_in4 : std_logic_vector(1 downto 0);
    signal VN639_in5 : std_logic_vector(1 downto 0);
    signal VN640_in0 : std_logic_vector(1 downto 0);
    signal VN640_in1 : std_logic_vector(1 downto 0);
    signal VN640_in2 : std_logic_vector(1 downto 0);
    signal VN640_in3 : std_logic_vector(1 downto 0);
    signal VN640_in4 : std_logic_vector(1 downto 0);
    signal VN640_in5 : std_logic_vector(1 downto 0);
    signal VN641_in0 : std_logic_vector(1 downto 0);
    signal VN641_in1 : std_logic_vector(1 downto 0);
    signal VN641_in2 : std_logic_vector(1 downto 0);
    signal VN641_in3 : std_logic_vector(1 downto 0);
    signal VN641_in4 : std_logic_vector(1 downto 0);
    signal VN641_in5 : std_logic_vector(1 downto 0);
    signal VN642_in0 : std_logic_vector(1 downto 0);
    signal VN642_in1 : std_logic_vector(1 downto 0);
    signal VN642_in2 : std_logic_vector(1 downto 0);
    signal VN642_in3 : std_logic_vector(1 downto 0);
    signal VN642_in4 : std_logic_vector(1 downto 0);
    signal VN642_in5 : std_logic_vector(1 downto 0);
    signal VN643_in0 : std_logic_vector(1 downto 0);
    signal VN643_in1 : std_logic_vector(1 downto 0);
    signal VN643_in2 : std_logic_vector(1 downto 0);
    signal VN643_in3 : std_logic_vector(1 downto 0);
    signal VN643_in4 : std_logic_vector(1 downto 0);
    signal VN643_in5 : std_logic_vector(1 downto 0);
    signal VN644_in0 : std_logic_vector(1 downto 0);
    signal VN644_in1 : std_logic_vector(1 downto 0);
    signal VN644_in2 : std_logic_vector(1 downto 0);
    signal VN644_in3 : std_logic_vector(1 downto 0);
    signal VN644_in4 : std_logic_vector(1 downto 0);
    signal VN644_in5 : std_logic_vector(1 downto 0);
    signal VN645_in0 : std_logic_vector(1 downto 0);
    signal VN645_in1 : std_logic_vector(1 downto 0);
    signal VN645_in2 : std_logic_vector(1 downto 0);
    signal VN645_in3 : std_logic_vector(1 downto 0);
    signal VN645_in4 : std_logic_vector(1 downto 0);
    signal VN645_in5 : std_logic_vector(1 downto 0);
    signal VN646_in0 : std_logic_vector(1 downto 0);
    signal VN646_in1 : std_logic_vector(1 downto 0);
    signal VN646_in2 : std_logic_vector(1 downto 0);
    signal VN646_in3 : std_logic_vector(1 downto 0);
    signal VN646_in4 : std_logic_vector(1 downto 0);
    signal VN646_in5 : std_logic_vector(1 downto 0);
    signal VN647_in0 : std_logic_vector(1 downto 0);
    signal VN647_in1 : std_logic_vector(1 downto 0);
    signal VN647_in2 : std_logic_vector(1 downto 0);
    signal VN647_in3 : std_logic_vector(1 downto 0);
    signal VN647_in4 : std_logic_vector(1 downto 0);
    signal VN647_in5 : std_logic_vector(1 downto 0);
    signal VN648_in0 : std_logic_vector(1 downto 0);
    signal VN648_in1 : std_logic_vector(1 downto 0);
    signal VN648_in2 : std_logic_vector(1 downto 0);
    signal VN648_in3 : std_logic_vector(1 downto 0);
    signal VN648_in4 : std_logic_vector(1 downto 0);
    signal VN648_in5 : std_logic_vector(1 downto 0);
    signal VN649_in0 : std_logic_vector(1 downto 0);
    signal VN649_in1 : std_logic_vector(1 downto 0);
    signal VN649_in2 : std_logic_vector(1 downto 0);
    signal VN649_in3 : std_logic_vector(1 downto 0);
    signal VN649_in4 : std_logic_vector(1 downto 0);
    signal VN649_in5 : std_logic_vector(1 downto 0);
    signal VN650_in0 : std_logic_vector(1 downto 0);
    signal VN650_in1 : std_logic_vector(1 downto 0);
    signal VN650_in2 : std_logic_vector(1 downto 0);
    signal VN650_in3 : std_logic_vector(1 downto 0);
    signal VN650_in4 : std_logic_vector(1 downto 0);
    signal VN650_in5 : std_logic_vector(1 downto 0);
    signal VN651_in0 : std_logic_vector(1 downto 0);
    signal VN651_in1 : std_logic_vector(1 downto 0);
    signal VN651_in2 : std_logic_vector(1 downto 0);
    signal VN651_in3 : std_logic_vector(1 downto 0);
    signal VN651_in4 : std_logic_vector(1 downto 0);
    signal VN651_in5 : std_logic_vector(1 downto 0);
    signal VN652_in0 : std_logic_vector(1 downto 0);
    signal VN652_in1 : std_logic_vector(1 downto 0);
    signal VN652_in2 : std_logic_vector(1 downto 0);
    signal VN652_in3 : std_logic_vector(1 downto 0);
    signal VN652_in4 : std_logic_vector(1 downto 0);
    signal VN652_in5 : std_logic_vector(1 downto 0);
    signal VN653_in0 : std_logic_vector(1 downto 0);
    signal VN653_in1 : std_logic_vector(1 downto 0);
    signal VN653_in2 : std_logic_vector(1 downto 0);
    signal VN653_in3 : std_logic_vector(1 downto 0);
    signal VN653_in4 : std_logic_vector(1 downto 0);
    signal VN653_in5 : std_logic_vector(1 downto 0);
    signal VN654_in0 : std_logic_vector(1 downto 0);
    signal VN654_in1 : std_logic_vector(1 downto 0);
    signal VN654_in2 : std_logic_vector(1 downto 0);
    signal VN654_in3 : std_logic_vector(1 downto 0);
    signal VN654_in4 : std_logic_vector(1 downto 0);
    signal VN654_in5 : std_logic_vector(1 downto 0);
    signal VN655_in0 : std_logic_vector(1 downto 0);
    signal VN655_in1 : std_logic_vector(1 downto 0);
    signal VN655_in2 : std_logic_vector(1 downto 0);
    signal VN655_in3 : std_logic_vector(1 downto 0);
    signal VN655_in4 : std_logic_vector(1 downto 0);
    signal VN655_in5 : std_logic_vector(1 downto 0);
    signal VN656_in0 : std_logic_vector(1 downto 0);
    signal VN656_in1 : std_logic_vector(1 downto 0);
    signal VN656_in2 : std_logic_vector(1 downto 0);
    signal VN656_in3 : std_logic_vector(1 downto 0);
    signal VN656_in4 : std_logic_vector(1 downto 0);
    signal VN656_in5 : std_logic_vector(1 downto 0);
    signal VN657_in0 : std_logic_vector(1 downto 0);
    signal VN657_in1 : std_logic_vector(1 downto 0);
    signal VN657_in2 : std_logic_vector(1 downto 0);
    signal VN657_in3 : std_logic_vector(1 downto 0);
    signal VN657_in4 : std_logic_vector(1 downto 0);
    signal VN657_in5 : std_logic_vector(1 downto 0);
    signal VN658_in0 : std_logic_vector(1 downto 0);
    signal VN658_in1 : std_logic_vector(1 downto 0);
    signal VN658_in2 : std_logic_vector(1 downto 0);
    signal VN658_in3 : std_logic_vector(1 downto 0);
    signal VN658_in4 : std_logic_vector(1 downto 0);
    signal VN658_in5 : std_logic_vector(1 downto 0);
    signal VN659_in0 : std_logic_vector(1 downto 0);
    signal VN659_in1 : std_logic_vector(1 downto 0);
    signal VN659_in2 : std_logic_vector(1 downto 0);
    signal VN659_in3 : std_logic_vector(1 downto 0);
    signal VN659_in4 : std_logic_vector(1 downto 0);
    signal VN659_in5 : std_logic_vector(1 downto 0);
    signal VN660_in0 : std_logic_vector(1 downto 0);
    signal VN660_in1 : std_logic_vector(1 downto 0);
    signal VN660_in2 : std_logic_vector(1 downto 0);
    signal VN660_in3 : std_logic_vector(1 downto 0);
    signal VN660_in4 : std_logic_vector(1 downto 0);
    signal VN660_in5 : std_logic_vector(1 downto 0);
    signal VN661_in0 : std_logic_vector(1 downto 0);
    signal VN661_in1 : std_logic_vector(1 downto 0);
    signal VN661_in2 : std_logic_vector(1 downto 0);
    signal VN661_in3 : std_logic_vector(1 downto 0);
    signal VN661_in4 : std_logic_vector(1 downto 0);
    signal VN661_in5 : std_logic_vector(1 downto 0);
    signal VN662_in0 : std_logic_vector(1 downto 0);
    signal VN662_in1 : std_logic_vector(1 downto 0);
    signal VN662_in2 : std_logic_vector(1 downto 0);
    signal VN662_in3 : std_logic_vector(1 downto 0);
    signal VN662_in4 : std_logic_vector(1 downto 0);
    signal VN662_in5 : std_logic_vector(1 downto 0);
    signal VN663_in0 : std_logic_vector(1 downto 0);
    signal VN663_in1 : std_logic_vector(1 downto 0);
    signal VN663_in2 : std_logic_vector(1 downto 0);
    signal VN663_in3 : std_logic_vector(1 downto 0);
    signal VN663_in4 : std_logic_vector(1 downto 0);
    signal VN663_in5 : std_logic_vector(1 downto 0);
    signal VN664_in0 : std_logic_vector(1 downto 0);
    signal VN664_in1 : std_logic_vector(1 downto 0);
    signal VN664_in2 : std_logic_vector(1 downto 0);
    signal VN664_in3 : std_logic_vector(1 downto 0);
    signal VN664_in4 : std_logic_vector(1 downto 0);
    signal VN664_in5 : std_logic_vector(1 downto 0);
    signal VN665_in0 : std_logic_vector(1 downto 0);
    signal VN665_in1 : std_logic_vector(1 downto 0);
    signal VN665_in2 : std_logic_vector(1 downto 0);
    signal VN665_in3 : std_logic_vector(1 downto 0);
    signal VN665_in4 : std_logic_vector(1 downto 0);
    signal VN665_in5 : std_logic_vector(1 downto 0);
    signal VN666_in0 : std_logic_vector(1 downto 0);
    signal VN666_in1 : std_logic_vector(1 downto 0);
    signal VN666_in2 : std_logic_vector(1 downto 0);
    signal VN666_in3 : std_logic_vector(1 downto 0);
    signal VN666_in4 : std_logic_vector(1 downto 0);
    signal VN666_in5 : std_logic_vector(1 downto 0);
    signal VN667_in0 : std_logic_vector(1 downto 0);
    signal VN667_in1 : std_logic_vector(1 downto 0);
    signal VN667_in2 : std_logic_vector(1 downto 0);
    signal VN667_in3 : std_logic_vector(1 downto 0);
    signal VN667_in4 : std_logic_vector(1 downto 0);
    signal VN667_in5 : std_logic_vector(1 downto 0);
    signal VN668_in0 : std_logic_vector(1 downto 0);
    signal VN668_in1 : std_logic_vector(1 downto 0);
    signal VN668_in2 : std_logic_vector(1 downto 0);
    signal VN668_in3 : std_logic_vector(1 downto 0);
    signal VN668_in4 : std_logic_vector(1 downto 0);
    signal VN668_in5 : std_logic_vector(1 downto 0);
    signal VN669_in0 : std_logic_vector(1 downto 0);
    signal VN669_in1 : std_logic_vector(1 downto 0);
    signal VN669_in2 : std_logic_vector(1 downto 0);
    signal VN669_in3 : std_logic_vector(1 downto 0);
    signal VN669_in4 : std_logic_vector(1 downto 0);
    signal VN669_in5 : std_logic_vector(1 downto 0);
    signal VN670_in0 : std_logic_vector(1 downto 0);
    signal VN670_in1 : std_logic_vector(1 downto 0);
    signal VN670_in2 : std_logic_vector(1 downto 0);
    signal VN670_in3 : std_logic_vector(1 downto 0);
    signal VN670_in4 : std_logic_vector(1 downto 0);
    signal VN670_in5 : std_logic_vector(1 downto 0);
    signal VN671_in0 : std_logic_vector(1 downto 0);
    signal VN671_in1 : std_logic_vector(1 downto 0);
    signal VN671_in2 : std_logic_vector(1 downto 0);
    signal VN671_in3 : std_logic_vector(1 downto 0);
    signal VN671_in4 : std_logic_vector(1 downto 0);
    signal VN671_in5 : std_logic_vector(1 downto 0);
    signal VN672_in0 : std_logic_vector(1 downto 0);
    signal VN672_in1 : std_logic_vector(1 downto 0);
    signal VN672_in2 : std_logic_vector(1 downto 0);
    signal VN672_in3 : std_logic_vector(1 downto 0);
    signal VN672_in4 : std_logic_vector(1 downto 0);
    signal VN672_in5 : std_logic_vector(1 downto 0);
    signal VN673_in0 : std_logic_vector(1 downto 0);
    signal VN673_in1 : std_logic_vector(1 downto 0);
    signal VN673_in2 : std_logic_vector(1 downto 0);
    signal VN673_in3 : std_logic_vector(1 downto 0);
    signal VN673_in4 : std_logic_vector(1 downto 0);
    signal VN673_in5 : std_logic_vector(1 downto 0);
    signal VN674_in0 : std_logic_vector(1 downto 0);
    signal VN674_in1 : std_logic_vector(1 downto 0);
    signal VN674_in2 : std_logic_vector(1 downto 0);
    signal VN674_in3 : std_logic_vector(1 downto 0);
    signal VN674_in4 : std_logic_vector(1 downto 0);
    signal VN674_in5 : std_logic_vector(1 downto 0);
    signal VN675_in0 : std_logic_vector(1 downto 0);
    signal VN675_in1 : std_logic_vector(1 downto 0);
    signal VN675_in2 : std_logic_vector(1 downto 0);
    signal VN675_in3 : std_logic_vector(1 downto 0);
    signal VN675_in4 : std_logic_vector(1 downto 0);
    signal VN675_in5 : std_logic_vector(1 downto 0);
    signal VN676_in0 : std_logic_vector(1 downto 0);
    signal VN676_in1 : std_logic_vector(1 downto 0);
    signal VN676_in2 : std_logic_vector(1 downto 0);
    signal VN676_in3 : std_logic_vector(1 downto 0);
    signal VN676_in4 : std_logic_vector(1 downto 0);
    signal VN676_in5 : std_logic_vector(1 downto 0);
    signal VN677_in0 : std_logic_vector(1 downto 0);
    signal VN677_in1 : std_logic_vector(1 downto 0);
    signal VN677_in2 : std_logic_vector(1 downto 0);
    signal VN677_in3 : std_logic_vector(1 downto 0);
    signal VN677_in4 : std_logic_vector(1 downto 0);
    signal VN677_in5 : std_logic_vector(1 downto 0);
    signal VN678_in0 : std_logic_vector(1 downto 0);
    signal VN678_in1 : std_logic_vector(1 downto 0);
    signal VN678_in2 : std_logic_vector(1 downto 0);
    signal VN678_in3 : std_logic_vector(1 downto 0);
    signal VN678_in4 : std_logic_vector(1 downto 0);
    signal VN678_in5 : std_logic_vector(1 downto 0);
    signal VN679_in0 : std_logic_vector(1 downto 0);
    signal VN679_in1 : std_logic_vector(1 downto 0);
    signal VN679_in2 : std_logic_vector(1 downto 0);
    signal VN679_in3 : std_logic_vector(1 downto 0);
    signal VN679_in4 : std_logic_vector(1 downto 0);
    signal VN679_in5 : std_logic_vector(1 downto 0);
    signal VN680_in0 : std_logic_vector(1 downto 0);
    signal VN680_in1 : std_logic_vector(1 downto 0);
    signal VN680_in2 : std_logic_vector(1 downto 0);
    signal VN680_in3 : std_logic_vector(1 downto 0);
    signal VN680_in4 : std_logic_vector(1 downto 0);
    signal VN680_in5 : std_logic_vector(1 downto 0);
    signal VN681_in0 : std_logic_vector(1 downto 0);
    signal VN681_in1 : std_logic_vector(1 downto 0);
    signal VN681_in2 : std_logic_vector(1 downto 0);
    signal VN681_in3 : std_logic_vector(1 downto 0);
    signal VN681_in4 : std_logic_vector(1 downto 0);
    signal VN681_in5 : std_logic_vector(1 downto 0);
    signal VN682_in0 : std_logic_vector(1 downto 0);
    signal VN682_in1 : std_logic_vector(1 downto 0);
    signal VN682_in2 : std_logic_vector(1 downto 0);
    signal VN682_in3 : std_logic_vector(1 downto 0);
    signal VN682_in4 : std_logic_vector(1 downto 0);
    signal VN682_in5 : std_logic_vector(1 downto 0);
    signal VN683_in0 : std_logic_vector(1 downto 0);
    signal VN683_in1 : std_logic_vector(1 downto 0);
    signal VN683_in2 : std_logic_vector(1 downto 0);
    signal VN683_in3 : std_logic_vector(1 downto 0);
    signal VN683_in4 : std_logic_vector(1 downto 0);
    signal VN683_in5 : std_logic_vector(1 downto 0);
    signal VN684_in0 : std_logic_vector(1 downto 0);
    signal VN684_in1 : std_logic_vector(1 downto 0);
    signal VN684_in2 : std_logic_vector(1 downto 0);
    signal VN684_in3 : std_logic_vector(1 downto 0);
    signal VN684_in4 : std_logic_vector(1 downto 0);
    signal VN684_in5 : std_logic_vector(1 downto 0);
    signal VN685_in0 : std_logic_vector(1 downto 0);
    signal VN685_in1 : std_logic_vector(1 downto 0);
    signal VN685_in2 : std_logic_vector(1 downto 0);
    signal VN685_in3 : std_logic_vector(1 downto 0);
    signal VN685_in4 : std_logic_vector(1 downto 0);
    signal VN685_in5 : std_logic_vector(1 downto 0);
    signal VN686_in0 : std_logic_vector(1 downto 0);
    signal VN686_in1 : std_logic_vector(1 downto 0);
    signal VN686_in2 : std_logic_vector(1 downto 0);
    signal VN686_in3 : std_logic_vector(1 downto 0);
    signal VN686_in4 : std_logic_vector(1 downto 0);
    signal VN686_in5 : std_logic_vector(1 downto 0);
    signal VN687_in0 : std_logic_vector(1 downto 0);
    signal VN687_in1 : std_logic_vector(1 downto 0);
    signal VN687_in2 : std_logic_vector(1 downto 0);
    signal VN687_in3 : std_logic_vector(1 downto 0);
    signal VN687_in4 : std_logic_vector(1 downto 0);
    signal VN687_in5 : std_logic_vector(1 downto 0);
    signal VN688_in0 : std_logic_vector(1 downto 0);
    signal VN688_in1 : std_logic_vector(1 downto 0);
    signal VN688_in2 : std_logic_vector(1 downto 0);
    signal VN688_in3 : std_logic_vector(1 downto 0);
    signal VN688_in4 : std_logic_vector(1 downto 0);
    signal VN688_in5 : std_logic_vector(1 downto 0);
    signal VN689_in0 : std_logic_vector(1 downto 0);
    signal VN689_in1 : std_logic_vector(1 downto 0);
    signal VN689_in2 : std_logic_vector(1 downto 0);
    signal VN689_in3 : std_logic_vector(1 downto 0);
    signal VN689_in4 : std_logic_vector(1 downto 0);
    signal VN689_in5 : std_logic_vector(1 downto 0);
    signal VN690_in0 : std_logic_vector(1 downto 0);
    signal VN690_in1 : std_logic_vector(1 downto 0);
    signal VN690_in2 : std_logic_vector(1 downto 0);
    signal VN690_in3 : std_logic_vector(1 downto 0);
    signal VN690_in4 : std_logic_vector(1 downto 0);
    signal VN690_in5 : std_logic_vector(1 downto 0);
    signal VN691_in0 : std_logic_vector(1 downto 0);
    signal VN691_in1 : std_logic_vector(1 downto 0);
    signal VN691_in2 : std_logic_vector(1 downto 0);
    signal VN691_in3 : std_logic_vector(1 downto 0);
    signal VN691_in4 : std_logic_vector(1 downto 0);
    signal VN691_in5 : std_logic_vector(1 downto 0);
    signal VN692_in0 : std_logic_vector(1 downto 0);
    signal VN692_in1 : std_logic_vector(1 downto 0);
    signal VN692_in2 : std_logic_vector(1 downto 0);
    signal VN692_in3 : std_logic_vector(1 downto 0);
    signal VN692_in4 : std_logic_vector(1 downto 0);
    signal VN692_in5 : std_logic_vector(1 downto 0);
    signal VN693_in0 : std_logic_vector(1 downto 0);
    signal VN693_in1 : std_logic_vector(1 downto 0);
    signal VN693_in2 : std_logic_vector(1 downto 0);
    signal VN693_in3 : std_logic_vector(1 downto 0);
    signal VN693_in4 : std_logic_vector(1 downto 0);
    signal VN693_in5 : std_logic_vector(1 downto 0);
    signal VN694_in0 : std_logic_vector(1 downto 0);
    signal VN694_in1 : std_logic_vector(1 downto 0);
    signal VN694_in2 : std_logic_vector(1 downto 0);
    signal VN694_in3 : std_logic_vector(1 downto 0);
    signal VN694_in4 : std_logic_vector(1 downto 0);
    signal VN694_in5 : std_logic_vector(1 downto 0);
    signal VN695_in0 : std_logic_vector(1 downto 0);
    signal VN695_in1 : std_logic_vector(1 downto 0);
    signal VN695_in2 : std_logic_vector(1 downto 0);
    signal VN695_in3 : std_logic_vector(1 downto 0);
    signal VN695_in4 : std_logic_vector(1 downto 0);
    signal VN695_in5 : std_logic_vector(1 downto 0);
    signal VN696_in0 : std_logic_vector(1 downto 0);
    signal VN696_in1 : std_logic_vector(1 downto 0);
    signal VN696_in2 : std_logic_vector(1 downto 0);
    signal VN696_in3 : std_logic_vector(1 downto 0);
    signal VN696_in4 : std_logic_vector(1 downto 0);
    signal VN696_in5 : std_logic_vector(1 downto 0);
    signal VN697_in0 : std_logic_vector(1 downto 0);
    signal VN697_in1 : std_logic_vector(1 downto 0);
    signal VN697_in2 : std_logic_vector(1 downto 0);
    signal VN697_in3 : std_logic_vector(1 downto 0);
    signal VN697_in4 : std_logic_vector(1 downto 0);
    signal VN697_in5 : std_logic_vector(1 downto 0);
    signal VN698_in0 : std_logic_vector(1 downto 0);
    signal VN698_in1 : std_logic_vector(1 downto 0);
    signal VN698_in2 : std_logic_vector(1 downto 0);
    signal VN698_in3 : std_logic_vector(1 downto 0);
    signal VN698_in4 : std_logic_vector(1 downto 0);
    signal VN698_in5 : std_logic_vector(1 downto 0);
    signal VN699_in0 : std_logic_vector(1 downto 0);
    signal VN699_in1 : std_logic_vector(1 downto 0);
    signal VN699_in2 : std_logic_vector(1 downto 0);
    signal VN699_in3 : std_logic_vector(1 downto 0);
    signal VN699_in4 : std_logic_vector(1 downto 0);
    signal VN699_in5 : std_logic_vector(1 downto 0);
    signal VN700_in0 : std_logic_vector(1 downto 0);
    signal VN700_in1 : std_logic_vector(1 downto 0);
    signal VN700_in2 : std_logic_vector(1 downto 0);
    signal VN700_in3 : std_logic_vector(1 downto 0);
    signal VN700_in4 : std_logic_vector(1 downto 0);
    signal VN700_in5 : std_logic_vector(1 downto 0);
    signal VN701_in0 : std_logic_vector(1 downto 0);
    signal VN701_in1 : std_logic_vector(1 downto 0);
    signal VN701_in2 : std_logic_vector(1 downto 0);
    signal VN701_in3 : std_logic_vector(1 downto 0);
    signal VN701_in4 : std_logic_vector(1 downto 0);
    signal VN701_in5 : std_logic_vector(1 downto 0);
    signal VN702_in0 : std_logic_vector(1 downto 0);
    signal VN702_in1 : std_logic_vector(1 downto 0);
    signal VN702_in2 : std_logic_vector(1 downto 0);
    signal VN702_in3 : std_logic_vector(1 downto 0);
    signal VN702_in4 : std_logic_vector(1 downto 0);
    signal VN702_in5 : std_logic_vector(1 downto 0);
    signal VN703_in0 : std_logic_vector(1 downto 0);
    signal VN703_in1 : std_logic_vector(1 downto 0);
    signal VN703_in2 : std_logic_vector(1 downto 0);
    signal VN703_in3 : std_logic_vector(1 downto 0);
    signal VN703_in4 : std_logic_vector(1 downto 0);
    signal VN703_in5 : std_logic_vector(1 downto 0);
    signal VN704_in0 : std_logic_vector(1 downto 0);
    signal VN704_in1 : std_logic_vector(1 downto 0);
    signal VN704_in2 : std_logic_vector(1 downto 0);
    signal VN704_in3 : std_logic_vector(1 downto 0);
    signal VN704_in4 : std_logic_vector(1 downto 0);
    signal VN704_in5 : std_logic_vector(1 downto 0);
    signal VN705_in0 : std_logic_vector(1 downto 0);
    signal VN705_in1 : std_logic_vector(1 downto 0);
    signal VN705_in2 : std_logic_vector(1 downto 0);
    signal VN705_in3 : std_logic_vector(1 downto 0);
    signal VN705_in4 : std_logic_vector(1 downto 0);
    signal VN705_in5 : std_logic_vector(1 downto 0);
    signal VN706_in0 : std_logic_vector(1 downto 0);
    signal VN706_in1 : std_logic_vector(1 downto 0);
    signal VN706_in2 : std_logic_vector(1 downto 0);
    signal VN706_in3 : std_logic_vector(1 downto 0);
    signal VN706_in4 : std_logic_vector(1 downto 0);
    signal VN706_in5 : std_logic_vector(1 downto 0);
    signal VN707_in0 : std_logic_vector(1 downto 0);
    signal VN707_in1 : std_logic_vector(1 downto 0);
    signal VN707_in2 : std_logic_vector(1 downto 0);
    signal VN707_in3 : std_logic_vector(1 downto 0);
    signal VN707_in4 : std_logic_vector(1 downto 0);
    signal VN707_in5 : std_logic_vector(1 downto 0);
    signal VN708_in0 : std_logic_vector(1 downto 0);
    signal VN708_in1 : std_logic_vector(1 downto 0);
    signal VN708_in2 : std_logic_vector(1 downto 0);
    signal VN708_in3 : std_logic_vector(1 downto 0);
    signal VN708_in4 : std_logic_vector(1 downto 0);
    signal VN708_in5 : std_logic_vector(1 downto 0);
    signal VN709_in0 : std_logic_vector(1 downto 0);
    signal VN709_in1 : std_logic_vector(1 downto 0);
    signal VN709_in2 : std_logic_vector(1 downto 0);
    signal VN709_in3 : std_logic_vector(1 downto 0);
    signal VN709_in4 : std_logic_vector(1 downto 0);
    signal VN709_in5 : std_logic_vector(1 downto 0);
    signal VN710_in0 : std_logic_vector(1 downto 0);
    signal VN710_in1 : std_logic_vector(1 downto 0);
    signal VN710_in2 : std_logic_vector(1 downto 0);
    signal VN710_in3 : std_logic_vector(1 downto 0);
    signal VN710_in4 : std_logic_vector(1 downto 0);
    signal VN710_in5 : std_logic_vector(1 downto 0);
    signal VN711_in0 : std_logic_vector(1 downto 0);
    signal VN711_in1 : std_logic_vector(1 downto 0);
    signal VN711_in2 : std_logic_vector(1 downto 0);
    signal VN711_in3 : std_logic_vector(1 downto 0);
    signal VN711_in4 : std_logic_vector(1 downto 0);
    signal VN711_in5 : std_logic_vector(1 downto 0);
    signal VN712_in0 : std_logic_vector(1 downto 0);
    signal VN712_in1 : std_logic_vector(1 downto 0);
    signal VN712_in2 : std_logic_vector(1 downto 0);
    signal VN712_in3 : std_logic_vector(1 downto 0);
    signal VN712_in4 : std_logic_vector(1 downto 0);
    signal VN712_in5 : std_logic_vector(1 downto 0);
    signal VN713_in0 : std_logic_vector(1 downto 0);
    signal VN713_in1 : std_logic_vector(1 downto 0);
    signal VN713_in2 : std_logic_vector(1 downto 0);
    signal VN713_in3 : std_logic_vector(1 downto 0);
    signal VN713_in4 : std_logic_vector(1 downto 0);
    signal VN713_in5 : std_logic_vector(1 downto 0);
    signal VN714_in0 : std_logic_vector(1 downto 0);
    signal VN714_in1 : std_logic_vector(1 downto 0);
    signal VN714_in2 : std_logic_vector(1 downto 0);
    signal VN714_in3 : std_logic_vector(1 downto 0);
    signal VN714_in4 : std_logic_vector(1 downto 0);
    signal VN714_in5 : std_logic_vector(1 downto 0);
    signal VN715_in0 : std_logic_vector(1 downto 0);
    signal VN715_in1 : std_logic_vector(1 downto 0);
    signal VN715_in2 : std_logic_vector(1 downto 0);
    signal VN715_in3 : std_logic_vector(1 downto 0);
    signal VN715_in4 : std_logic_vector(1 downto 0);
    signal VN715_in5 : std_logic_vector(1 downto 0);
    signal VN716_in0 : std_logic_vector(1 downto 0);
    signal VN716_in1 : std_logic_vector(1 downto 0);
    signal VN716_in2 : std_logic_vector(1 downto 0);
    signal VN716_in3 : std_logic_vector(1 downto 0);
    signal VN716_in4 : std_logic_vector(1 downto 0);
    signal VN716_in5 : std_logic_vector(1 downto 0);
    signal VN717_in0 : std_logic_vector(1 downto 0);
    signal VN717_in1 : std_logic_vector(1 downto 0);
    signal VN717_in2 : std_logic_vector(1 downto 0);
    signal VN717_in3 : std_logic_vector(1 downto 0);
    signal VN717_in4 : std_logic_vector(1 downto 0);
    signal VN717_in5 : std_logic_vector(1 downto 0);
    signal VN718_in0 : std_logic_vector(1 downto 0);
    signal VN718_in1 : std_logic_vector(1 downto 0);
    signal VN718_in2 : std_logic_vector(1 downto 0);
    signal VN718_in3 : std_logic_vector(1 downto 0);
    signal VN718_in4 : std_logic_vector(1 downto 0);
    signal VN718_in5 : std_logic_vector(1 downto 0);
    signal VN719_in0 : std_logic_vector(1 downto 0);
    signal VN719_in1 : std_logic_vector(1 downto 0);
    signal VN719_in2 : std_logic_vector(1 downto 0);
    signal VN719_in3 : std_logic_vector(1 downto 0);
    signal VN719_in4 : std_logic_vector(1 downto 0);
    signal VN719_in5 : std_logic_vector(1 downto 0);
    signal VN720_in0 : std_logic_vector(1 downto 0);
    signal VN720_in1 : std_logic_vector(1 downto 0);
    signal VN720_in2 : std_logic_vector(1 downto 0);
    signal VN720_in3 : std_logic_vector(1 downto 0);
    signal VN720_in4 : std_logic_vector(1 downto 0);
    signal VN720_in5 : std_logic_vector(1 downto 0);
    signal VN721_in0 : std_logic_vector(1 downto 0);
    signal VN721_in1 : std_logic_vector(1 downto 0);
    signal VN721_in2 : std_logic_vector(1 downto 0);
    signal VN721_in3 : std_logic_vector(1 downto 0);
    signal VN721_in4 : std_logic_vector(1 downto 0);
    signal VN721_in5 : std_logic_vector(1 downto 0);
    signal VN722_in0 : std_logic_vector(1 downto 0);
    signal VN722_in1 : std_logic_vector(1 downto 0);
    signal VN722_in2 : std_logic_vector(1 downto 0);
    signal VN722_in3 : std_logic_vector(1 downto 0);
    signal VN722_in4 : std_logic_vector(1 downto 0);
    signal VN722_in5 : std_logic_vector(1 downto 0);
    signal VN723_in0 : std_logic_vector(1 downto 0);
    signal VN723_in1 : std_logic_vector(1 downto 0);
    signal VN723_in2 : std_logic_vector(1 downto 0);
    signal VN723_in3 : std_logic_vector(1 downto 0);
    signal VN723_in4 : std_logic_vector(1 downto 0);
    signal VN723_in5 : std_logic_vector(1 downto 0);
    signal VN724_in0 : std_logic_vector(1 downto 0);
    signal VN724_in1 : std_logic_vector(1 downto 0);
    signal VN724_in2 : std_logic_vector(1 downto 0);
    signal VN724_in3 : std_logic_vector(1 downto 0);
    signal VN724_in4 : std_logic_vector(1 downto 0);
    signal VN724_in5 : std_logic_vector(1 downto 0);
    signal VN725_in0 : std_logic_vector(1 downto 0);
    signal VN725_in1 : std_logic_vector(1 downto 0);
    signal VN725_in2 : std_logic_vector(1 downto 0);
    signal VN725_in3 : std_logic_vector(1 downto 0);
    signal VN725_in4 : std_logic_vector(1 downto 0);
    signal VN725_in5 : std_logic_vector(1 downto 0);
    signal VN726_in0 : std_logic_vector(1 downto 0);
    signal VN726_in1 : std_logic_vector(1 downto 0);
    signal VN726_in2 : std_logic_vector(1 downto 0);
    signal VN726_in3 : std_logic_vector(1 downto 0);
    signal VN726_in4 : std_logic_vector(1 downto 0);
    signal VN726_in5 : std_logic_vector(1 downto 0);
    signal VN727_in0 : std_logic_vector(1 downto 0);
    signal VN727_in1 : std_logic_vector(1 downto 0);
    signal VN727_in2 : std_logic_vector(1 downto 0);
    signal VN727_in3 : std_logic_vector(1 downto 0);
    signal VN727_in4 : std_logic_vector(1 downto 0);
    signal VN727_in5 : std_logic_vector(1 downto 0);
    signal VN728_in0 : std_logic_vector(1 downto 0);
    signal VN728_in1 : std_logic_vector(1 downto 0);
    signal VN728_in2 : std_logic_vector(1 downto 0);
    signal VN728_in3 : std_logic_vector(1 downto 0);
    signal VN728_in4 : std_logic_vector(1 downto 0);
    signal VN728_in5 : std_logic_vector(1 downto 0);
    signal VN729_in0 : std_logic_vector(1 downto 0);
    signal VN729_in1 : std_logic_vector(1 downto 0);
    signal VN729_in2 : std_logic_vector(1 downto 0);
    signal VN729_in3 : std_logic_vector(1 downto 0);
    signal VN729_in4 : std_logic_vector(1 downto 0);
    signal VN729_in5 : std_logic_vector(1 downto 0);
    signal VN730_in0 : std_logic_vector(1 downto 0);
    signal VN730_in1 : std_logic_vector(1 downto 0);
    signal VN730_in2 : std_logic_vector(1 downto 0);
    signal VN730_in3 : std_logic_vector(1 downto 0);
    signal VN730_in4 : std_logic_vector(1 downto 0);
    signal VN730_in5 : std_logic_vector(1 downto 0);
    signal VN731_in0 : std_logic_vector(1 downto 0);
    signal VN731_in1 : std_logic_vector(1 downto 0);
    signal VN731_in2 : std_logic_vector(1 downto 0);
    signal VN731_in3 : std_logic_vector(1 downto 0);
    signal VN731_in4 : std_logic_vector(1 downto 0);
    signal VN731_in5 : std_logic_vector(1 downto 0);
    signal VN732_in0 : std_logic_vector(1 downto 0);
    signal VN732_in1 : std_logic_vector(1 downto 0);
    signal VN732_in2 : std_logic_vector(1 downto 0);
    signal VN732_in3 : std_logic_vector(1 downto 0);
    signal VN732_in4 : std_logic_vector(1 downto 0);
    signal VN732_in5 : std_logic_vector(1 downto 0);
    signal VN733_in0 : std_logic_vector(1 downto 0);
    signal VN733_in1 : std_logic_vector(1 downto 0);
    signal VN733_in2 : std_logic_vector(1 downto 0);
    signal VN733_in3 : std_logic_vector(1 downto 0);
    signal VN733_in4 : std_logic_vector(1 downto 0);
    signal VN733_in5 : std_logic_vector(1 downto 0);
    signal VN734_in0 : std_logic_vector(1 downto 0);
    signal VN734_in1 : std_logic_vector(1 downto 0);
    signal VN734_in2 : std_logic_vector(1 downto 0);
    signal VN734_in3 : std_logic_vector(1 downto 0);
    signal VN734_in4 : std_logic_vector(1 downto 0);
    signal VN734_in5 : std_logic_vector(1 downto 0);
    signal VN735_in0 : std_logic_vector(1 downto 0);
    signal VN735_in1 : std_logic_vector(1 downto 0);
    signal VN735_in2 : std_logic_vector(1 downto 0);
    signal VN735_in3 : std_logic_vector(1 downto 0);
    signal VN735_in4 : std_logic_vector(1 downto 0);
    signal VN735_in5 : std_logic_vector(1 downto 0);
    signal VN736_in0 : std_logic_vector(1 downto 0);
    signal VN736_in1 : std_logic_vector(1 downto 0);
    signal VN736_in2 : std_logic_vector(1 downto 0);
    signal VN736_in3 : std_logic_vector(1 downto 0);
    signal VN736_in4 : std_logic_vector(1 downto 0);
    signal VN736_in5 : std_logic_vector(1 downto 0);
    signal VN737_in0 : std_logic_vector(1 downto 0);
    signal VN737_in1 : std_logic_vector(1 downto 0);
    signal VN737_in2 : std_logic_vector(1 downto 0);
    signal VN737_in3 : std_logic_vector(1 downto 0);
    signal VN737_in4 : std_logic_vector(1 downto 0);
    signal VN737_in5 : std_logic_vector(1 downto 0);
    signal VN738_in0 : std_logic_vector(1 downto 0);
    signal VN738_in1 : std_logic_vector(1 downto 0);
    signal VN738_in2 : std_logic_vector(1 downto 0);
    signal VN738_in3 : std_logic_vector(1 downto 0);
    signal VN738_in4 : std_logic_vector(1 downto 0);
    signal VN738_in5 : std_logic_vector(1 downto 0);
    signal VN739_in0 : std_logic_vector(1 downto 0);
    signal VN739_in1 : std_logic_vector(1 downto 0);
    signal VN739_in2 : std_logic_vector(1 downto 0);
    signal VN739_in3 : std_logic_vector(1 downto 0);
    signal VN739_in4 : std_logic_vector(1 downto 0);
    signal VN739_in5 : std_logic_vector(1 downto 0);
    signal VN740_in0 : std_logic_vector(1 downto 0);
    signal VN740_in1 : std_logic_vector(1 downto 0);
    signal VN740_in2 : std_logic_vector(1 downto 0);
    signal VN740_in3 : std_logic_vector(1 downto 0);
    signal VN740_in4 : std_logic_vector(1 downto 0);
    signal VN740_in5 : std_logic_vector(1 downto 0);
    signal VN741_in0 : std_logic_vector(1 downto 0);
    signal VN741_in1 : std_logic_vector(1 downto 0);
    signal VN741_in2 : std_logic_vector(1 downto 0);
    signal VN741_in3 : std_logic_vector(1 downto 0);
    signal VN741_in4 : std_logic_vector(1 downto 0);
    signal VN741_in5 : std_logic_vector(1 downto 0);
    signal VN742_in0 : std_logic_vector(1 downto 0);
    signal VN742_in1 : std_logic_vector(1 downto 0);
    signal VN742_in2 : std_logic_vector(1 downto 0);
    signal VN742_in3 : std_logic_vector(1 downto 0);
    signal VN742_in4 : std_logic_vector(1 downto 0);
    signal VN742_in5 : std_logic_vector(1 downto 0);
    signal VN743_in0 : std_logic_vector(1 downto 0);
    signal VN743_in1 : std_logic_vector(1 downto 0);
    signal VN743_in2 : std_logic_vector(1 downto 0);
    signal VN743_in3 : std_logic_vector(1 downto 0);
    signal VN743_in4 : std_logic_vector(1 downto 0);
    signal VN743_in5 : std_logic_vector(1 downto 0);
    signal VN744_in0 : std_logic_vector(1 downto 0);
    signal VN744_in1 : std_logic_vector(1 downto 0);
    signal VN744_in2 : std_logic_vector(1 downto 0);
    signal VN744_in3 : std_logic_vector(1 downto 0);
    signal VN744_in4 : std_logic_vector(1 downto 0);
    signal VN744_in5 : std_logic_vector(1 downto 0);
    signal VN745_in0 : std_logic_vector(1 downto 0);
    signal VN745_in1 : std_logic_vector(1 downto 0);
    signal VN745_in2 : std_logic_vector(1 downto 0);
    signal VN745_in3 : std_logic_vector(1 downto 0);
    signal VN745_in4 : std_logic_vector(1 downto 0);
    signal VN745_in5 : std_logic_vector(1 downto 0);
    signal VN746_in0 : std_logic_vector(1 downto 0);
    signal VN746_in1 : std_logic_vector(1 downto 0);
    signal VN746_in2 : std_logic_vector(1 downto 0);
    signal VN746_in3 : std_logic_vector(1 downto 0);
    signal VN746_in4 : std_logic_vector(1 downto 0);
    signal VN746_in5 : std_logic_vector(1 downto 0);
    signal VN747_in0 : std_logic_vector(1 downto 0);
    signal VN747_in1 : std_logic_vector(1 downto 0);
    signal VN747_in2 : std_logic_vector(1 downto 0);
    signal VN747_in3 : std_logic_vector(1 downto 0);
    signal VN747_in4 : std_logic_vector(1 downto 0);
    signal VN747_in5 : std_logic_vector(1 downto 0);
    signal VN748_in0 : std_logic_vector(1 downto 0);
    signal VN748_in1 : std_logic_vector(1 downto 0);
    signal VN748_in2 : std_logic_vector(1 downto 0);
    signal VN748_in3 : std_logic_vector(1 downto 0);
    signal VN748_in4 : std_logic_vector(1 downto 0);
    signal VN748_in5 : std_logic_vector(1 downto 0);
    signal VN749_in0 : std_logic_vector(1 downto 0);
    signal VN749_in1 : std_logic_vector(1 downto 0);
    signal VN749_in2 : std_logic_vector(1 downto 0);
    signal VN749_in3 : std_logic_vector(1 downto 0);
    signal VN749_in4 : std_logic_vector(1 downto 0);
    signal VN749_in5 : std_logic_vector(1 downto 0);
    signal VN750_in0 : std_logic_vector(1 downto 0);
    signal VN750_in1 : std_logic_vector(1 downto 0);
    signal VN750_in2 : std_logic_vector(1 downto 0);
    signal VN750_in3 : std_logic_vector(1 downto 0);
    signal VN750_in4 : std_logic_vector(1 downto 0);
    signal VN750_in5 : std_logic_vector(1 downto 0);
    signal VN751_in0 : std_logic_vector(1 downto 0);
    signal VN751_in1 : std_logic_vector(1 downto 0);
    signal VN751_in2 : std_logic_vector(1 downto 0);
    signal VN751_in3 : std_logic_vector(1 downto 0);
    signal VN751_in4 : std_logic_vector(1 downto 0);
    signal VN751_in5 : std_logic_vector(1 downto 0);
    signal VN752_in0 : std_logic_vector(1 downto 0);
    signal VN752_in1 : std_logic_vector(1 downto 0);
    signal VN752_in2 : std_logic_vector(1 downto 0);
    signal VN752_in3 : std_logic_vector(1 downto 0);
    signal VN752_in4 : std_logic_vector(1 downto 0);
    signal VN752_in5 : std_logic_vector(1 downto 0);
    signal VN753_in0 : std_logic_vector(1 downto 0);
    signal VN753_in1 : std_logic_vector(1 downto 0);
    signal VN753_in2 : std_logic_vector(1 downto 0);
    signal VN753_in3 : std_logic_vector(1 downto 0);
    signal VN753_in4 : std_logic_vector(1 downto 0);
    signal VN753_in5 : std_logic_vector(1 downto 0);
    signal VN754_in0 : std_logic_vector(1 downto 0);
    signal VN754_in1 : std_logic_vector(1 downto 0);
    signal VN754_in2 : std_logic_vector(1 downto 0);
    signal VN754_in3 : std_logic_vector(1 downto 0);
    signal VN754_in4 : std_logic_vector(1 downto 0);
    signal VN754_in5 : std_logic_vector(1 downto 0);
    signal VN755_in0 : std_logic_vector(1 downto 0);
    signal VN755_in1 : std_logic_vector(1 downto 0);
    signal VN755_in2 : std_logic_vector(1 downto 0);
    signal VN755_in3 : std_logic_vector(1 downto 0);
    signal VN755_in4 : std_logic_vector(1 downto 0);
    signal VN755_in5 : std_logic_vector(1 downto 0);
    signal VN756_in0 : std_logic_vector(1 downto 0);
    signal VN756_in1 : std_logic_vector(1 downto 0);
    signal VN756_in2 : std_logic_vector(1 downto 0);
    signal VN756_in3 : std_logic_vector(1 downto 0);
    signal VN756_in4 : std_logic_vector(1 downto 0);
    signal VN756_in5 : std_logic_vector(1 downto 0);
    signal VN757_in0 : std_logic_vector(1 downto 0);
    signal VN757_in1 : std_logic_vector(1 downto 0);
    signal VN757_in2 : std_logic_vector(1 downto 0);
    signal VN757_in3 : std_logic_vector(1 downto 0);
    signal VN757_in4 : std_logic_vector(1 downto 0);
    signal VN757_in5 : std_logic_vector(1 downto 0);
    signal VN758_in0 : std_logic_vector(1 downto 0);
    signal VN758_in1 : std_logic_vector(1 downto 0);
    signal VN758_in2 : std_logic_vector(1 downto 0);
    signal VN758_in3 : std_logic_vector(1 downto 0);
    signal VN758_in4 : std_logic_vector(1 downto 0);
    signal VN758_in5 : std_logic_vector(1 downto 0);
    signal VN759_in0 : std_logic_vector(1 downto 0);
    signal VN759_in1 : std_logic_vector(1 downto 0);
    signal VN759_in2 : std_logic_vector(1 downto 0);
    signal VN759_in3 : std_logic_vector(1 downto 0);
    signal VN759_in4 : std_logic_vector(1 downto 0);
    signal VN759_in5 : std_logic_vector(1 downto 0);
    signal VN760_in0 : std_logic_vector(1 downto 0);
    signal VN760_in1 : std_logic_vector(1 downto 0);
    signal VN760_in2 : std_logic_vector(1 downto 0);
    signal VN760_in3 : std_logic_vector(1 downto 0);
    signal VN760_in4 : std_logic_vector(1 downto 0);
    signal VN760_in5 : std_logic_vector(1 downto 0);
    signal VN761_in0 : std_logic_vector(1 downto 0);
    signal VN761_in1 : std_logic_vector(1 downto 0);
    signal VN761_in2 : std_logic_vector(1 downto 0);
    signal VN761_in3 : std_logic_vector(1 downto 0);
    signal VN761_in4 : std_logic_vector(1 downto 0);
    signal VN761_in5 : std_logic_vector(1 downto 0);
    signal VN762_in0 : std_logic_vector(1 downto 0);
    signal VN762_in1 : std_logic_vector(1 downto 0);
    signal VN762_in2 : std_logic_vector(1 downto 0);
    signal VN762_in3 : std_logic_vector(1 downto 0);
    signal VN762_in4 : std_logic_vector(1 downto 0);
    signal VN762_in5 : std_logic_vector(1 downto 0);
    signal VN763_in0 : std_logic_vector(1 downto 0);
    signal VN763_in1 : std_logic_vector(1 downto 0);
    signal VN763_in2 : std_logic_vector(1 downto 0);
    signal VN763_in3 : std_logic_vector(1 downto 0);
    signal VN763_in4 : std_logic_vector(1 downto 0);
    signal VN763_in5 : std_logic_vector(1 downto 0);
    signal VN764_in0 : std_logic_vector(1 downto 0);
    signal VN764_in1 : std_logic_vector(1 downto 0);
    signal VN764_in2 : std_logic_vector(1 downto 0);
    signal VN764_in3 : std_logic_vector(1 downto 0);
    signal VN764_in4 : std_logic_vector(1 downto 0);
    signal VN764_in5 : std_logic_vector(1 downto 0);
    signal VN765_in0 : std_logic_vector(1 downto 0);
    signal VN765_in1 : std_logic_vector(1 downto 0);
    signal VN765_in2 : std_logic_vector(1 downto 0);
    signal VN765_in3 : std_logic_vector(1 downto 0);
    signal VN765_in4 : std_logic_vector(1 downto 0);
    signal VN765_in5 : std_logic_vector(1 downto 0);
    signal VN766_in0 : std_logic_vector(1 downto 0);
    signal VN766_in1 : std_logic_vector(1 downto 0);
    signal VN766_in2 : std_logic_vector(1 downto 0);
    signal VN766_in3 : std_logic_vector(1 downto 0);
    signal VN766_in4 : std_logic_vector(1 downto 0);
    signal VN766_in5 : std_logic_vector(1 downto 0);
    signal VN767_in0 : std_logic_vector(1 downto 0);
    signal VN767_in1 : std_logic_vector(1 downto 0);
    signal VN767_in2 : std_logic_vector(1 downto 0);
    signal VN767_in3 : std_logic_vector(1 downto 0);
    signal VN767_in4 : std_logic_vector(1 downto 0);
    signal VN767_in5 : std_logic_vector(1 downto 0);
    signal VN768_in0 : std_logic_vector(1 downto 0);
    signal VN768_in1 : std_logic_vector(1 downto 0);
    signal VN768_in2 : std_logic_vector(1 downto 0);
    signal VN768_in3 : std_logic_vector(1 downto 0);
    signal VN768_in4 : std_logic_vector(1 downto 0);
    signal VN768_in5 : std_logic_vector(1 downto 0);
    signal VN769_in0 : std_logic_vector(1 downto 0);
    signal VN769_in1 : std_logic_vector(1 downto 0);
    signal VN769_in2 : std_logic_vector(1 downto 0);
    signal VN769_in3 : std_logic_vector(1 downto 0);
    signal VN769_in4 : std_logic_vector(1 downto 0);
    signal VN769_in5 : std_logic_vector(1 downto 0);
    signal VN770_in0 : std_logic_vector(1 downto 0);
    signal VN770_in1 : std_logic_vector(1 downto 0);
    signal VN770_in2 : std_logic_vector(1 downto 0);
    signal VN770_in3 : std_logic_vector(1 downto 0);
    signal VN770_in4 : std_logic_vector(1 downto 0);
    signal VN770_in5 : std_logic_vector(1 downto 0);
    signal VN771_in0 : std_logic_vector(1 downto 0);
    signal VN771_in1 : std_logic_vector(1 downto 0);
    signal VN771_in2 : std_logic_vector(1 downto 0);
    signal VN771_in3 : std_logic_vector(1 downto 0);
    signal VN771_in4 : std_logic_vector(1 downto 0);
    signal VN771_in5 : std_logic_vector(1 downto 0);
    signal VN772_in0 : std_logic_vector(1 downto 0);
    signal VN772_in1 : std_logic_vector(1 downto 0);
    signal VN772_in2 : std_logic_vector(1 downto 0);
    signal VN772_in3 : std_logic_vector(1 downto 0);
    signal VN772_in4 : std_logic_vector(1 downto 0);
    signal VN772_in5 : std_logic_vector(1 downto 0);
    signal VN773_in0 : std_logic_vector(1 downto 0);
    signal VN773_in1 : std_logic_vector(1 downto 0);
    signal VN773_in2 : std_logic_vector(1 downto 0);
    signal VN773_in3 : std_logic_vector(1 downto 0);
    signal VN773_in4 : std_logic_vector(1 downto 0);
    signal VN773_in5 : std_logic_vector(1 downto 0);
    signal VN774_in0 : std_logic_vector(1 downto 0);
    signal VN774_in1 : std_logic_vector(1 downto 0);
    signal VN774_in2 : std_logic_vector(1 downto 0);
    signal VN774_in3 : std_logic_vector(1 downto 0);
    signal VN774_in4 : std_logic_vector(1 downto 0);
    signal VN774_in5 : std_logic_vector(1 downto 0);
    signal VN775_in0 : std_logic_vector(1 downto 0);
    signal VN775_in1 : std_logic_vector(1 downto 0);
    signal VN775_in2 : std_logic_vector(1 downto 0);
    signal VN775_in3 : std_logic_vector(1 downto 0);
    signal VN775_in4 : std_logic_vector(1 downto 0);
    signal VN775_in5 : std_logic_vector(1 downto 0);
    signal VN776_in0 : std_logic_vector(1 downto 0);
    signal VN776_in1 : std_logic_vector(1 downto 0);
    signal VN776_in2 : std_logic_vector(1 downto 0);
    signal VN776_in3 : std_logic_vector(1 downto 0);
    signal VN776_in4 : std_logic_vector(1 downto 0);
    signal VN776_in5 : std_logic_vector(1 downto 0);
    signal VN777_in0 : std_logic_vector(1 downto 0);
    signal VN777_in1 : std_logic_vector(1 downto 0);
    signal VN777_in2 : std_logic_vector(1 downto 0);
    signal VN777_in3 : std_logic_vector(1 downto 0);
    signal VN777_in4 : std_logic_vector(1 downto 0);
    signal VN777_in5 : std_logic_vector(1 downto 0);
    signal VN778_in0 : std_logic_vector(1 downto 0);
    signal VN778_in1 : std_logic_vector(1 downto 0);
    signal VN778_in2 : std_logic_vector(1 downto 0);
    signal VN778_in3 : std_logic_vector(1 downto 0);
    signal VN778_in4 : std_logic_vector(1 downto 0);
    signal VN778_in5 : std_logic_vector(1 downto 0);
    signal VN779_in0 : std_logic_vector(1 downto 0);
    signal VN779_in1 : std_logic_vector(1 downto 0);
    signal VN779_in2 : std_logic_vector(1 downto 0);
    signal VN779_in3 : std_logic_vector(1 downto 0);
    signal VN779_in4 : std_logic_vector(1 downto 0);
    signal VN779_in5 : std_logic_vector(1 downto 0);
    signal VN780_in0 : std_logic_vector(1 downto 0);
    signal VN780_in1 : std_logic_vector(1 downto 0);
    signal VN780_in2 : std_logic_vector(1 downto 0);
    signal VN780_in3 : std_logic_vector(1 downto 0);
    signal VN780_in4 : std_logic_vector(1 downto 0);
    signal VN780_in5 : std_logic_vector(1 downto 0);
    signal VN781_in0 : std_logic_vector(1 downto 0);
    signal VN781_in1 : std_logic_vector(1 downto 0);
    signal VN781_in2 : std_logic_vector(1 downto 0);
    signal VN781_in3 : std_logic_vector(1 downto 0);
    signal VN781_in4 : std_logic_vector(1 downto 0);
    signal VN781_in5 : std_logic_vector(1 downto 0);
    signal VN782_in0 : std_logic_vector(1 downto 0);
    signal VN782_in1 : std_logic_vector(1 downto 0);
    signal VN782_in2 : std_logic_vector(1 downto 0);
    signal VN782_in3 : std_logic_vector(1 downto 0);
    signal VN782_in4 : std_logic_vector(1 downto 0);
    signal VN782_in5 : std_logic_vector(1 downto 0);
    signal VN783_in0 : std_logic_vector(1 downto 0);
    signal VN783_in1 : std_logic_vector(1 downto 0);
    signal VN783_in2 : std_logic_vector(1 downto 0);
    signal VN783_in3 : std_logic_vector(1 downto 0);
    signal VN783_in4 : std_logic_vector(1 downto 0);
    signal VN783_in5 : std_logic_vector(1 downto 0);
    signal VN784_in0 : std_logic_vector(1 downto 0);
    signal VN784_in1 : std_logic_vector(1 downto 0);
    signal VN784_in2 : std_logic_vector(1 downto 0);
    signal VN784_in3 : std_logic_vector(1 downto 0);
    signal VN784_in4 : std_logic_vector(1 downto 0);
    signal VN784_in5 : std_logic_vector(1 downto 0);
    signal VN785_in0 : std_logic_vector(1 downto 0);
    signal VN785_in1 : std_logic_vector(1 downto 0);
    signal VN785_in2 : std_logic_vector(1 downto 0);
    signal VN785_in3 : std_logic_vector(1 downto 0);
    signal VN785_in4 : std_logic_vector(1 downto 0);
    signal VN785_in5 : std_logic_vector(1 downto 0);
    signal VN786_in0 : std_logic_vector(1 downto 0);
    signal VN786_in1 : std_logic_vector(1 downto 0);
    signal VN786_in2 : std_logic_vector(1 downto 0);
    signal VN786_in3 : std_logic_vector(1 downto 0);
    signal VN786_in4 : std_logic_vector(1 downto 0);
    signal VN786_in5 : std_logic_vector(1 downto 0);
    signal VN787_in0 : std_logic_vector(1 downto 0);
    signal VN787_in1 : std_logic_vector(1 downto 0);
    signal VN787_in2 : std_logic_vector(1 downto 0);
    signal VN787_in3 : std_logic_vector(1 downto 0);
    signal VN787_in4 : std_logic_vector(1 downto 0);
    signal VN787_in5 : std_logic_vector(1 downto 0);
    signal VN788_in0 : std_logic_vector(1 downto 0);
    signal VN788_in1 : std_logic_vector(1 downto 0);
    signal VN788_in2 : std_logic_vector(1 downto 0);
    signal VN788_in3 : std_logic_vector(1 downto 0);
    signal VN788_in4 : std_logic_vector(1 downto 0);
    signal VN788_in5 : std_logic_vector(1 downto 0);
    signal VN789_in0 : std_logic_vector(1 downto 0);
    signal VN789_in1 : std_logic_vector(1 downto 0);
    signal VN789_in2 : std_logic_vector(1 downto 0);
    signal VN789_in3 : std_logic_vector(1 downto 0);
    signal VN789_in4 : std_logic_vector(1 downto 0);
    signal VN789_in5 : std_logic_vector(1 downto 0);
    signal VN790_in0 : std_logic_vector(1 downto 0);
    signal VN790_in1 : std_logic_vector(1 downto 0);
    signal VN790_in2 : std_logic_vector(1 downto 0);
    signal VN790_in3 : std_logic_vector(1 downto 0);
    signal VN790_in4 : std_logic_vector(1 downto 0);
    signal VN790_in5 : std_logic_vector(1 downto 0);
    signal VN791_in0 : std_logic_vector(1 downto 0);
    signal VN791_in1 : std_logic_vector(1 downto 0);
    signal VN791_in2 : std_logic_vector(1 downto 0);
    signal VN791_in3 : std_logic_vector(1 downto 0);
    signal VN791_in4 : std_logic_vector(1 downto 0);
    signal VN791_in5 : std_logic_vector(1 downto 0);
    signal VN792_in0 : std_logic_vector(1 downto 0);
    signal VN792_in1 : std_logic_vector(1 downto 0);
    signal VN792_in2 : std_logic_vector(1 downto 0);
    signal VN792_in3 : std_logic_vector(1 downto 0);
    signal VN792_in4 : std_logic_vector(1 downto 0);
    signal VN792_in5 : std_logic_vector(1 downto 0);
    signal VN793_in0 : std_logic_vector(1 downto 0);
    signal VN793_in1 : std_logic_vector(1 downto 0);
    signal VN793_in2 : std_logic_vector(1 downto 0);
    signal VN793_in3 : std_logic_vector(1 downto 0);
    signal VN793_in4 : std_logic_vector(1 downto 0);
    signal VN793_in5 : std_logic_vector(1 downto 0);
    signal VN794_in0 : std_logic_vector(1 downto 0);
    signal VN794_in1 : std_logic_vector(1 downto 0);
    signal VN794_in2 : std_logic_vector(1 downto 0);
    signal VN794_in3 : std_logic_vector(1 downto 0);
    signal VN794_in4 : std_logic_vector(1 downto 0);
    signal VN794_in5 : std_logic_vector(1 downto 0);
    signal VN795_in0 : std_logic_vector(1 downto 0);
    signal VN795_in1 : std_logic_vector(1 downto 0);
    signal VN795_in2 : std_logic_vector(1 downto 0);
    signal VN795_in3 : std_logic_vector(1 downto 0);
    signal VN795_in4 : std_logic_vector(1 downto 0);
    signal VN795_in5 : std_logic_vector(1 downto 0);
    signal VN796_in0 : std_logic_vector(1 downto 0);
    signal VN796_in1 : std_logic_vector(1 downto 0);
    signal VN796_in2 : std_logic_vector(1 downto 0);
    signal VN796_in3 : std_logic_vector(1 downto 0);
    signal VN796_in4 : std_logic_vector(1 downto 0);
    signal VN796_in5 : std_logic_vector(1 downto 0);
    signal VN797_in0 : std_logic_vector(1 downto 0);
    signal VN797_in1 : std_logic_vector(1 downto 0);
    signal VN797_in2 : std_logic_vector(1 downto 0);
    signal VN797_in3 : std_logic_vector(1 downto 0);
    signal VN797_in4 : std_logic_vector(1 downto 0);
    signal VN797_in5 : std_logic_vector(1 downto 0);
    signal VN798_in0 : std_logic_vector(1 downto 0);
    signal VN798_in1 : std_logic_vector(1 downto 0);
    signal VN798_in2 : std_logic_vector(1 downto 0);
    signal VN798_in3 : std_logic_vector(1 downto 0);
    signal VN798_in4 : std_logic_vector(1 downto 0);
    signal VN798_in5 : std_logic_vector(1 downto 0);
    signal VN799_in0 : std_logic_vector(1 downto 0);
    signal VN799_in1 : std_logic_vector(1 downto 0);
    signal VN799_in2 : std_logic_vector(1 downto 0);
    signal VN799_in3 : std_logic_vector(1 downto 0);
    signal VN799_in4 : std_logic_vector(1 downto 0);
    signal VN799_in5 : std_logic_vector(1 downto 0);
    signal VN800_in0 : std_logic_vector(1 downto 0);
    signal VN800_in1 : std_logic_vector(1 downto 0);
    signal VN800_in2 : std_logic_vector(1 downto 0);
    signal VN800_in3 : std_logic_vector(1 downto 0);
    signal VN800_in4 : std_logic_vector(1 downto 0);
    signal VN800_in5 : std_logic_vector(1 downto 0);
    signal VN801_in0 : std_logic_vector(1 downto 0);
    signal VN801_in1 : std_logic_vector(1 downto 0);
    signal VN801_in2 : std_logic_vector(1 downto 0);
    signal VN801_in3 : std_logic_vector(1 downto 0);
    signal VN801_in4 : std_logic_vector(1 downto 0);
    signal VN801_in5 : std_logic_vector(1 downto 0);
    signal VN802_in0 : std_logic_vector(1 downto 0);
    signal VN802_in1 : std_logic_vector(1 downto 0);
    signal VN802_in2 : std_logic_vector(1 downto 0);
    signal VN802_in3 : std_logic_vector(1 downto 0);
    signal VN802_in4 : std_logic_vector(1 downto 0);
    signal VN802_in5 : std_logic_vector(1 downto 0);
    signal VN803_in0 : std_logic_vector(1 downto 0);
    signal VN803_in1 : std_logic_vector(1 downto 0);
    signal VN803_in2 : std_logic_vector(1 downto 0);
    signal VN803_in3 : std_logic_vector(1 downto 0);
    signal VN803_in4 : std_logic_vector(1 downto 0);
    signal VN803_in5 : std_logic_vector(1 downto 0);
    signal VN804_in0 : std_logic_vector(1 downto 0);
    signal VN804_in1 : std_logic_vector(1 downto 0);
    signal VN804_in2 : std_logic_vector(1 downto 0);
    signal VN804_in3 : std_logic_vector(1 downto 0);
    signal VN804_in4 : std_logic_vector(1 downto 0);
    signal VN804_in5 : std_logic_vector(1 downto 0);
    signal VN805_in0 : std_logic_vector(1 downto 0);
    signal VN805_in1 : std_logic_vector(1 downto 0);
    signal VN805_in2 : std_logic_vector(1 downto 0);
    signal VN805_in3 : std_logic_vector(1 downto 0);
    signal VN805_in4 : std_logic_vector(1 downto 0);
    signal VN805_in5 : std_logic_vector(1 downto 0);
    signal VN806_in0 : std_logic_vector(1 downto 0);
    signal VN806_in1 : std_logic_vector(1 downto 0);
    signal VN806_in2 : std_logic_vector(1 downto 0);
    signal VN806_in3 : std_logic_vector(1 downto 0);
    signal VN806_in4 : std_logic_vector(1 downto 0);
    signal VN806_in5 : std_logic_vector(1 downto 0);
    signal VN807_in0 : std_logic_vector(1 downto 0);
    signal VN807_in1 : std_logic_vector(1 downto 0);
    signal VN807_in2 : std_logic_vector(1 downto 0);
    signal VN807_in3 : std_logic_vector(1 downto 0);
    signal VN807_in4 : std_logic_vector(1 downto 0);
    signal VN807_in5 : std_logic_vector(1 downto 0);
    signal VN808_in0 : std_logic_vector(1 downto 0);
    signal VN808_in1 : std_logic_vector(1 downto 0);
    signal VN808_in2 : std_logic_vector(1 downto 0);
    signal VN808_in3 : std_logic_vector(1 downto 0);
    signal VN808_in4 : std_logic_vector(1 downto 0);
    signal VN808_in5 : std_logic_vector(1 downto 0);
    signal VN809_in0 : std_logic_vector(1 downto 0);
    signal VN809_in1 : std_logic_vector(1 downto 0);
    signal VN809_in2 : std_logic_vector(1 downto 0);
    signal VN809_in3 : std_logic_vector(1 downto 0);
    signal VN809_in4 : std_logic_vector(1 downto 0);
    signal VN809_in5 : std_logic_vector(1 downto 0);
    signal VN810_in0 : std_logic_vector(1 downto 0);
    signal VN810_in1 : std_logic_vector(1 downto 0);
    signal VN810_in2 : std_logic_vector(1 downto 0);
    signal VN810_in3 : std_logic_vector(1 downto 0);
    signal VN810_in4 : std_logic_vector(1 downto 0);
    signal VN810_in5 : std_logic_vector(1 downto 0);
    signal VN811_in0 : std_logic_vector(1 downto 0);
    signal VN811_in1 : std_logic_vector(1 downto 0);
    signal VN811_in2 : std_logic_vector(1 downto 0);
    signal VN811_in3 : std_logic_vector(1 downto 0);
    signal VN811_in4 : std_logic_vector(1 downto 0);
    signal VN811_in5 : std_logic_vector(1 downto 0);
    signal VN812_in0 : std_logic_vector(1 downto 0);
    signal VN812_in1 : std_logic_vector(1 downto 0);
    signal VN812_in2 : std_logic_vector(1 downto 0);
    signal VN812_in3 : std_logic_vector(1 downto 0);
    signal VN812_in4 : std_logic_vector(1 downto 0);
    signal VN812_in5 : std_logic_vector(1 downto 0);
    signal VN813_in0 : std_logic_vector(1 downto 0);
    signal VN813_in1 : std_logic_vector(1 downto 0);
    signal VN813_in2 : std_logic_vector(1 downto 0);
    signal VN813_in3 : std_logic_vector(1 downto 0);
    signal VN813_in4 : std_logic_vector(1 downto 0);
    signal VN813_in5 : std_logic_vector(1 downto 0);
    signal VN814_in0 : std_logic_vector(1 downto 0);
    signal VN814_in1 : std_logic_vector(1 downto 0);
    signal VN814_in2 : std_logic_vector(1 downto 0);
    signal VN814_in3 : std_logic_vector(1 downto 0);
    signal VN814_in4 : std_logic_vector(1 downto 0);
    signal VN814_in5 : std_logic_vector(1 downto 0);
    signal VN815_in0 : std_logic_vector(1 downto 0);
    signal VN815_in1 : std_logic_vector(1 downto 0);
    signal VN815_in2 : std_logic_vector(1 downto 0);
    signal VN815_in3 : std_logic_vector(1 downto 0);
    signal VN815_in4 : std_logic_vector(1 downto 0);
    signal VN815_in5 : std_logic_vector(1 downto 0);
    signal VN816_in0 : std_logic_vector(1 downto 0);
    signal VN816_in1 : std_logic_vector(1 downto 0);
    signal VN816_in2 : std_logic_vector(1 downto 0);
    signal VN816_in3 : std_logic_vector(1 downto 0);
    signal VN816_in4 : std_logic_vector(1 downto 0);
    signal VN816_in5 : std_logic_vector(1 downto 0);
    signal VN817_in0 : std_logic_vector(1 downto 0);
    signal VN817_in1 : std_logic_vector(1 downto 0);
    signal VN817_in2 : std_logic_vector(1 downto 0);
    signal VN817_in3 : std_logic_vector(1 downto 0);
    signal VN817_in4 : std_logic_vector(1 downto 0);
    signal VN817_in5 : std_logic_vector(1 downto 0);
    signal VN818_in0 : std_logic_vector(1 downto 0);
    signal VN818_in1 : std_logic_vector(1 downto 0);
    signal VN818_in2 : std_logic_vector(1 downto 0);
    signal VN818_in3 : std_logic_vector(1 downto 0);
    signal VN818_in4 : std_logic_vector(1 downto 0);
    signal VN818_in5 : std_logic_vector(1 downto 0);
    signal VN819_in0 : std_logic_vector(1 downto 0);
    signal VN819_in1 : std_logic_vector(1 downto 0);
    signal VN819_in2 : std_logic_vector(1 downto 0);
    signal VN819_in3 : std_logic_vector(1 downto 0);
    signal VN819_in4 : std_logic_vector(1 downto 0);
    signal VN819_in5 : std_logic_vector(1 downto 0);
    signal VN820_in0 : std_logic_vector(1 downto 0);
    signal VN820_in1 : std_logic_vector(1 downto 0);
    signal VN820_in2 : std_logic_vector(1 downto 0);
    signal VN820_in3 : std_logic_vector(1 downto 0);
    signal VN820_in4 : std_logic_vector(1 downto 0);
    signal VN820_in5 : std_logic_vector(1 downto 0);
    signal VN821_in0 : std_logic_vector(1 downto 0);
    signal VN821_in1 : std_logic_vector(1 downto 0);
    signal VN821_in2 : std_logic_vector(1 downto 0);
    signal VN821_in3 : std_logic_vector(1 downto 0);
    signal VN821_in4 : std_logic_vector(1 downto 0);
    signal VN821_in5 : std_logic_vector(1 downto 0);
    signal VN822_in0 : std_logic_vector(1 downto 0);
    signal VN822_in1 : std_logic_vector(1 downto 0);
    signal VN822_in2 : std_logic_vector(1 downto 0);
    signal VN822_in3 : std_logic_vector(1 downto 0);
    signal VN822_in4 : std_logic_vector(1 downto 0);
    signal VN822_in5 : std_logic_vector(1 downto 0);
    signal VN823_in0 : std_logic_vector(1 downto 0);
    signal VN823_in1 : std_logic_vector(1 downto 0);
    signal VN823_in2 : std_logic_vector(1 downto 0);
    signal VN823_in3 : std_logic_vector(1 downto 0);
    signal VN823_in4 : std_logic_vector(1 downto 0);
    signal VN823_in5 : std_logic_vector(1 downto 0);
    signal VN824_in0 : std_logic_vector(1 downto 0);
    signal VN824_in1 : std_logic_vector(1 downto 0);
    signal VN824_in2 : std_logic_vector(1 downto 0);
    signal VN824_in3 : std_logic_vector(1 downto 0);
    signal VN824_in4 : std_logic_vector(1 downto 0);
    signal VN824_in5 : std_logic_vector(1 downto 0);
    signal VN825_in0 : std_logic_vector(1 downto 0);
    signal VN825_in1 : std_logic_vector(1 downto 0);
    signal VN825_in2 : std_logic_vector(1 downto 0);
    signal VN825_in3 : std_logic_vector(1 downto 0);
    signal VN825_in4 : std_logic_vector(1 downto 0);
    signal VN825_in5 : std_logic_vector(1 downto 0);
    signal VN826_in0 : std_logic_vector(1 downto 0);
    signal VN826_in1 : std_logic_vector(1 downto 0);
    signal VN826_in2 : std_logic_vector(1 downto 0);
    signal VN826_in3 : std_logic_vector(1 downto 0);
    signal VN826_in4 : std_logic_vector(1 downto 0);
    signal VN826_in5 : std_logic_vector(1 downto 0);
    signal VN827_in0 : std_logic_vector(1 downto 0);
    signal VN827_in1 : std_logic_vector(1 downto 0);
    signal VN827_in2 : std_logic_vector(1 downto 0);
    signal VN827_in3 : std_logic_vector(1 downto 0);
    signal VN827_in4 : std_logic_vector(1 downto 0);
    signal VN827_in5 : std_logic_vector(1 downto 0);
    signal VN828_in0 : std_logic_vector(1 downto 0);
    signal VN828_in1 : std_logic_vector(1 downto 0);
    signal VN828_in2 : std_logic_vector(1 downto 0);
    signal VN828_in3 : std_logic_vector(1 downto 0);
    signal VN828_in4 : std_logic_vector(1 downto 0);
    signal VN828_in5 : std_logic_vector(1 downto 0);
    signal VN829_in0 : std_logic_vector(1 downto 0);
    signal VN829_in1 : std_logic_vector(1 downto 0);
    signal VN829_in2 : std_logic_vector(1 downto 0);
    signal VN829_in3 : std_logic_vector(1 downto 0);
    signal VN829_in4 : std_logic_vector(1 downto 0);
    signal VN829_in5 : std_logic_vector(1 downto 0);
    signal VN830_in0 : std_logic_vector(1 downto 0);
    signal VN830_in1 : std_logic_vector(1 downto 0);
    signal VN830_in2 : std_logic_vector(1 downto 0);
    signal VN830_in3 : std_logic_vector(1 downto 0);
    signal VN830_in4 : std_logic_vector(1 downto 0);
    signal VN830_in5 : std_logic_vector(1 downto 0);
    signal VN831_in0 : std_logic_vector(1 downto 0);
    signal VN831_in1 : std_logic_vector(1 downto 0);
    signal VN831_in2 : std_logic_vector(1 downto 0);
    signal VN831_in3 : std_logic_vector(1 downto 0);
    signal VN831_in4 : std_logic_vector(1 downto 0);
    signal VN831_in5 : std_logic_vector(1 downto 0);
    signal VN832_in0 : std_logic_vector(1 downto 0);
    signal VN832_in1 : std_logic_vector(1 downto 0);
    signal VN832_in2 : std_logic_vector(1 downto 0);
    signal VN832_in3 : std_logic_vector(1 downto 0);
    signal VN832_in4 : std_logic_vector(1 downto 0);
    signal VN832_in5 : std_logic_vector(1 downto 0);
    signal VN833_in0 : std_logic_vector(1 downto 0);
    signal VN833_in1 : std_logic_vector(1 downto 0);
    signal VN833_in2 : std_logic_vector(1 downto 0);
    signal VN833_in3 : std_logic_vector(1 downto 0);
    signal VN833_in4 : std_logic_vector(1 downto 0);
    signal VN833_in5 : std_logic_vector(1 downto 0);
    signal VN834_in0 : std_logic_vector(1 downto 0);
    signal VN834_in1 : std_logic_vector(1 downto 0);
    signal VN834_in2 : std_logic_vector(1 downto 0);
    signal VN834_in3 : std_logic_vector(1 downto 0);
    signal VN834_in4 : std_logic_vector(1 downto 0);
    signal VN834_in5 : std_logic_vector(1 downto 0);
    signal VN835_in0 : std_logic_vector(1 downto 0);
    signal VN835_in1 : std_logic_vector(1 downto 0);
    signal VN835_in2 : std_logic_vector(1 downto 0);
    signal VN835_in3 : std_logic_vector(1 downto 0);
    signal VN835_in4 : std_logic_vector(1 downto 0);
    signal VN835_in5 : std_logic_vector(1 downto 0);
    signal VN836_in0 : std_logic_vector(1 downto 0);
    signal VN836_in1 : std_logic_vector(1 downto 0);
    signal VN836_in2 : std_logic_vector(1 downto 0);
    signal VN836_in3 : std_logic_vector(1 downto 0);
    signal VN836_in4 : std_logic_vector(1 downto 0);
    signal VN836_in5 : std_logic_vector(1 downto 0);
    signal VN837_in0 : std_logic_vector(1 downto 0);
    signal VN837_in1 : std_logic_vector(1 downto 0);
    signal VN837_in2 : std_logic_vector(1 downto 0);
    signal VN837_in3 : std_logic_vector(1 downto 0);
    signal VN837_in4 : std_logic_vector(1 downto 0);
    signal VN837_in5 : std_logic_vector(1 downto 0);
    signal VN838_in0 : std_logic_vector(1 downto 0);
    signal VN838_in1 : std_logic_vector(1 downto 0);
    signal VN838_in2 : std_logic_vector(1 downto 0);
    signal VN838_in3 : std_logic_vector(1 downto 0);
    signal VN838_in4 : std_logic_vector(1 downto 0);
    signal VN838_in5 : std_logic_vector(1 downto 0);
    signal VN839_in0 : std_logic_vector(1 downto 0);
    signal VN839_in1 : std_logic_vector(1 downto 0);
    signal VN839_in2 : std_logic_vector(1 downto 0);
    signal VN839_in3 : std_logic_vector(1 downto 0);
    signal VN839_in4 : std_logic_vector(1 downto 0);
    signal VN839_in5 : std_logic_vector(1 downto 0);
    signal VN840_in0 : std_logic_vector(1 downto 0);
    signal VN840_in1 : std_logic_vector(1 downto 0);
    signal VN840_in2 : std_logic_vector(1 downto 0);
    signal VN840_in3 : std_logic_vector(1 downto 0);
    signal VN840_in4 : std_logic_vector(1 downto 0);
    signal VN840_in5 : std_logic_vector(1 downto 0);
    signal VN841_in0 : std_logic_vector(1 downto 0);
    signal VN841_in1 : std_logic_vector(1 downto 0);
    signal VN841_in2 : std_logic_vector(1 downto 0);
    signal VN841_in3 : std_logic_vector(1 downto 0);
    signal VN841_in4 : std_logic_vector(1 downto 0);
    signal VN841_in5 : std_logic_vector(1 downto 0);
    signal VN842_in0 : std_logic_vector(1 downto 0);
    signal VN842_in1 : std_logic_vector(1 downto 0);
    signal VN842_in2 : std_logic_vector(1 downto 0);
    signal VN842_in3 : std_logic_vector(1 downto 0);
    signal VN842_in4 : std_logic_vector(1 downto 0);
    signal VN842_in5 : std_logic_vector(1 downto 0);
    signal VN843_in0 : std_logic_vector(1 downto 0);
    signal VN843_in1 : std_logic_vector(1 downto 0);
    signal VN843_in2 : std_logic_vector(1 downto 0);
    signal VN843_in3 : std_logic_vector(1 downto 0);
    signal VN843_in4 : std_logic_vector(1 downto 0);
    signal VN843_in5 : std_logic_vector(1 downto 0);
    signal VN844_in0 : std_logic_vector(1 downto 0);
    signal VN844_in1 : std_logic_vector(1 downto 0);
    signal VN844_in2 : std_logic_vector(1 downto 0);
    signal VN844_in3 : std_logic_vector(1 downto 0);
    signal VN844_in4 : std_logic_vector(1 downto 0);
    signal VN844_in5 : std_logic_vector(1 downto 0);
    signal VN845_in0 : std_logic_vector(1 downto 0);
    signal VN845_in1 : std_logic_vector(1 downto 0);
    signal VN845_in2 : std_logic_vector(1 downto 0);
    signal VN845_in3 : std_logic_vector(1 downto 0);
    signal VN845_in4 : std_logic_vector(1 downto 0);
    signal VN845_in5 : std_logic_vector(1 downto 0);
    signal VN846_in0 : std_logic_vector(1 downto 0);
    signal VN846_in1 : std_logic_vector(1 downto 0);
    signal VN846_in2 : std_logic_vector(1 downto 0);
    signal VN846_in3 : std_logic_vector(1 downto 0);
    signal VN846_in4 : std_logic_vector(1 downto 0);
    signal VN846_in5 : std_logic_vector(1 downto 0);
    signal VN847_in0 : std_logic_vector(1 downto 0);
    signal VN847_in1 : std_logic_vector(1 downto 0);
    signal VN847_in2 : std_logic_vector(1 downto 0);
    signal VN847_in3 : std_logic_vector(1 downto 0);
    signal VN847_in4 : std_logic_vector(1 downto 0);
    signal VN847_in5 : std_logic_vector(1 downto 0);
    signal VN848_in0 : std_logic_vector(1 downto 0);
    signal VN848_in1 : std_logic_vector(1 downto 0);
    signal VN848_in2 : std_logic_vector(1 downto 0);
    signal VN848_in3 : std_logic_vector(1 downto 0);
    signal VN848_in4 : std_logic_vector(1 downto 0);
    signal VN848_in5 : std_logic_vector(1 downto 0);
    signal VN849_in0 : std_logic_vector(1 downto 0);
    signal VN849_in1 : std_logic_vector(1 downto 0);
    signal VN849_in2 : std_logic_vector(1 downto 0);
    signal VN849_in3 : std_logic_vector(1 downto 0);
    signal VN849_in4 : std_logic_vector(1 downto 0);
    signal VN849_in5 : std_logic_vector(1 downto 0);
    signal VN850_in0 : std_logic_vector(1 downto 0);
    signal VN850_in1 : std_logic_vector(1 downto 0);
    signal VN850_in2 : std_logic_vector(1 downto 0);
    signal VN850_in3 : std_logic_vector(1 downto 0);
    signal VN850_in4 : std_logic_vector(1 downto 0);
    signal VN850_in5 : std_logic_vector(1 downto 0);
    signal VN851_in0 : std_logic_vector(1 downto 0);
    signal VN851_in1 : std_logic_vector(1 downto 0);
    signal VN851_in2 : std_logic_vector(1 downto 0);
    signal VN851_in3 : std_logic_vector(1 downto 0);
    signal VN851_in4 : std_logic_vector(1 downto 0);
    signal VN851_in5 : std_logic_vector(1 downto 0);
    signal VN852_in0 : std_logic_vector(1 downto 0);
    signal VN852_in1 : std_logic_vector(1 downto 0);
    signal VN852_in2 : std_logic_vector(1 downto 0);
    signal VN852_in3 : std_logic_vector(1 downto 0);
    signal VN852_in4 : std_logic_vector(1 downto 0);
    signal VN852_in5 : std_logic_vector(1 downto 0);
    signal VN853_in0 : std_logic_vector(1 downto 0);
    signal VN853_in1 : std_logic_vector(1 downto 0);
    signal VN853_in2 : std_logic_vector(1 downto 0);
    signal VN853_in3 : std_logic_vector(1 downto 0);
    signal VN853_in4 : std_logic_vector(1 downto 0);
    signal VN853_in5 : std_logic_vector(1 downto 0);
    signal VN854_in0 : std_logic_vector(1 downto 0);
    signal VN854_in1 : std_logic_vector(1 downto 0);
    signal VN854_in2 : std_logic_vector(1 downto 0);
    signal VN854_in3 : std_logic_vector(1 downto 0);
    signal VN854_in4 : std_logic_vector(1 downto 0);
    signal VN854_in5 : std_logic_vector(1 downto 0);
    signal VN855_in0 : std_logic_vector(1 downto 0);
    signal VN855_in1 : std_logic_vector(1 downto 0);
    signal VN855_in2 : std_logic_vector(1 downto 0);
    signal VN855_in3 : std_logic_vector(1 downto 0);
    signal VN855_in4 : std_logic_vector(1 downto 0);
    signal VN855_in5 : std_logic_vector(1 downto 0);
    signal VN856_in0 : std_logic_vector(1 downto 0);
    signal VN856_in1 : std_logic_vector(1 downto 0);
    signal VN856_in2 : std_logic_vector(1 downto 0);
    signal VN856_in3 : std_logic_vector(1 downto 0);
    signal VN856_in4 : std_logic_vector(1 downto 0);
    signal VN856_in5 : std_logic_vector(1 downto 0);
    signal VN857_in0 : std_logic_vector(1 downto 0);
    signal VN857_in1 : std_logic_vector(1 downto 0);
    signal VN857_in2 : std_logic_vector(1 downto 0);
    signal VN857_in3 : std_logic_vector(1 downto 0);
    signal VN857_in4 : std_logic_vector(1 downto 0);
    signal VN857_in5 : std_logic_vector(1 downto 0);
    signal VN858_in0 : std_logic_vector(1 downto 0);
    signal VN858_in1 : std_logic_vector(1 downto 0);
    signal VN858_in2 : std_logic_vector(1 downto 0);
    signal VN858_in3 : std_logic_vector(1 downto 0);
    signal VN858_in4 : std_logic_vector(1 downto 0);
    signal VN858_in5 : std_logic_vector(1 downto 0);
    signal VN859_in0 : std_logic_vector(1 downto 0);
    signal VN859_in1 : std_logic_vector(1 downto 0);
    signal VN859_in2 : std_logic_vector(1 downto 0);
    signal VN859_in3 : std_logic_vector(1 downto 0);
    signal VN859_in4 : std_logic_vector(1 downto 0);
    signal VN859_in5 : std_logic_vector(1 downto 0);
    signal VN860_in0 : std_logic_vector(1 downto 0);
    signal VN860_in1 : std_logic_vector(1 downto 0);
    signal VN860_in2 : std_logic_vector(1 downto 0);
    signal VN860_in3 : std_logic_vector(1 downto 0);
    signal VN860_in4 : std_logic_vector(1 downto 0);
    signal VN860_in5 : std_logic_vector(1 downto 0);
    signal VN861_in0 : std_logic_vector(1 downto 0);
    signal VN861_in1 : std_logic_vector(1 downto 0);
    signal VN861_in2 : std_logic_vector(1 downto 0);
    signal VN861_in3 : std_logic_vector(1 downto 0);
    signal VN861_in4 : std_logic_vector(1 downto 0);
    signal VN861_in5 : std_logic_vector(1 downto 0);
    signal VN862_in0 : std_logic_vector(1 downto 0);
    signal VN862_in1 : std_logic_vector(1 downto 0);
    signal VN862_in2 : std_logic_vector(1 downto 0);
    signal VN862_in3 : std_logic_vector(1 downto 0);
    signal VN862_in4 : std_logic_vector(1 downto 0);
    signal VN862_in5 : std_logic_vector(1 downto 0);
    signal VN863_in0 : std_logic_vector(1 downto 0);
    signal VN863_in1 : std_logic_vector(1 downto 0);
    signal VN863_in2 : std_logic_vector(1 downto 0);
    signal VN863_in3 : std_logic_vector(1 downto 0);
    signal VN863_in4 : std_logic_vector(1 downto 0);
    signal VN863_in5 : std_logic_vector(1 downto 0);
    signal VN864_in0 : std_logic_vector(1 downto 0);
    signal VN864_in1 : std_logic_vector(1 downto 0);
    signal VN864_in2 : std_logic_vector(1 downto 0);
    signal VN864_in3 : std_logic_vector(1 downto 0);
    signal VN864_in4 : std_logic_vector(1 downto 0);
    signal VN864_in5 : std_logic_vector(1 downto 0);
    signal VN865_in0 : std_logic_vector(1 downto 0);
    signal VN865_in1 : std_logic_vector(1 downto 0);
    signal VN865_in2 : std_logic_vector(1 downto 0);
    signal VN865_in3 : std_logic_vector(1 downto 0);
    signal VN865_in4 : std_logic_vector(1 downto 0);
    signal VN865_in5 : std_logic_vector(1 downto 0);
    signal VN866_in0 : std_logic_vector(1 downto 0);
    signal VN866_in1 : std_logic_vector(1 downto 0);
    signal VN866_in2 : std_logic_vector(1 downto 0);
    signal VN866_in3 : std_logic_vector(1 downto 0);
    signal VN866_in4 : std_logic_vector(1 downto 0);
    signal VN866_in5 : std_logic_vector(1 downto 0);
    signal VN867_in0 : std_logic_vector(1 downto 0);
    signal VN867_in1 : std_logic_vector(1 downto 0);
    signal VN867_in2 : std_logic_vector(1 downto 0);
    signal VN867_in3 : std_logic_vector(1 downto 0);
    signal VN867_in4 : std_logic_vector(1 downto 0);
    signal VN867_in5 : std_logic_vector(1 downto 0);
    signal VN868_in0 : std_logic_vector(1 downto 0);
    signal VN868_in1 : std_logic_vector(1 downto 0);
    signal VN868_in2 : std_logic_vector(1 downto 0);
    signal VN868_in3 : std_logic_vector(1 downto 0);
    signal VN868_in4 : std_logic_vector(1 downto 0);
    signal VN868_in5 : std_logic_vector(1 downto 0);
    signal VN869_in0 : std_logic_vector(1 downto 0);
    signal VN869_in1 : std_logic_vector(1 downto 0);
    signal VN869_in2 : std_logic_vector(1 downto 0);
    signal VN869_in3 : std_logic_vector(1 downto 0);
    signal VN869_in4 : std_logic_vector(1 downto 0);
    signal VN869_in5 : std_logic_vector(1 downto 0);
    signal VN870_in0 : std_logic_vector(1 downto 0);
    signal VN870_in1 : std_logic_vector(1 downto 0);
    signal VN870_in2 : std_logic_vector(1 downto 0);
    signal VN870_in3 : std_logic_vector(1 downto 0);
    signal VN870_in4 : std_logic_vector(1 downto 0);
    signal VN870_in5 : std_logic_vector(1 downto 0);
    signal VN871_in0 : std_logic_vector(1 downto 0);
    signal VN871_in1 : std_logic_vector(1 downto 0);
    signal VN871_in2 : std_logic_vector(1 downto 0);
    signal VN871_in3 : std_logic_vector(1 downto 0);
    signal VN871_in4 : std_logic_vector(1 downto 0);
    signal VN871_in5 : std_logic_vector(1 downto 0);
    signal VN872_in0 : std_logic_vector(1 downto 0);
    signal VN872_in1 : std_logic_vector(1 downto 0);
    signal VN872_in2 : std_logic_vector(1 downto 0);
    signal VN872_in3 : std_logic_vector(1 downto 0);
    signal VN872_in4 : std_logic_vector(1 downto 0);
    signal VN872_in5 : std_logic_vector(1 downto 0);
    signal VN873_in0 : std_logic_vector(1 downto 0);
    signal VN873_in1 : std_logic_vector(1 downto 0);
    signal VN873_in2 : std_logic_vector(1 downto 0);
    signal VN873_in3 : std_logic_vector(1 downto 0);
    signal VN873_in4 : std_logic_vector(1 downto 0);
    signal VN873_in5 : std_logic_vector(1 downto 0);
    signal VN874_in0 : std_logic_vector(1 downto 0);
    signal VN874_in1 : std_logic_vector(1 downto 0);
    signal VN874_in2 : std_logic_vector(1 downto 0);
    signal VN874_in3 : std_logic_vector(1 downto 0);
    signal VN874_in4 : std_logic_vector(1 downto 0);
    signal VN874_in5 : std_logic_vector(1 downto 0);
    signal VN875_in0 : std_logic_vector(1 downto 0);
    signal VN875_in1 : std_logic_vector(1 downto 0);
    signal VN875_in2 : std_logic_vector(1 downto 0);
    signal VN875_in3 : std_logic_vector(1 downto 0);
    signal VN875_in4 : std_logic_vector(1 downto 0);
    signal VN875_in5 : std_logic_vector(1 downto 0);
    signal VN876_in0 : std_logic_vector(1 downto 0);
    signal VN876_in1 : std_logic_vector(1 downto 0);
    signal VN876_in2 : std_logic_vector(1 downto 0);
    signal VN876_in3 : std_logic_vector(1 downto 0);
    signal VN876_in4 : std_logic_vector(1 downto 0);
    signal VN876_in5 : std_logic_vector(1 downto 0);
    signal VN877_in0 : std_logic_vector(1 downto 0);
    signal VN877_in1 : std_logic_vector(1 downto 0);
    signal VN877_in2 : std_logic_vector(1 downto 0);
    signal VN877_in3 : std_logic_vector(1 downto 0);
    signal VN877_in4 : std_logic_vector(1 downto 0);
    signal VN877_in5 : std_logic_vector(1 downto 0);
    signal VN878_in0 : std_logic_vector(1 downto 0);
    signal VN878_in1 : std_logic_vector(1 downto 0);
    signal VN878_in2 : std_logic_vector(1 downto 0);
    signal VN878_in3 : std_logic_vector(1 downto 0);
    signal VN878_in4 : std_logic_vector(1 downto 0);
    signal VN878_in5 : std_logic_vector(1 downto 0);
    signal VN879_in0 : std_logic_vector(1 downto 0);
    signal VN879_in1 : std_logic_vector(1 downto 0);
    signal VN879_in2 : std_logic_vector(1 downto 0);
    signal VN879_in3 : std_logic_vector(1 downto 0);
    signal VN879_in4 : std_logic_vector(1 downto 0);
    signal VN879_in5 : std_logic_vector(1 downto 0);
    signal VN880_in0 : std_logic_vector(1 downto 0);
    signal VN880_in1 : std_logic_vector(1 downto 0);
    signal VN880_in2 : std_logic_vector(1 downto 0);
    signal VN880_in3 : std_logic_vector(1 downto 0);
    signal VN880_in4 : std_logic_vector(1 downto 0);
    signal VN880_in5 : std_logic_vector(1 downto 0);
    signal VN881_in0 : std_logic_vector(1 downto 0);
    signal VN881_in1 : std_logic_vector(1 downto 0);
    signal VN881_in2 : std_logic_vector(1 downto 0);
    signal VN881_in3 : std_logic_vector(1 downto 0);
    signal VN881_in4 : std_logic_vector(1 downto 0);
    signal VN881_in5 : std_logic_vector(1 downto 0);
    signal VN882_in0 : std_logic_vector(1 downto 0);
    signal VN882_in1 : std_logic_vector(1 downto 0);
    signal VN882_in2 : std_logic_vector(1 downto 0);
    signal VN882_in3 : std_logic_vector(1 downto 0);
    signal VN882_in4 : std_logic_vector(1 downto 0);
    signal VN882_in5 : std_logic_vector(1 downto 0);
    signal VN883_in0 : std_logic_vector(1 downto 0);
    signal VN883_in1 : std_logic_vector(1 downto 0);
    signal VN883_in2 : std_logic_vector(1 downto 0);
    signal VN883_in3 : std_logic_vector(1 downto 0);
    signal VN883_in4 : std_logic_vector(1 downto 0);
    signal VN883_in5 : std_logic_vector(1 downto 0);
    signal VN884_in0 : std_logic_vector(1 downto 0);
    signal VN884_in1 : std_logic_vector(1 downto 0);
    signal VN884_in2 : std_logic_vector(1 downto 0);
    signal VN884_in3 : std_logic_vector(1 downto 0);
    signal VN884_in4 : std_logic_vector(1 downto 0);
    signal VN884_in5 : std_logic_vector(1 downto 0);
    signal VN885_in0 : std_logic_vector(1 downto 0);
    signal VN885_in1 : std_logic_vector(1 downto 0);
    signal VN885_in2 : std_logic_vector(1 downto 0);
    signal VN885_in3 : std_logic_vector(1 downto 0);
    signal VN885_in4 : std_logic_vector(1 downto 0);
    signal VN885_in5 : std_logic_vector(1 downto 0);
    signal VN886_in0 : std_logic_vector(1 downto 0);
    signal VN886_in1 : std_logic_vector(1 downto 0);
    signal VN886_in2 : std_logic_vector(1 downto 0);
    signal VN886_in3 : std_logic_vector(1 downto 0);
    signal VN886_in4 : std_logic_vector(1 downto 0);
    signal VN886_in5 : std_logic_vector(1 downto 0);
    signal VN887_in0 : std_logic_vector(1 downto 0);
    signal VN887_in1 : std_logic_vector(1 downto 0);
    signal VN887_in2 : std_logic_vector(1 downto 0);
    signal VN887_in3 : std_logic_vector(1 downto 0);
    signal VN887_in4 : std_logic_vector(1 downto 0);
    signal VN887_in5 : std_logic_vector(1 downto 0);
    signal VN888_in0 : std_logic_vector(1 downto 0);
    signal VN888_in1 : std_logic_vector(1 downto 0);
    signal VN888_in2 : std_logic_vector(1 downto 0);
    signal VN888_in3 : std_logic_vector(1 downto 0);
    signal VN888_in4 : std_logic_vector(1 downto 0);
    signal VN888_in5 : std_logic_vector(1 downto 0);
    signal VN889_in0 : std_logic_vector(1 downto 0);
    signal VN889_in1 : std_logic_vector(1 downto 0);
    signal VN889_in2 : std_logic_vector(1 downto 0);
    signal VN889_in3 : std_logic_vector(1 downto 0);
    signal VN889_in4 : std_logic_vector(1 downto 0);
    signal VN889_in5 : std_logic_vector(1 downto 0);
    signal VN890_in0 : std_logic_vector(1 downto 0);
    signal VN890_in1 : std_logic_vector(1 downto 0);
    signal VN890_in2 : std_logic_vector(1 downto 0);
    signal VN890_in3 : std_logic_vector(1 downto 0);
    signal VN890_in4 : std_logic_vector(1 downto 0);
    signal VN890_in5 : std_logic_vector(1 downto 0);
    signal VN891_in0 : std_logic_vector(1 downto 0);
    signal VN891_in1 : std_logic_vector(1 downto 0);
    signal VN891_in2 : std_logic_vector(1 downto 0);
    signal VN891_in3 : std_logic_vector(1 downto 0);
    signal VN891_in4 : std_logic_vector(1 downto 0);
    signal VN891_in5 : std_logic_vector(1 downto 0);
    signal VN892_in0 : std_logic_vector(1 downto 0);
    signal VN892_in1 : std_logic_vector(1 downto 0);
    signal VN892_in2 : std_logic_vector(1 downto 0);
    signal VN892_in3 : std_logic_vector(1 downto 0);
    signal VN892_in4 : std_logic_vector(1 downto 0);
    signal VN892_in5 : std_logic_vector(1 downto 0);
    signal VN893_in0 : std_logic_vector(1 downto 0);
    signal VN893_in1 : std_logic_vector(1 downto 0);
    signal VN893_in2 : std_logic_vector(1 downto 0);
    signal VN893_in3 : std_logic_vector(1 downto 0);
    signal VN893_in4 : std_logic_vector(1 downto 0);
    signal VN893_in5 : std_logic_vector(1 downto 0);
    signal VN894_in0 : std_logic_vector(1 downto 0);
    signal VN894_in1 : std_logic_vector(1 downto 0);
    signal VN894_in2 : std_logic_vector(1 downto 0);
    signal VN894_in3 : std_logic_vector(1 downto 0);
    signal VN894_in4 : std_logic_vector(1 downto 0);
    signal VN894_in5 : std_logic_vector(1 downto 0);
    signal VN895_in0 : std_logic_vector(1 downto 0);
    signal VN895_in1 : std_logic_vector(1 downto 0);
    signal VN895_in2 : std_logic_vector(1 downto 0);
    signal VN895_in3 : std_logic_vector(1 downto 0);
    signal VN895_in4 : std_logic_vector(1 downto 0);
    signal VN895_in5 : std_logic_vector(1 downto 0);
    signal VN896_in0 : std_logic_vector(1 downto 0);
    signal VN896_in1 : std_logic_vector(1 downto 0);
    signal VN896_in2 : std_logic_vector(1 downto 0);
    signal VN896_in3 : std_logic_vector(1 downto 0);
    signal VN896_in4 : std_logic_vector(1 downto 0);
    signal VN896_in5 : std_logic_vector(1 downto 0);
    signal VN897_in0 : std_logic_vector(1 downto 0);
    signal VN897_in1 : std_logic_vector(1 downto 0);
    signal VN897_in2 : std_logic_vector(1 downto 0);
    signal VN897_in3 : std_logic_vector(1 downto 0);
    signal VN897_in4 : std_logic_vector(1 downto 0);
    signal VN897_in5 : std_logic_vector(1 downto 0);
    signal VN898_in0 : std_logic_vector(1 downto 0);
    signal VN898_in1 : std_logic_vector(1 downto 0);
    signal VN898_in2 : std_logic_vector(1 downto 0);
    signal VN898_in3 : std_logic_vector(1 downto 0);
    signal VN898_in4 : std_logic_vector(1 downto 0);
    signal VN898_in5 : std_logic_vector(1 downto 0);
    signal VN899_in0 : std_logic_vector(1 downto 0);
    signal VN899_in1 : std_logic_vector(1 downto 0);
    signal VN899_in2 : std_logic_vector(1 downto 0);
    signal VN899_in3 : std_logic_vector(1 downto 0);
    signal VN899_in4 : std_logic_vector(1 downto 0);
    signal VN899_in5 : std_logic_vector(1 downto 0);
    signal VN900_in0 : std_logic_vector(1 downto 0);
    signal VN900_in1 : std_logic_vector(1 downto 0);
    signal VN900_in2 : std_logic_vector(1 downto 0);
    signal VN900_in3 : std_logic_vector(1 downto 0);
    signal VN900_in4 : std_logic_vector(1 downto 0);
    signal VN900_in5 : std_logic_vector(1 downto 0);
    signal VN901_in0 : std_logic_vector(1 downto 0);
    signal VN901_in1 : std_logic_vector(1 downto 0);
    signal VN901_in2 : std_logic_vector(1 downto 0);
    signal VN901_in3 : std_logic_vector(1 downto 0);
    signal VN901_in4 : std_logic_vector(1 downto 0);
    signal VN901_in5 : std_logic_vector(1 downto 0);
    signal VN902_in0 : std_logic_vector(1 downto 0);
    signal VN902_in1 : std_logic_vector(1 downto 0);
    signal VN902_in2 : std_logic_vector(1 downto 0);
    signal VN902_in3 : std_logic_vector(1 downto 0);
    signal VN902_in4 : std_logic_vector(1 downto 0);
    signal VN902_in5 : std_logic_vector(1 downto 0);
    signal VN903_in0 : std_logic_vector(1 downto 0);
    signal VN903_in1 : std_logic_vector(1 downto 0);
    signal VN903_in2 : std_logic_vector(1 downto 0);
    signal VN903_in3 : std_logic_vector(1 downto 0);
    signal VN903_in4 : std_logic_vector(1 downto 0);
    signal VN903_in5 : std_logic_vector(1 downto 0);
    signal VN904_in0 : std_logic_vector(1 downto 0);
    signal VN904_in1 : std_logic_vector(1 downto 0);
    signal VN904_in2 : std_logic_vector(1 downto 0);
    signal VN904_in3 : std_logic_vector(1 downto 0);
    signal VN904_in4 : std_logic_vector(1 downto 0);
    signal VN904_in5 : std_logic_vector(1 downto 0);
    signal VN905_in0 : std_logic_vector(1 downto 0);
    signal VN905_in1 : std_logic_vector(1 downto 0);
    signal VN905_in2 : std_logic_vector(1 downto 0);
    signal VN905_in3 : std_logic_vector(1 downto 0);
    signal VN905_in4 : std_logic_vector(1 downto 0);
    signal VN905_in5 : std_logic_vector(1 downto 0);
    signal VN906_in0 : std_logic_vector(1 downto 0);
    signal VN906_in1 : std_logic_vector(1 downto 0);
    signal VN906_in2 : std_logic_vector(1 downto 0);
    signal VN906_in3 : std_logic_vector(1 downto 0);
    signal VN906_in4 : std_logic_vector(1 downto 0);
    signal VN906_in5 : std_logic_vector(1 downto 0);
    signal VN907_in0 : std_logic_vector(1 downto 0);
    signal VN907_in1 : std_logic_vector(1 downto 0);
    signal VN907_in2 : std_logic_vector(1 downto 0);
    signal VN907_in3 : std_logic_vector(1 downto 0);
    signal VN907_in4 : std_logic_vector(1 downto 0);
    signal VN907_in5 : std_logic_vector(1 downto 0);
    signal VN908_in0 : std_logic_vector(1 downto 0);
    signal VN908_in1 : std_logic_vector(1 downto 0);
    signal VN908_in2 : std_logic_vector(1 downto 0);
    signal VN908_in3 : std_logic_vector(1 downto 0);
    signal VN908_in4 : std_logic_vector(1 downto 0);
    signal VN908_in5 : std_logic_vector(1 downto 0);
    signal VN909_in0 : std_logic_vector(1 downto 0);
    signal VN909_in1 : std_logic_vector(1 downto 0);
    signal VN909_in2 : std_logic_vector(1 downto 0);
    signal VN909_in3 : std_logic_vector(1 downto 0);
    signal VN909_in4 : std_logic_vector(1 downto 0);
    signal VN909_in5 : std_logic_vector(1 downto 0);
    signal VN910_in0 : std_logic_vector(1 downto 0);
    signal VN910_in1 : std_logic_vector(1 downto 0);
    signal VN910_in2 : std_logic_vector(1 downto 0);
    signal VN910_in3 : std_logic_vector(1 downto 0);
    signal VN910_in4 : std_logic_vector(1 downto 0);
    signal VN910_in5 : std_logic_vector(1 downto 0);
    signal VN911_in0 : std_logic_vector(1 downto 0);
    signal VN911_in1 : std_logic_vector(1 downto 0);
    signal VN911_in2 : std_logic_vector(1 downto 0);
    signal VN911_in3 : std_logic_vector(1 downto 0);
    signal VN911_in4 : std_logic_vector(1 downto 0);
    signal VN911_in5 : std_logic_vector(1 downto 0);
    signal VN912_in0 : std_logic_vector(1 downto 0);
    signal VN912_in1 : std_logic_vector(1 downto 0);
    signal VN912_in2 : std_logic_vector(1 downto 0);
    signal VN912_in3 : std_logic_vector(1 downto 0);
    signal VN912_in4 : std_logic_vector(1 downto 0);
    signal VN912_in5 : std_logic_vector(1 downto 0);
    signal VN913_in0 : std_logic_vector(1 downto 0);
    signal VN913_in1 : std_logic_vector(1 downto 0);
    signal VN913_in2 : std_logic_vector(1 downto 0);
    signal VN913_in3 : std_logic_vector(1 downto 0);
    signal VN913_in4 : std_logic_vector(1 downto 0);
    signal VN913_in5 : std_logic_vector(1 downto 0);
    signal VN914_in0 : std_logic_vector(1 downto 0);
    signal VN914_in1 : std_logic_vector(1 downto 0);
    signal VN914_in2 : std_logic_vector(1 downto 0);
    signal VN914_in3 : std_logic_vector(1 downto 0);
    signal VN914_in4 : std_logic_vector(1 downto 0);
    signal VN914_in5 : std_logic_vector(1 downto 0);
    signal VN915_in0 : std_logic_vector(1 downto 0);
    signal VN915_in1 : std_logic_vector(1 downto 0);
    signal VN915_in2 : std_logic_vector(1 downto 0);
    signal VN915_in3 : std_logic_vector(1 downto 0);
    signal VN915_in4 : std_logic_vector(1 downto 0);
    signal VN915_in5 : std_logic_vector(1 downto 0);
    signal VN916_in0 : std_logic_vector(1 downto 0);
    signal VN916_in1 : std_logic_vector(1 downto 0);
    signal VN916_in2 : std_logic_vector(1 downto 0);
    signal VN916_in3 : std_logic_vector(1 downto 0);
    signal VN916_in4 : std_logic_vector(1 downto 0);
    signal VN916_in5 : std_logic_vector(1 downto 0);
    signal VN917_in0 : std_logic_vector(1 downto 0);
    signal VN917_in1 : std_logic_vector(1 downto 0);
    signal VN917_in2 : std_logic_vector(1 downto 0);
    signal VN917_in3 : std_logic_vector(1 downto 0);
    signal VN917_in4 : std_logic_vector(1 downto 0);
    signal VN917_in5 : std_logic_vector(1 downto 0);
    signal VN918_in0 : std_logic_vector(1 downto 0);
    signal VN918_in1 : std_logic_vector(1 downto 0);
    signal VN918_in2 : std_logic_vector(1 downto 0);
    signal VN918_in3 : std_logic_vector(1 downto 0);
    signal VN918_in4 : std_logic_vector(1 downto 0);
    signal VN918_in5 : std_logic_vector(1 downto 0);
    signal VN919_in0 : std_logic_vector(1 downto 0);
    signal VN919_in1 : std_logic_vector(1 downto 0);
    signal VN919_in2 : std_logic_vector(1 downto 0);
    signal VN919_in3 : std_logic_vector(1 downto 0);
    signal VN919_in4 : std_logic_vector(1 downto 0);
    signal VN919_in5 : std_logic_vector(1 downto 0);
    signal VN920_in0 : std_logic_vector(1 downto 0);
    signal VN920_in1 : std_logic_vector(1 downto 0);
    signal VN920_in2 : std_logic_vector(1 downto 0);
    signal VN920_in3 : std_logic_vector(1 downto 0);
    signal VN920_in4 : std_logic_vector(1 downto 0);
    signal VN920_in5 : std_logic_vector(1 downto 0);
    signal VN921_in0 : std_logic_vector(1 downto 0);
    signal VN921_in1 : std_logic_vector(1 downto 0);
    signal VN921_in2 : std_logic_vector(1 downto 0);
    signal VN921_in3 : std_logic_vector(1 downto 0);
    signal VN921_in4 : std_logic_vector(1 downto 0);
    signal VN921_in5 : std_logic_vector(1 downto 0);
    signal VN922_in0 : std_logic_vector(1 downto 0);
    signal VN922_in1 : std_logic_vector(1 downto 0);
    signal VN922_in2 : std_logic_vector(1 downto 0);
    signal VN922_in3 : std_logic_vector(1 downto 0);
    signal VN922_in4 : std_logic_vector(1 downto 0);
    signal VN922_in5 : std_logic_vector(1 downto 0);
    signal VN923_in0 : std_logic_vector(1 downto 0);
    signal VN923_in1 : std_logic_vector(1 downto 0);
    signal VN923_in2 : std_logic_vector(1 downto 0);
    signal VN923_in3 : std_logic_vector(1 downto 0);
    signal VN923_in4 : std_logic_vector(1 downto 0);
    signal VN923_in5 : std_logic_vector(1 downto 0);
    signal VN924_in0 : std_logic_vector(1 downto 0);
    signal VN924_in1 : std_logic_vector(1 downto 0);
    signal VN924_in2 : std_logic_vector(1 downto 0);
    signal VN924_in3 : std_logic_vector(1 downto 0);
    signal VN924_in4 : std_logic_vector(1 downto 0);
    signal VN924_in5 : std_logic_vector(1 downto 0);
    signal VN925_in0 : std_logic_vector(1 downto 0);
    signal VN925_in1 : std_logic_vector(1 downto 0);
    signal VN925_in2 : std_logic_vector(1 downto 0);
    signal VN925_in3 : std_logic_vector(1 downto 0);
    signal VN925_in4 : std_logic_vector(1 downto 0);
    signal VN925_in5 : std_logic_vector(1 downto 0);
    signal VN926_in0 : std_logic_vector(1 downto 0);
    signal VN926_in1 : std_logic_vector(1 downto 0);
    signal VN926_in2 : std_logic_vector(1 downto 0);
    signal VN926_in3 : std_logic_vector(1 downto 0);
    signal VN926_in4 : std_logic_vector(1 downto 0);
    signal VN926_in5 : std_logic_vector(1 downto 0);
    signal VN927_in0 : std_logic_vector(1 downto 0);
    signal VN927_in1 : std_logic_vector(1 downto 0);
    signal VN927_in2 : std_logic_vector(1 downto 0);
    signal VN927_in3 : std_logic_vector(1 downto 0);
    signal VN927_in4 : std_logic_vector(1 downto 0);
    signal VN927_in5 : std_logic_vector(1 downto 0);
    signal VN928_in0 : std_logic_vector(1 downto 0);
    signal VN928_in1 : std_logic_vector(1 downto 0);
    signal VN928_in2 : std_logic_vector(1 downto 0);
    signal VN928_in3 : std_logic_vector(1 downto 0);
    signal VN928_in4 : std_logic_vector(1 downto 0);
    signal VN928_in5 : std_logic_vector(1 downto 0);
    signal VN929_in0 : std_logic_vector(1 downto 0);
    signal VN929_in1 : std_logic_vector(1 downto 0);
    signal VN929_in2 : std_logic_vector(1 downto 0);
    signal VN929_in3 : std_logic_vector(1 downto 0);
    signal VN929_in4 : std_logic_vector(1 downto 0);
    signal VN929_in5 : std_logic_vector(1 downto 0);
    signal VN930_in0 : std_logic_vector(1 downto 0);
    signal VN930_in1 : std_logic_vector(1 downto 0);
    signal VN930_in2 : std_logic_vector(1 downto 0);
    signal VN930_in3 : std_logic_vector(1 downto 0);
    signal VN930_in4 : std_logic_vector(1 downto 0);
    signal VN930_in5 : std_logic_vector(1 downto 0);
    signal VN931_in0 : std_logic_vector(1 downto 0);
    signal VN931_in1 : std_logic_vector(1 downto 0);
    signal VN931_in2 : std_logic_vector(1 downto 0);
    signal VN931_in3 : std_logic_vector(1 downto 0);
    signal VN931_in4 : std_logic_vector(1 downto 0);
    signal VN931_in5 : std_logic_vector(1 downto 0);
    signal VN932_in0 : std_logic_vector(1 downto 0);
    signal VN932_in1 : std_logic_vector(1 downto 0);
    signal VN932_in2 : std_logic_vector(1 downto 0);
    signal VN932_in3 : std_logic_vector(1 downto 0);
    signal VN932_in4 : std_logic_vector(1 downto 0);
    signal VN932_in5 : std_logic_vector(1 downto 0);
    signal VN933_in0 : std_logic_vector(1 downto 0);
    signal VN933_in1 : std_logic_vector(1 downto 0);
    signal VN933_in2 : std_logic_vector(1 downto 0);
    signal VN933_in3 : std_logic_vector(1 downto 0);
    signal VN933_in4 : std_logic_vector(1 downto 0);
    signal VN933_in5 : std_logic_vector(1 downto 0);
    signal VN934_in0 : std_logic_vector(1 downto 0);
    signal VN934_in1 : std_logic_vector(1 downto 0);
    signal VN934_in2 : std_logic_vector(1 downto 0);
    signal VN934_in3 : std_logic_vector(1 downto 0);
    signal VN934_in4 : std_logic_vector(1 downto 0);
    signal VN934_in5 : std_logic_vector(1 downto 0);
    signal VN935_in0 : std_logic_vector(1 downto 0);
    signal VN935_in1 : std_logic_vector(1 downto 0);
    signal VN935_in2 : std_logic_vector(1 downto 0);
    signal VN935_in3 : std_logic_vector(1 downto 0);
    signal VN935_in4 : std_logic_vector(1 downto 0);
    signal VN935_in5 : std_logic_vector(1 downto 0);
    signal VN936_in0 : std_logic_vector(1 downto 0);
    signal VN936_in1 : std_logic_vector(1 downto 0);
    signal VN936_in2 : std_logic_vector(1 downto 0);
    signal VN936_in3 : std_logic_vector(1 downto 0);
    signal VN936_in4 : std_logic_vector(1 downto 0);
    signal VN936_in5 : std_logic_vector(1 downto 0);
    signal VN937_in0 : std_logic_vector(1 downto 0);
    signal VN937_in1 : std_logic_vector(1 downto 0);
    signal VN937_in2 : std_logic_vector(1 downto 0);
    signal VN937_in3 : std_logic_vector(1 downto 0);
    signal VN937_in4 : std_logic_vector(1 downto 0);
    signal VN937_in5 : std_logic_vector(1 downto 0);
    signal VN938_in0 : std_logic_vector(1 downto 0);
    signal VN938_in1 : std_logic_vector(1 downto 0);
    signal VN938_in2 : std_logic_vector(1 downto 0);
    signal VN938_in3 : std_logic_vector(1 downto 0);
    signal VN938_in4 : std_logic_vector(1 downto 0);
    signal VN938_in5 : std_logic_vector(1 downto 0);
    signal VN939_in0 : std_logic_vector(1 downto 0);
    signal VN939_in1 : std_logic_vector(1 downto 0);
    signal VN939_in2 : std_logic_vector(1 downto 0);
    signal VN939_in3 : std_logic_vector(1 downto 0);
    signal VN939_in4 : std_logic_vector(1 downto 0);
    signal VN939_in5 : std_logic_vector(1 downto 0);
    signal VN940_in0 : std_logic_vector(1 downto 0);
    signal VN940_in1 : std_logic_vector(1 downto 0);
    signal VN940_in2 : std_logic_vector(1 downto 0);
    signal VN940_in3 : std_logic_vector(1 downto 0);
    signal VN940_in4 : std_logic_vector(1 downto 0);
    signal VN940_in5 : std_logic_vector(1 downto 0);
    signal VN941_in0 : std_logic_vector(1 downto 0);
    signal VN941_in1 : std_logic_vector(1 downto 0);
    signal VN941_in2 : std_logic_vector(1 downto 0);
    signal VN941_in3 : std_logic_vector(1 downto 0);
    signal VN941_in4 : std_logic_vector(1 downto 0);
    signal VN941_in5 : std_logic_vector(1 downto 0);
    signal VN942_in0 : std_logic_vector(1 downto 0);
    signal VN942_in1 : std_logic_vector(1 downto 0);
    signal VN942_in2 : std_logic_vector(1 downto 0);
    signal VN942_in3 : std_logic_vector(1 downto 0);
    signal VN942_in4 : std_logic_vector(1 downto 0);
    signal VN942_in5 : std_logic_vector(1 downto 0);
    signal VN943_in0 : std_logic_vector(1 downto 0);
    signal VN943_in1 : std_logic_vector(1 downto 0);
    signal VN943_in2 : std_logic_vector(1 downto 0);
    signal VN943_in3 : std_logic_vector(1 downto 0);
    signal VN943_in4 : std_logic_vector(1 downto 0);
    signal VN943_in5 : std_logic_vector(1 downto 0);
    signal VN944_in0 : std_logic_vector(1 downto 0);
    signal VN944_in1 : std_logic_vector(1 downto 0);
    signal VN944_in2 : std_logic_vector(1 downto 0);
    signal VN944_in3 : std_logic_vector(1 downto 0);
    signal VN944_in4 : std_logic_vector(1 downto 0);
    signal VN944_in5 : std_logic_vector(1 downto 0);
    signal VN945_in0 : std_logic_vector(1 downto 0);
    signal VN945_in1 : std_logic_vector(1 downto 0);
    signal VN945_in2 : std_logic_vector(1 downto 0);
    signal VN945_in3 : std_logic_vector(1 downto 0);
    signal VN945_in4 : std_logic_vector(1 downto 0);
    signal VN945_in5 : std_logic_vector(1 downto 0);
    signal VN946_in0 : std_logic_vector(1 downto 0);
    signal VN946_in1 : std_logic_vector(1 downto 0);
    signal VN946_in2 : std_logic_vector(1 downto 0);
    signal VN946_in3 : std_logic_vector(1 downto 0);
    signal VN946_in4 : std_logic_vector(1 downto 0);
    signal VN946_in5 : std_logic_vector(1 downto 0);
    signal VN947_in0 : std_logic_vector(1 downto 0);
    signal VN947_in1 : std_logic_vector(1 downto 0);
    signal VN947_in2 : std_logic_vector(1 downto 0);
    signal VN947_in3 : std_logic_vector(1 downto 0);
    signal VN947_in4 : std_logic_vector(1 downto 0);
    signal VN947_in5 : std_logic_vector(1 downto 0);
    signal VN948_in0 : std_logic_vector(1 downto 0);
    signal VN948_in1 : std_logic_vector(1 downto 0);
    signal VN948_in2 : std_logic_vector(1 downto 0);
    signal VN948_in3 : std_logic_vector(1 downto 0);
    signal VN948_in4 : std_logic_vector(1 downto 0);
    signal VN948_in5 : std_logic_vector(1 downto 0);
    signal VN949_in0 : std_logic_vector(1 downto 0);
    signal VN949_in1 : std_logic_vector(1 downto 0);
    signal VN949_in2 : std_logic_vector(1 downto 0);
    signal VN949_in3 : std_logic_vector(1 downto 0);
    signal VN949_in4 : std_logic_vector(1 downto 0);
    signal VN949_in5 : std_logic_vector(1 downto 0);
    signal VN950_in0 : std_logic_vector(1 downto 0);
    signal VN950_in1 : std_logic_vector(1 downto 0);
    signal VN950_in2 : std_logic_vector(1 downto 0);
    signal VN950_in3 : std_logic_vector(1 downto 0);
    signal VN950_in4 : std_logic_vector(1 downto 0);
    signal VN950_in5 : std_logic_vector(1 downto 0);
    signal VN951_in0 : std_logic_vector(1 downto 0);
    signal VN951_in1 : std_logic_vector(1 downto 0);
    signal VN951_in2 : std_logic_vector(1 downto 0);
    signal VN951_in3 : std_logic_vector(1 downto 0);
    signal VN951_in4 : std_logic_vector(1 downto 0);
    signal VN951_in5 : std_logic_vector(1 downto 0);
    signal VN952_in0 : std_logic_vector(1 downto 0);
    signal VN952_in1 : std_logic_vector(1 downto 0);
    signal VN952_in2 : std_logic_vector(1 downto 0);
    signal VN952_in3 : std_logic_vector(1 downto 0);
    signal VN952_in4 : std_logic_vector(1 downto 0);
    signal VN952_in5 : std_logic_vector(1 downto 0);
    signal VN953_in0 : std_logic_vector(1 downto 0);
    signal VN953_in1 : std_logic_vector(1 downto 0);
    signal VN953_in2 : std_logic_vector(1 downto 0);
    signal VN953_in3 : std_logic_vector(1 downto 0);
    signal VN953_in4 : std_logic_vector(1 downto 0);
    signal VN953_in5 : std_logic_vector(1 downto 0);
    signal VN954_in0 : std_logic_vector(1 downto 0);
    signal VN954_in1 : std_logic_vector(1 downto 0);
    signal VN954_in2 : std_logic_vector(1 downto 0);
    signal VN954_in3 : std_logic_vector(1 downto 0);
    signal VN954_in4 : std_logic_vector(1 downto 0);
    signal VN954_in5 : std_logic_vector(1 downto 0);
    signal VN955_in0 : std_logic_vector(1 downto 0);
    signal VN955_in1 : std_logic_vector(1 downto 0);
    signal VN955_in2 : std_logic_vector(1 downto 0);
    signal VN955_in3 : std_logic_vector(1 downto 0);
    signal VN955_in4 : std_logic_vector(1 downto 0);
    signal VN955_in5 : std_logic_vector(1 downto 0);
    signal VN956_in0 : std_logic_vector(1 downto 0);
    signal VN956_in1 : std_logic_vector(1 downto 0);
    signal VN956_in2 : std_logic_vector(1 downto 0);
    signal VN956_in3 : std_logic_vector(1 downto 0);
    signal VN956_in4 : std_logic_vector(1 downto 0);
    signal VN956_in5 : std_logic_vector(1 downto 0);
    signal VN957_in0 : std_logic_vector(1 downto 0);
    signal VN957_in1 : std_logic_vector(1 downto 0);
    signal VN957_in2 : std_logic_vector(1 downto 0);
    signal VN957_in3 : std_logic_vector(1 downto 0);
    signal VN957_in4 : std_logic_vector(1 downto 0);
    signal VN957_in5 : std_logic_vector(1 downto 0);
    signal VN958_in0 : std_logic_vector(1 downto 0);
    signal VN958_in1 : std_logic_vector(1 downto 0);
    signal VN958_in2 : std_logic_vector(1 downto 0);
    signal VN958_in3 : std_logic_vector(1 downto 0);
    signal VN958_in4 : std_logic_vector(1 downto 0);
    signal VN958_in5 : std_logic_vector(1 downto 0);
    signal VN959_in0 : std_logic_vector(1 downto 0);
    signal VN959_in1 : std_logic_vector(1 downto 0);
    signal VN959_in2 : std_logic_vector(1 downto 0);
    signal VN959_in3 : std_logic_vector(1 downto 0);
    signal VN959_in4 : std_logic_vector(1 downto 0);
    signal VN959_in5 : std_logic_vector(1 downto 0);
    signal VN960_in0 : std_logic_vector(1 downto 0);
    signal VN960_in1 : std_logic_vector(1 downto 0);
    signal VN960_in2 : std_logic_vector(1 downto 0);
    signal VN960_in3 : std_logic_vector(1 downto 0);
    signal VN960_in4 : std_logic_vector(1 downto 0);
    signal VN960_in5 : std_logic_vector(1 downto 0);
    signal VN961_in0 : std_logic_vector(1 downto 0);
    signal VN961_in1 : std_logic_vector(1 downto 0);
    signal VN961_in2 : std_logic_vector(1 downto 0);
    signal VN961_in3 : std_logic_vector(1 downto 0);
    signal VN961_in4 : std_logic_vector(1 downto 0);
    signal VN961_in5 : std_logic_vector(1 downto 0);
    signal VN962_in0 : std_logic_vector(1 downto 0);
    signal VN962_in1 : std_logic_vector(1 downto 0);
    signal VN962_in2 : std_logic_vector(1 downto 0);
    signal VN962_in3 : std_logic_vector(1 downto 0);
    signal VN962_in4 : std_logic_vector(1 downto 0);
    signal VN962_in5 : std_logic_vector(1 downto 0);
    signal VN963_in0 : std_logic_vector(1 downto 0);
    signal VN963_in1 : std_logic_vector(1 downto 0);
    signal VN963_in2 : std_logic_vector(1 downto 0);
    signal VN963_in3 : std_logic_vector(1 downto 0);
    signal VN963_in4 : std_logic_vector(1 downto 0);
    signal VN963_in5 : std_logic_vector(1 downto 0);
    signal VN964_in0 : std_logic_vector(1 downto 0);
    signal VN964_in1 : std_logic_vector(1 downto 0);
    signal VN964_in2 : std_logic_vector(1 downto 0);
    signal VN964_in3 : std_logic_vector(1 downto 0);
    signal VN964_in4 : std_logic_vector(1 downto 0);
    signal VN964_in5 : std_logic_vector(1 downto 0);
    signal VN965_in0 : std_logic_vector(1 downto 0);
    signal VN965_in1 : std_logic_vector(1 downto 0);
    signal VN965_in2 : std_logic_vector(1 downto 0);
    signal VN965_in3 : std_logic_vector(1 downto 0);
    signal VN965_in4 : std_logic_vector(1 downto 0);
    signal VN965_in5 : std_logic_vector(1 downto 0);
    signal VN966_in0 : std_logic_vector(1 downto 0);
    signal VN966_in1 : std_logic_vector(1 downto 0);
    signal VN966_in2 : std_logic_vector(1 downto 0);
    signal VN966_in3 : std_logic_vector(1 downto 0);
    signal VN966_in4 : std_logic_vector(1 downto 0);
    signal VN966_in5 : std_logic_vector(1 downto 0);
    signal VN967_in0 : std_logic_vector(1 downto 0);
    signal VN967_in1 : std_logic_vector(1 downto 0);
    signal VN967_in2 : std_logic_vector(1 downto 0);
    signal VN967_in3 : std_logic_vector(1 downto 0);
    signal VN967_in4 : std_logic_vector(1 downto 0);
    signal VN967_in5 : std_logic_vector(1 downto 0);
    signal VN968_in0 : std_logic_vector(1 downto 0);
    signal VN968_in1 : std_logic_vector(1 downto 0);
    signal VN968_in2 : std_logic_vector(1 downto 0);
    signal VN968_in3 : std_logic_vector(1 downto 0);
    signal VN968_in4 : std_logic_vector(1 downto 0);
    signal VN968_in5 : std_logic_vector(1 downto 0);
    signal VN969_in0 : std_logic_vector(1 downto 0);
    signal VN969_in1 : std_logic_vector(1 downto 0);
    signal VN969_in2 : std_logic_vector(1 downto 0);
    signal VN969_in3 : std_logic_vector(1 downto 0);
    signal VN969_in4 : std_logic_vector(1 downto 0);
    signal VN969_in5 : std_logic_vector(1 downto 0);
    signal VN970_in0 : std_logic_vector(1 downto 0);
    signal VN970_in1 : std_logic_vector(1 downto 0);
    signal VN970_in2 : std_logic_vector(1 downto 0);
    signal VN970_in3 : std_logic_vector(1 downto 0);
    signal VN970_in4 : std_logic_vector(1 downto 0);
    signal VN970_in5 : std_logic_vector(1 downto 0);
    signal VN971_in0 : std_logic_vector(1 downto 0);
    signal VN971_in1 : std_logic_vector(1 downto 0);
    signal VN971_in2 : std_logic_vector(1 downto 0);
    signal VN971_in3 : std_logic_vector(1 downto 0);
    signal VN971_in4 : std_logic_vector(1 downto 0);
    signal VN971_in5 : std_logic_vector(1 downto 0);
    signal VN972_in0 : std_logic_vector(1 downto 0);
    signal VN972_in1 : std_logic_vector(1 downto 0);
    signal VN972_in2 : std_logic_vector(1 downto 0);
    signal VN972_in3 : std_logic_vector(1 downto 0);
    signal VN972_in4 : std_logic_vector(1 downto 0);
    signal VN972_in5 : std_logic_vector(1 downto 0);
    signal VN973_in0 : std_logic_vector(1 downto 0);
    signal VN973_in1 : std_logic_vector(1 downto 0);
    signal VN973_in2 : std_logic_vector(1 downto 0);
    signal VN973_in3 : std_logic_vector(1 downto 0);
    signal VN973_in4 : std_logic_vector(1 downto 0);
    signal VN973_in5 : std_logic_vector(1 downto 0);
    signal VN974_in0 : std_logic_vector(1 downto 0);
    signal VN974_in1 : std_logic_vector(1 downto 0);
    signal VN974_in2 : std_logic_vector(1 downto 0);
    signal VN974_in3 : std_logic_vector(1 downto 0);
    signal VN974_in4 : std_logic_vector(1 downto 0);
    signal VN974_in5 : std_logic_vector(1 downto 0);
    signal VN975_in0 : std_logic_vector(1 downto 0);
    signal VN975_in1 : std_logic_vector(1 downto 0);
    signal VN975_in2 : std_logic_vector(1 downto 0);
    signal VN975_in3 : std_logic_vector(1 downto 0);
    signal VN975_in4 : std_logic_vector(1 downto 0);
    signal VN975_in5 : std_logic_vector(1 downto 0);
    signal VN976_in0 : std_logic_vector(1 downto 0);
    signal VN976_in1 : std_logic_vector(1 downto 0);
    signal VN976_in2 : std_logic_vector(1 downto 0);
    signal VN976_in3 : std_logic_vector(1 downto 0);
    signal VN976_in4 : std_logic_vector(1 downto 0);
    signal VN976_in5 : std_logic_vector(1 downto 0);
    signal VN977_in0 : std_logic_vector(1 downto 0);
    signal VN977_in1 : std_logic_vector(1 downto 0);
    signal VN977_in2 : std_logic_vector(1 downto 0);
    signal VN977_in3 : std_logic_vector(1 downto 0);
    signal VN977_in4 : std_logic_vector(1 downto 0);
    signal VN977_in5 : std_logic_vector(1 downto 0);
    signal VN978_in0 : std_logic_vector(1 downto 0);
    signal VN978_in1 : std_logic_vector(1 downto 0);
    signal VN978_in2 : std_logic_vector(1 downto 0);
    signal VN978_in3 : std_logic_vector(1 downto 0);
    signal VN978_in4 : std_logic_vector(1 downto 0);
    signal VN978_in5 : std_logic_vector(1 downto 0);
    signal VN979_in0 : std_logic_vector(1 downto 0);
    signal VN979_in1 : std_logic_vector(1 downto 0);
    signal VN979_in2 : std_logic_vector(1 downto 0);
    signal VN979_in3 : std_logic_vector(1 downto 0);
    signal VN979_in4 : std_logic_vector(1 downto 0);
    signal VN979_in5 : std_logic_vector(1 downto 0);
    signal VN980_in0 : std_logic_vector(1 downto 0);
    signal VN980_in1 : std_logic_vector(1 downto 0);
    signal VN980_in2 : std_logic_vector(1 downto 0);
    signal VN980_in3 : std_logic_vector(1 downto 0);
    signal VN980_in4 : std_logic_vector(1 downto 0);
    signal VN980_in5 : std_logic_vector(1 downto 0);
    signal VN981_in0 : std_logic_vector(1 downto 0);
    signal VN981_in1 : std_logic_vector(1 downto 0);
    signal VN981_in2 : std_logic_vector(1 downto 0);
    signal VN981_in3 : std_logic_vector(1 downto 0);
    signal VN981_in4 : std_logic_vector(1 downto 0);
    signal VN981_in5 : std_logic_vector(1 downto 0);
    signal VN982_in0 : std_logic_vector(1 downto 0);
    signal VN982_in1 : std_logic_vector(1 downto 0);
    signal VN982_in2 : std_logic_vector(1 downto 0);
    signal VN982_in3 : std_logic_vector(1 downto 0);
    signal VN982_in4 : std_logic_vector(1 downto 0);
    signal VN982_in5 : std_logic_vector(1 downto 0);
    signal VN983_in0 : std_logic_vector(1 downto 0);
    signal VN983_in1 : std_logic_vector(1 downto 0);
    signal VN983_in2 : std_logic_vector(1 downto 0);
    signal VN983_in3 : std_logic_vector(1 downto 0);
    signal VN983_in4 : std_logic_vector(1 downto 0);
    signal VN983_in5 : std_logic_vector(1 downto 0);
    signal VN984_in0 : std_logic_vector(1 downto 0);
    signal VN984_in1 : std_logic_vector(1 downto 0);
    signal VN984_in2 : std_logic_vector(1 downto 0);
    signal VN984_in3 : std_logic_vector(1 downto 0);
    signal VN984_in4 : std_logic_vector(1 downto 0);
    signal VN984_in5 : std_logic_vector(1 downto 0);
    signal VN985_in0 : std_logic_vector(1 downto 0);
    signal VN985_in1 : std_logic_vector(1 downto 0);
    signal VN985_in2 : std_logic_vector(1 downto 0);
    signal VN985_in3 : std_logic_vector(1 downto 0);
    signal VN985_in4 : std_logic_vector(1 downto 0);
    signal VN985_in5 : std_logic_vector(1 downto 0);
    signal VN986_in0 : std_logic_vector(1 downto 0);
    signal VN986_in1 : std_logic_vector(1 downto 0);
    signal VN986_in2 : std_logic_vector(1 downto 0);
    signal VN986_in3 : std_logic_vector(1 downto 0);
    signal VN986_in4 : std_logic_vector(1 downto 0);
    signal VN986_in5 : std_logic_vector(1 downto 0);
    signal VN987_in0 : std_logic_vector(1 downto 0);
    signal VN987_in1 : std_logic_vector(1 downto 0);
    signal VN987_in2 : std_logic_vector(1 downto 0);
    signal VN987_in3 : std_logic_vector(1 downto 0);
    signal VN987_in4 : std_logic_vector(1 downto 0);
    signal VN987_in5 : std_logic_vector(1 downto 0);
    signal VN988_in0 : std_logic_vector(1 downto 0);
    signal VN988_in1 : std_logic_vector(1 downto 0);
    signal VN988_in2 : std_logic_vector(1 downto 0);
    signal VN988_in3 : std_logic_vector(1 downto 0);
    signal VN988_in4 : std_logic_vector(1 downto 0);
    signal VN988_in5 : std_logic_vector(1 downto 0);
    signal VN989_in0 : std_logic_vector(1 downto 0);
    signal VN989_in1 : std_logic_vector(1 downto 0);
    signal VN989_in2 : std_logic_vector(1 downto 0);
    signal VN989_in3 : std_logic_vector(1 downto 0);
    signal VN989_in4 : std_logic_vector(1 downto 0);
    signal VN989_in5 : std_logic_vector(1 downto 0);
    signal VN990_in0 : std_logic_vector(1 downto 0);
    signal VN990_in1 : std_logic_vector(1 downto 0);
    signal VN990_in2 : std_logic_vector(1 downto 0);
    signal VN990_in3 : std_logic_vector(1 downto 0);
    signal VN990_in4 : std_logic_vector(1 downto 0);
    signal VN990_in5 : std_logic_vector(1 downto 0);
    signal VN991_in0 : std_logic_vector(1 downto 0);
    signal VN991_in1 : std_logic_vector(1 downto 0);
    signal VN991_in2 : std_logic_vector(1 downto 0);
    signal VN991_in3 : std_logic_vector(1 downto 0);
    signal VN991_in4 : std_logic_vector(1 downto 0);
    signal VN991_in5 : std_logic_vector(1 downto 0);
    signal VN992_in0 : std_logic_vector(1 downto 0);
    signal VN992_in1 : std_logic_vector(1 downto 0);
    signal VN992_in2 : std_logic_vector(1 downto 0);
    signal VN992_in3 : std_logic_vector(1 downto 0);
    signal VN992_in4 : std_logic_vector(1 downto 0);
    signal VN992_in5 : std_logic_vector(1 downto 0);
    signal VN993_in0 : std_logic_vector(1 downto 0);
    signal VN993_in1 : std_logic_vector(1 downto 0);
    signal VN993_in2 : std_logic_vector(1 downto 0);
    signal VN993_in3 : std_logic_vector(1 downto 0);
    signal VN993_in4 : std_logic_vector(1 downto 0);
    signal VN993_in5 : std_logic_vector(1 downto 0);
    signal VN994_in0 : std_logic_vector(1 downto 0);
    signal VN994_in1 : std_logic_vector(1 downto 0);
    signal VN994_in2 : std_logic_vector(1 downto 0);
    signal VN994_in3 : std_logic_vector(1 downto 0);
    signal VN994_in4 : std_logic_vector(1 downto 0);
    signal VN994_in5 : std_logic_vector(1 downto 0);
    signal VN995_in0 : std_logic_vector(1 downto 0);
    signal VN995_in1 : std_logic_vector(1 downto 0);
    signal VN995_in2 : std_logic_vector(1 downto 0);
    signal VN995_in3 : std_logic_vector(1 downto 0);
    signal VN995_in4 : std_logic_vector(1 downto 0);
    signal VN995_in5 : std_logic_vector(1 downto 0);
    signal VN996_in0 : std_logic_vector(1 downto 0);
    signal VN996_in1 : std_logic_vector(1 downto 0);
    signal VN996_in2 : std_logic_vector(1 downto 0);
    signal VN996_in3 : std_logic_vector(1 downto 0);
    signal VN996_in4 : std_logic_vector(1 downto 0);
    signal VN996_in5 : std_logic_vector(1 downto 0);
    signal VN997_in0 : std_logic_vector(1 downto 0);
    signal VN997_in1 : std_logic_vector(1 downto 0);
    signal VN997_in2 : std_logic_vector(1 downto 0);
    signal VN997_in3 : std_logic_vector(1 downto 0);
    signal VN997_in4 : std_logic_vector(1 downto 0);
    signal VN997_in5 : std_logic_vector(1 downto 0);
    signal VN998_in0 : std_logic_vector(1 downto 0);
    signal VN998_in1 : std_logic_vector(1 downto 0);
    signal VN998_in2 : std_logic_vector(1 downto 0);
    signal VN998_in3 : std_logic_vector(1 downto 0);
    signal VN998_in4 : std_logic_vector(1 downto 0);
    signal VN998_in5 : std_logic_vector(1 downto 0);
    signal VN999_in0 : std_logic_vector(1 downto 0);
    signal VN999_in1 : std_logic_vector(1 downto 0);
    signal VN999_in2 : std_logic_vector(1 downto 0);
    signal VN999_in3 : std_logic_vector(1 downto 0);
    signal VN999_in4 : std_logic_vector(1 downto 0);
    signal VN999_in5 : std_logic_vector(1 downto 0);
    signal VN1000_in0 : std_logic_vector(1 downto 0);
    signal VN1000_in1 : std_logic_vector(1 downto 0);
    signal VN1000_in2 : std_logic_vector(1 downto 0);
    signal VN1000_in3 : std_logic_vector(1 downto 0);
    signal VN1000_in4 : std_logic_vector(1 downto 0);
    signal VN1000_in5 : std_logic_vector(1 downto 0);
    signal VN1001_in0 : std_logic_vector(1 downto 0);
    signal VN1001_in1 : std_logic_vector(1 downto 0);
    signal VN1001_in2 : std_logic_vector(1 downto 0);
    signal VN1001_in3 : std_logic_vector(1 downto 0);
    signal VN1001_in4 : std_logic_vector(1 downto 0);
    signal VN1001_in5 : std_logic_vector(1 downto 0);
    signal VN1002_in0 : std_logic_vector(1 downto 0);
    signal VN1002_in1 : std_logic_vector(1 downto 0);
    signal VN1002_in2 : std_logic_vector(1 downto 0);
    signal VN1002_in3 : std_logic_vector(1 downto 0);
    signal VN1002_in4 : std_logic_vector(1 downto 0);
    signal VN1002_in5 : std_logic_vector(1 downto 0);
    signal VN1003_in0 : std_logic_vector(1 downto 0);
    signal VN1003_in1 : std_logic_vector(1 downto 0);
    signal VN1003_in2 : std_logic_vector(1 downto 0);
    signal VN1003_in3 : std_logic_vector(1 downto 0);
    signal VN1003_in4 : std_logic_vector(1 downto 0);
    signal VN1003_in5 : std_logic_vector(1 downto 0);
    signal VN1004_in0 : std_logic_vector(1 downto 0);
    signal VN1004_in1 : std_logic_vector(1 downto 0);
    signal VN1004_in2 : std_logic_vector(1 downto 0);
    signal VN1004_in3 : std_logic_vector(1 downto 0);
    signal VN1004_in4 : std_logic_vector(1 downto 0);
    signal VN1004_in5 : std_logic_vector(1 downto 0);
    signal VN1005_in0 : std_logic_vector(1 downto 0);
    signal VN1005_in1 : std_logic_vector(1 downto 0);
    signal VN1005_in2 : std_logic_vector(1 downto 0);
    signal VN1005_in3 : std_logic_vector(1 downto 0);
    signal VN1005_in4 : std_logic_vector(1 downto 0);
    signal VN1005_in5 : std_logic_vector(1 downto 0);
    signal VN1006_in0 : std_logic_vector(1 downto 0);
    signal VN1006_in1 : std_logic_vector(1 downto 0);
    signal VN1006_in2 : std_logic_vector(1 downto 0);
    signal VN1006_in3 : std_logic_vector(1 downto 0);
    signal VN1006_in4 : std_logic_vector(1 downto 0);
    signal VN1006_in5 : std_logic_vector(1 downto 0);
    signal VN1007_in0 : std_logic_vector(1 downto 0);
    signal VN1007_in1 : std_logic_vector(1 downto 0);
    signal VN1007_in2 : std_logic_vector(1 downto 0);
    signal VN1007_in3 : std_logic_vector(1 downto 0);
    signal VN1007_in4 : std_logic_vector(1 downto 0);
    signal VN1007_in5 : std_logic_vector(1 downto 0);
    signal VN1008_in0 : std_logic_vector(1 downto 0);
    signal VN1008_in1 : std_logic_vector(1 downto 0);
    signal VN1008_in2 : std_logic_vector(1 downto 0);
    signal VN1008_in3 : std_logic_vector(1 downto 0);
    signal VN1008_in4 : std_logic_vector(1 downto 0);
    signal VN1008_in5 : std_logic_vector(1 downto 0);
    signal VN1009_in0 : std_logic_vector(1 downto 0);
    signal VN1009_in1 : std_logic_vector(1 downto 0);
    signal VN1009_in2 : std_logic_vector(1 downto 0);
    signal VN1009_in3 : std_logic_vector(1 downto 0);
    signal VN1009_in4 : std_logic_vector(1 downto 0);
    signal VN1009_in5 : std_logic_vector(1 downto 0);
    signal VN1010_in0 : std_logic_vector(1 downto 0);
    signal VN1010_in1 : std_logic_vector(1 downto 0);
    signal VN1010_in2 : std_logic_vector(1 downto 0);
    signal VN1010_in3 : std_logic_vector(1 downto 0);
    signal VN1010_in4 : std_logic_vector(1 downto 0);
    signal VN1010_in5 : std_logic_vector(1 downto 0);
    signal VN1011_in0 : std_logic_vector(1 downto 0);
    signal VN1011_in1 : std_logic_vector(1 downto 0);
    signal VN1011_in2 : std_logic_vector(1 downto 0);
    signal VN1011_in3 : std_logic_vector(1 downto 0);
    signal VN1011_in4 : std_logic_vector(1 downto 0);
    signal VN1011_in5 : std_logic_vector(1 downto 0);
    signal VN1012_in0 : std_logic_vector(1 downto 0);
    signal VN1012_in1 : std_logic_vector(1 downto 0);
    signal VN1012_in2 : std_logic_vector(1 downto 0);
    signal VN1012_in3 : std_logic_vector(1 downto 0);
    signal VN1012_in4 : std_logic_vector(1 downto 0);
    signal VN1012_in5 : std_logic_vector(1 downto 0);
    signal VN1013_in0 : std_logic_vector(1 downto 0);
    signal VN1013_in1 : std_logic_vector(1 downto 0);
    signal VN1013_in2 : std_logic_vector(1 downto 0);
    signal VN1013_in3 : std_logic_vector(1 downto 0);
    signal VN1013_in4 : std_logic_vector(1 downto 0);
    signal VN1013_in5 : std_logic_vector(1 downto 0);
    signal VN1014_in0 : std_logic_vector(1 downto 0);
    signal VN1014_in1 : std_logic_vector(1 downto 0);
    signal VN1014_in2 : std_logic_vector(1 downto 0);
    signal VN1014_in3 : std_logic_vector(1 downto 0);
    signal VN1014_in4 : std_logic_vector(1 downto 0);
    signal VN1014_in5 : std_logic_vector(1 downto 0);
    signal VN1015_in0 : std_logic_vector(1 downto 0);
    signal VN1015_in1 : std_logic_vector(1 downto 0);
    signal VN1015_in2 : std_logic_vector(1 downto 0);
    signal VN1015_in3 : std_logic_vector(1 downto 0);
    signal VN1015_in4 : std_logic_vector(1 downto 0);
    signal VN1015_in5 : std_logic_vector(1 downto 0);
    signal VN1016_in0 : std_logic_vector(1 downto 0);
    signal VN1016_in1 : std_logic_vector(1 downto 0);
    signal VN1016_in2 : std_logic_vector(1 downto 0);
    signal VN1016_in3 : std_logic_vector(1 downto 0);
    signal VN1016_in4 : std_logic_vector(1 downto 0);
    signal VN1016_in5 : std_logic_vector(1 downto 0);
    signal VN1017_in0 : std_logic_vector(1 downto 0);
    signal VN1017_in1 : std_logic_vector(1 downto 0);
    signal VN1017_in2 : std_logic_vector(1 downto 0);
    signal VN1017_in3 : std_logic_vector(1 downto 0);
    signal VN1017_in4 : std_logic_vector(1 downto 0);
    signal VN1017_in5 : std_logic_vector(1 downto 0);
    signal VN1018_in0 : std_logic_vector(1 downto 0);
    signal VN1018_in1 : std_logic_vector(1 downto 0);
    signal VN1018_in2 : std_logic_vector(1 downto 0);
    signal VN1018_in3 : std_logic_vector(1 downto 0);
    signal VN1018_in4 : std_logic_vector(1 downto 0);
    signal VN1018_in5 : std_logic_vector(1 downto 0);
    signal VN1019_in0 : std_logic_vector(1 downto 0);
    signal VN1019_in1 : std_logic_vector(1 downto 0);
    signal VN1019_in2 : std_logic_vector(1 downto 0);
    signal VN1019_in3 : std_logic_vector(1 downto 0);
    signal VN1019_in4 : std_logic_vector(1 downto 0);
    signal VN1019_in5 : std_logic_vector(1 downto 0);
    signal VN1020_in0 : std_logic_vector(1 downto 0);
    signal VN1020_in1 : std_logic_vector(1 downto 0);
    signal VN1020_in2 : std_logic_vector(1 downto 0);
    signal VN1020_in3 : std_logic_vector(1 downto 0);
    signal VN1020_in4 : std_logic_vector(1 downto 0);
    signal VN1020_in5 : std_logic_vector(1 downto 0);
    signal VN1021_in0 : std_logic_vector(1 downto 0);
    signal VN1021_in1 : std_logic_vector(1 downto 0);
    signal VN1021_in2 : std_logic_vector(1 downto 0);
    signal VN1021_in3 : std_logic_vector(1 downto 0);
    signal VN1021_in4 : std_logic_vector(1 downto 0);
    signal VN1021_in5 : std_logic_vector(1 downto 0);
    signal VN1022_in0 : std_logic_vector(1 downto 0);
    signal VN1022_in1 : std_logic_vector(1 downto 0);
    signal VN1022_in2 : std_logic_vector(1 downto 0);
    signal VN1022_in3 : std_logic_vector(1 downto 0);
    signal VN1022_in4 : std_logic_vector(1 downto 0);
    signal VN1022_in5 : std_logic_vector(1 downto 0);
    signal VN1023_in0 : std_logic_vector(1 downto 0);
    signal VN1023_in1 : std_logic_vector(1 downto 0);
    signal VN1023_in2 : std_logic_vector(1 downto 0);
    signal VN1023_in3 : std_logic_vector(1 downto 0);
    signal VN1023_in4 : std_logic_vector(1 downto 0);
    signal VN1023_in5 : std_logic_vector(1 downto 0);
    signal VN1024_in0 : std_logic_vector(1 downto 0);
    signal VN1024_in1 : std_logic_vector(1 downto 0);
    signal VN1024_in2 : std_logic_vector(1 downto 0);
    signal VN1024_in3 : std_logic_vector(1 downto 0);
    signal VN1024_in4 : std_logic_vector(1 downto 0);
    signal VN1024_in5 : std_logic_vector(1 downto 0);
    signal VN1025_in0 : std_logic_vector(1 downto 0);
    signal VN1025_in1 : std_logic_vector(1 downto 0);
    signal VN1025_in2 : std_logic_vector(1 downto 0);
    signal VN1025_in3 : std_logic_vector(1 downto 0);
    signal VN1025_in4 : std_logic_vector(1 downto 0);
    signal VN1025_in5 : std_logic_vector(1 downto 0);
    signal VN1026_in0 : std_logic_vector(1 downto 0);
    signal VN1026_in1 : std_logic_vector(1 downto 0);
    signal VN1026_in2 : std_logic_vector(1 downto 0);
    signal VN1026_in3 : std_logic_vector(1 downto 0);
    signal VN1026_in4 : std_logic_vector(1 downto 0);
    signal VN1026_in5 : std_logic_vector(1 downto 0);
    signal VN1027_in0 : std_logic_vector(1 downto 0);
    signal VN1027_in1 : std_logic_vector(1 downto 0);
    signal VN1027_in2 : std_logic_vector(1 downto 0);
    signal VN1027_in3 : std_logic_vector(1 downto 0);
    signal VN1027_in4 : std_logic_vector(1 downto 0);
    signal VN1027_in5 : std_logic_vector(1 downto 0);
    signal VN1028_in0 : std_logic_vector(1 downto 0);
    signal VN1028_in1 : std_logic_vector(1 downto 0);
    signal VN1028_in2 : std_logic_vector(1 downto 0);
    signal VN1028_in3 : std_logic_vector(1 downto 0);
    signal VN1028_in4 : std_logic_vector(1 downto 0);
    signal VN1028_in5 : std_logic_vector(1 downto 0);
    signal VN1029_in0 : std_logic_vector(1 downto 0);
    signal VN1029_in1 : std_logic_vector(1 downto 0);
    signal VN1029_in2 : std_logic_vector(1 downto 0);
    signal VN1029_in3 : std_logic_vector(1 downto 0);
    signal VN1029_in4 : std_logic_vector(1 downto 0);
    signal VN1029_in5 : std_logic_vector(1 downto 0);
    signal VN1030_in0 : std_logic_vector(1 downto 0);
    signal VN1030_in1 : std_logic_vector(1 downto 0);
    signal VN1030_in2 : std_logic_vector(1 downto 0);
    signal VN1030_in3 : std_logic_vector(1 downto 0);
    signal VN1030_in4 : std_logic_vector(1 downto 0);
    signal VN1030_in5 : std_logic_vector(1 downto 0);
    signal VN1031_in0 : std_logic_vector(1 downto 0);
    signal VN1031_in1 : std_logic_vector(1 downto 0);
    signal VN1031_in2 : std_logic_vector(1 downto 0);
    signal VN1031_in3 : std_logic_vector(1 downto 0);
    signal VN1031_in4 : std_logic_vector(1 downto 0);
    signal VN1031_in5 : std_logic_vector(1 downto 0);
    signal VN1032_in0 : std_logic_vector(1 downto 0);
    signal VN1032_in1 : std_logic_vector(1 downto 0);
    signal VN1032_in2 : std_logic_vector(1 downto 0);
    signal VN1032_in3 : std_logic_vector(1 downto 0);
    signal VN1032_in4 : std_logic_vector(1 downto 0);
    signal VN1032_in5 : std_logic_vector(1 downto 0);
    signal VN1033_in0 : std_logic_vector(1 downto 0);
    signal VN1033_in1 : std_logic_vector(1 downto 0);
    signal VN1033_in2 : std_logic_vector(1 downto 0);
    signal VN1033_in3 : std_logic_vector(1 downto 0);
    signal VN1033_in4 : std_logic_vector(1 downto 0);
    signal VN1033_in5 : std_logic_vector(1 downto 0);
    signal VN1034_in0 : std_logic_vector(1 downto 0);
    signal VN1034_in1 : std_logic_vector(1 downto 0);
    signal VN1034_in2 : std_logic_vector(1 downto 0);
    signal VN1034_in3 : std_logic_vector(1 downto 0);
    signal VN1034_in4 : std_logic_vector(1 downto 0);
    signal VN1034_in5 : std_logic_vector(1 downto 0);
    signal VN1035_in0 : std_logic_vector(1 downto 0);
    signal VN1035_in1 : std_logic_vector(1 downto 0);
    signal VN1035_in2 : std_logic_vector(1 downto 0);
    signal VN1035_in3 : std_logic_vector(1 downto 0);
    signal VN1035_in4 : std_logic_vector(1 downto 0);
    signal VN1035_in5 : std_logic_vector(1 downto 0);
    signal VN1036_in0 : std_logic_vector(1 downto 0);
    signal VN1036_in1 : std_logic_vector(1 downto 0);
    signal VN1036_in2 : std_logic_vector(1 downto 0);
    signal VN1036_in3 : std_logic_vector(1 downto 0);
    signal VN1036_in4 : std_logic_vector(1 downto 0);
    signal VN1036_in5 : std_logic_vector(1 downto 0);
    signal VN1037_in0 : std_logic_vector(1 downto 0);
    signal VN1037_in1 : std_logic_vector(1 downto 0);
    signal VN1037_in2 : std_logic_vector(1 downto 0);
    signal VN1037_in3 : std_logic_vector(1 downto 0);
    signal VN1037_in4 : std_logic_vector(1 downto 0);
    signal VN1037_in5 : std_logic_vector(1 downto 0);
    signal VN1038_in0 : std_logic_vector(1 downto 0);
    signal VN1038_in1 : std_logic_vector(1 downto 0);
    signal VN1038_in2 : std_logic_vector(1 downto 0);
    signal VN1038_in3 : std_logic_vector(1 downto 0);
    signal VN1038_in4 : std_logic_vector(1 downto 0);
    signal VN1038_in5 : std_logic_vector(1 downto 0);
    signal VN1039_in0 : std_logic_vector(1 downto 0);
    signal VN1039_in1 : std_logic_vector(1 downto 0);
    signal VN1039_in2 : std_logic_vector(1 downto 0);
    signal VN1039_in3 : std_logic_vector(1 downto 0);
    signal VN1039_in4 : std_logic_vector(1 downto 0);
    signal VN1039_in5 : std_logic_vector(1 downto 0);
    signal VN1040_in0 : std_logic_vector(1 downto 0);
    signal VN1040_in1 : std_logic_vector(1 downto 0);
    signal VN1040_in2 : std_logic_vector(1 downto 0);
    signal VN1040_in3 : std_logic_vector(1 downto 0);
    signal VN1040_in4 : std_logic_vector(1 downto 0);
    signal VN1040_in5 : std_logic_vector(1 downto 0);
    signal VN1041_in0 : std_logic_vector(1 downto 0);
    signal VN1041_in1 : std_logic_vector(1 downto 0);
    signal VN1041_in2 : std_logic_vector(1 downto 0);
    signal VN1041_in3 : std_logic_vector(1 downto 0);
    signal VN1041_in4 : std_logic_vector(1 downto 0);
    signal VN1041_in5 : std_logic_vector(1 downto 0);
    signal VN1042_in0 : std_logic_vector(1 downto 0);
    signal VN1042_in1 : std_logic_vector(1 downto 0);
    signal VN1042_in2 : std_logic_vector(1 downto 0);
    signal VN1042_in3 : std_logic_vector(1 downto 0);
    signal VN1042_in4 : std_logic_vector(1 downto 0);
    signal VN1042_in5 : std_logic_vector(1 downto 0);
    signal VN1043_in0 : std_logic_vector(1 downto 0);
    signal VN1043_in1 : std_logic_vector(1 downto 0);
    signal VN1043_in2 : std_logic_vector(1 downto 0);
    signal VN1043_in3 : std_logic_vector(1 downto 0);
    signal VN1043_in4 : std_logic_vector(1 downto 0);
    signal VN1043_in5 : std_logic_vector(1 downto 0);
    signal VN1044_in0 : std_logic_vector(1 downto 0);
    signal VN1044_in1 : std_logic_vector(1 downto 0);
    signal VN1044_in2 : std_logic_vector(1 downto 0);
    signal VN1044_in3 : std_logic_vector(1 downto 0);
    signal VN1044_in4 : std_logic_vector(1 downto 0);
    signal VN1044_in5 : std_logic_vector(1 downto 0);
    signal VN1045_in0 : std_logic_vector(1 downto 0);
    signal VN1045_in1 : std_logic_vector(1 downto 0);
    signal VN1045_in2 : std_logic_vector(1 downto 0);
    signal VN1045_in3 : std_logic_vector(1 downto 0);
    signal VN1045_in4 : std_logic_vector(1 downto 0);
    signal VN1045_in5 : std_logic_vector(1 downto 0);
    signal VN1046_in0 : std_logic_vector(1 downto 0);
    signal VN1046_in1 : std_logic_vector(1 downto 0);
    signal VN1046_in2 : std_logic_vector(1 downto 0);
    signal VN1046_in3 : std_logic_vector(1 downto 0);
    signal VN1046_in4 : std_logic_vector(1 downto 0);
    signal VN1046_in5 : std_logic_vector(1 downto 0);
    signal VN1047_in0 : std_logic_vector(1 downto 0);
    signal VN1047_in1 : std_logic_vector(1 downto 0);
    signal VN1047_in2 : std_logic_vector(1 downto 0);
    signal VN1047_in3 : std_logic_vector(1 downto 0);
    signal VN1047_in4 : std_logic_vector(1 downto 0);
    signal VN1047_in5 : std_logic_vector(1 downto 0);
    signal VN1048_in0 : std_logic_vector(1 downto 0);
    signal VN1048_in1 : std_logic_vector(1 downto 0);
    signal VN1048_in2 : std_logic_vector(1 downto 0);
    signal VN1048_in3 : std_logic_vector(1 downto 0);
    signal VN1048_in4 : std_logic_vector(1 downto 0);
    signal VN1048_in5 : std_logic_vector(1 downto 0);
    signal VN1049_in0 : std_logic_vector(1 downto 0);
    signal VN1049_in1 : std_logic_vector(1 downto 0);
    signal VN1049_in2 : std_logic_vector(1 downto 0);
    signal VN1049_in3 : std_logic_vector(1 downto 0);
    signal VN1049_in4 : std_logic_vector(1 downto 0);
    signal VN1049_in5 : std_logic_vector(1 downto 0);
    signal VN1050_in0 : std_logic_vector(1 downto 0);
    signal VN1050_in1 : std_logic_vector(1 downto 0);
    signal VN1050_in2 : std_logic_vector(1 downto 0);
    signal VN1050_in3 : std_logic_vector(1 downto 0);
    signal VN1050_in4 : std_logic_vector(1 downto 0);
    signal VN1050_in5 : std_logic_vector(1 downto 0);
    signal VN1051_in0 : std_logic_vector(1 downto 0);
    signal VN1051_in1 : std_logic_vector(1 downto 0);
    signal VN1051_in2 : std_logic_vector(1 downto 0);
    signal VN1051_in3 : std_logic_vector(1 downto 0);
    signal VN1051_in4 : std_logic_vector(1 downto 0);
    signal VN1051_in5 : std_logic_vector(1 downto 0);
    signal VN1052_in0 : std_logic_vector(1 downto 0);
    signal VN1052_in1 : std_logic_vector(1 downto 0);
    signal VN1052_in2 : std_logic_vector(1 downto 0);
    signal VN1052_in3 : std_logic_vector(1 downto 0);
    signal VN1052_in4 : std_logic_vector(1 downto 0);
    signal VN1052_in5 : std_logic_vector(1 downto 0);
    signal VN1053_in0 : std_logic_vector(1 downto 0);
    signal VN1053_in1 : std_logic_vector(1 downto 0);
    signal VN1053_in2 : std_logic_vector(1 downto 0);
    signal VN1053_in3 : std_logic_vector(1 downto 0);
    signal VN1053_in4 : std_logic_vector(1 downto 0);
    signal VN1053_in5 : std_logic_vector(1 downto 0);
    signal VN1054_in0 : std_logic_vector(1 downto 0);
    signal VN1054_in1 : std_logic_vector(1 downto 0);
    signal VN1054_in2 : std_logic_vector(1 downto 0);
    signal VN1054_in3 : std_logic_vector(1 downto 0);
    signal VN1054_in4 : std_logic_vector(1 downto 0);
    signal VN1054_in5 : std_logic_vector(1 downto 0);
    signal VN1055_in0 : std_logic_vector(1 downto 0);
    signal VN1055_in1 : std_logic_vector(1 downto 0);
    signal VN1055_in2 : std_logic_vector(1 downto 0);
    signal VN1055_in3 : std_logic_vector(1 downto 0);
    signal VN1055_in4 : std_logic_vector(1 downto 0);
    signal VN1055_in5 : std_logic_vector(1 downto 0);
    signal VN1056_in0 : std_logic_vector(1 downto 0);
    signal VN1056_in1 : std_logic_vector(1 downto 0);
    signal VN1056_in2 : std_logic_vector(1 downto 0);
    signal VN1056_in3 : std_logic_vector(1 downto 0);
    signal VN1056_in4 : std_logic_vector(1 downto 0);
    signal VN1056_in5 : std_logic_vector(1 downto 0);
    signal VN1057_in0 : std_logic_vector(1 downto 0);
    signal VN1057_in1 : std_logic_vector(1 downto 0);
    signal VN1057_in2 : std_logic_vector(1 downto 0);
    signal VN1057_in3 : std_logic_vector(1 downto 0);
    signal VN1057_in4 : std_logic_vector(1 downto 0);
    signal VN1057_in5 : std_logic_vector(1 downto 0);
    signal VN1058_in0 : std_logic_vector(1 downto 0);
    signal VN1058_in1 : std_logic_vector(1 downto 0);
    signal VN1058_in2 : std_logic_vector(1 downto 0);
    signal VN1058_in3 : std_logic_vector(1 downto 0);
    signal VN1058_in4 : std_logic_vector(1 downto 0);
    signal VN1058_in5 : std_logic_vector(1 downto 0);
    signal VN1059_in0 : std_logic_vector(1 downto 0);
    signal VN1059_in1 : std_logic_vector(1 downto 0);
    signal VN1059_in2 : std_logic_vector(1 downto 0);
    signal VN1059_in3 : std_logic_vector(1 downto 0);
    signal VN1059_in4 : std_logic_vector(1 downto 0);
    signal VN1059_in5 : std_logic_vector(1 downto 0);
    signal VN1060_in0 : std_logic_vector(1 downto 0);
    signal VN1060_in1 : std_logic_vector(1 downto 0);
    signal VN1060_in2 : std_logic_vector(1 downto 0);
    signal VN1060_in3 : std_logic_vector(1 downto 0);
    signal VN1060_in4 : std_logic_vector(1 downto 0);
    signal VN1060_in5 : std_logic_vector(1 downto 0);
    signal VN1061_in0 : std_logic_vector(1 downto 0);
    signal VN1061_in1 : std_logic_vector(1 downto 0);
    signal VN1061_in2 : std_logic_vector(1 downto 0);
    signal VN1061_in3 : std_logic_vector(1 downto 0);
    signal VN1061_in4 : std_logic_vector(1 downto 0);
    signal VN1061_in5 : std_logic_vector(1 downto 0);
    signal VN1062_in0 : std_logic_vector(1 downto 0);
    signal VN1062_in1 : std_logic_vector(1 downto 0);
    signal VN1062_in2 : std_logic_vector(1 downto 0);
    signal VN1062_in3 : std_logic_vector(1 downto 0);
    signal VN1062_in4 : std_logic_vector(1 downto 0);
    signal VN1062_in5 : std_logic_vector(1 downto 0);
    signal VN1063_in0 : std_logic_vector(1 downto 0);
    signal VN1063_in1 : std_logic_vector(1 downto 0);
    signal VN1063_in2 : std_logic_vector(1 downto 0);
    signal VN1063_in3 : std_logic_vector(1 downto 0);
    signal VN1063_in4 : std_logic_vector(1 downto 0);
    signal VN1063_in5 : std_logic_vector(1 downto 0);
    signal VN1064_in0 : std_logic_vector(1 downto 0);
    signal VN1064_in1 : std_logic_vector(1 downto 0);
    signal VN1064_in2 : std_logic_vector(1 downto 0);
    signal VN1064_in3 : std_logic_vector(1 downto 0);
    signal VN1064_in4 : std_logic_vector(1 downto 0);
    signal VN1064_in5 : std_logic_vector(1 downto 0);
    signal VN1065_in0 : std_logic_vector(1 downto 0);
    signal VN1065_in1 : std_logic_vector(1 downto 0);
    signal VN1065_in2 : std_logic_vector(1 downto 0);
    signal VN1065_in3 : std_logic_vector(1 downto 0);
    signal VN1065_in4 : std_logic_vector(1 downto 0);
    signal VN1065_in5 : std_logic_vector(1 downto 0);
    signal VN1066_in0 : std_logic_vector(1 downto 0);
    signal VN1066_in1 : std_logic_vector(1 downto 0);
    signal VN1066_in2 : std_logic_vector(1 downto 0);
    signal VN1066_in3 : std_logic_vector(1 downto 0);
    signal VN1066_in4 : std_logic_vector(1 downto 0);
    signal VN1066_in5 : std_logic_vector(1 downto 0);
    signal VN1067_in0 : std_logic_vector(1 downto 0);
    signal VN1067_in1 : std_logic_vector(1 downto 0);
    signal VN1067_in2 : std_logic_vector(1 downto 0);
    signal VN1067_in3 : std_logic_vector(1 downto 0);
    signal VN1067_in4 : std_logic_vector(1 downto 0);
    signal VN1067_in5 : std_logic_vector(1 downto 0);
    signal VN1068_in0 : std_logic_vector(1 downto 0);
    signal VN1068_in1 : std_logic_vector(1 downto 0);
    signal VN1068_in2 : std_logic_vector(1 downto 0);
    signal VN1068_in3 : std_logic_vector(1 downto 0);
    signal VN1068_in4 : std_logic_vector(1 downto 0);
    signal VN1068_in5 : std_logic_vector(1 downto 0);
    signal VN1069_in0 : std_logic_vector(1 downto 0);
    signal VN1069_in1 : std_logic_vector(1 downto 0);
    signal VN1069_in2 : std_logic_vector(1 downto 0);
    signal VN1069_in3 : std_logic_vector(1 downto 0);
    signal VN1069_in4 : std_logic_vector(1 downto 0);
    signal VN1069_in5 : std_logic_vector(1 downto 0);
    signal VN1070_in0 : std_logic_vector(1 downto 0);
    signal VN1070_in1 : std_logic_vector(1 downto 0);
    signal VN1070_in2 : std_logic_vector(1 downto 0);
    signal VN1070_in3 : std_logic_vector(1 downto 0);
    signal VN1070_in4 : std_logic_vector(1 downto 0);
    signal VN1070_in5 : std_logic_vector(1 downto 0);
    signal VN1071_in0 : std_logic_vector(1 downto 0);
    signal VN1071_in1 : std_logic_vector(1 downto 0);
    signal VN1071_in2 : std_logic_vector(1 downto 0);
    signal VN1071_in3 : std_logic_vector(1 downto 0);
    signal VN1071_in4 : std_logic_vector(1 downto 0);
    signal VN1071_in5 : std_logic_vector(1 downto 0);
    signal VN1072_in0 : std_logic_vector(1 downto 0);
    signal VN1072_in1 : std_logic_vector(1 downto 0);
    signal VN1072_in2 : std_logic_vector(1 downto 0);
    signal VN1072_in3 : std_logic_vector(1 downto 0);
    signal VN1072_in4 : std_logic_vector(1 downto 0);
    signal VN1072_in5 : std_logic_vector(1 downto 0);
    signal VN1073_in0 : std_logic_vector(1 downto 0);
    signal VN1073_in1 : std_logic_vector(1 downto 0);
    signal VN1073_in2 : std_logic_vector(1 downto 0);
    signal VN1073_in3 : std_logic_vector(1 downto 0);
    signal VN1073_in4 : std_logic_vector(1 downto 0);
    signal VN1073_in5 : std_logic_vector(1 downto 0);
    signal VN1074_in0 : std_logic_vector(1 downto 0);
    signal VN1074_in1 : std_logic_vector(1 downto 0);
    signal VN1074_in2 : std_logic_vector(1 downto 0);
    signal VN1074_in3 : std_logic_vector(1 downto 0);
    signal VN1074_in4 : std_logic_vector(1 downto 0);
    signal VN1074_in5 : std_logic_vector(1 downto 0);
    signal VN1075_in0 : std_logic_vector(1 downto 0);
    signal VN1075_in1 : std_logic_vector(1 downto 0);
    signal VN1075_in2 : std_logic_vector(1 downto 0);
    signal VN1075_in3 : std_logic_vector(1 downto 0);
    signal VN1075_in4 : std_logic_vector(1 downto 0);
    signal VN1075_in5 : std_logic_vector(1 downto 0);
    signal VN1076_in0 : std_logic_vector(1 downto 0);
    signal VN1076_in1 : std_logic_vector(1 downto 0);
    signal VN1076_in2 : std_logic_vector(1 downto 0);
    signal VN1076_in3 : std_logic_vector(1 downto 0);
    signal VN1076_in4 : std_logic_vector(1 downto 0);
    signal VN1076_in5 : std_logic_vector(1 downto 0);
    signal VN1077_in0 : std_logic_vector(1 downto 0);
    signal VN1077_in1 : std_logic_vector(1 downto 0);
    signal VN1077_in2 : std_logic_vector(1 downto 0);
    signal VN1077_in3 : std_logic_vector(1 downto 0);
    signal VN1077_in4 : std_logic_vector(1 downto 0);
    signal VN1077_in5 : std_logic_vector(1 downto 0);
    signal VN1078_in0 : std_logic_vector(1 downto 0);
    signal VN1078_in1 : std_logic_vector(1 downto 0);
    signal VN1078_in2 : std_logic_vector(1 downto 0);
    signal VN1078_in3 : std_logic_vector(1 downto 0);
    signal VN1078_in4 : std_logic_vector(1 downto 0);
    signal VN1078_in5 : std_logic_vector(1 downto 0);
    signal VN1079_in0 : std_logic_vector(1 downto 0);
    signal VN1079_in1 : std_logic_vector(1 downto 0);
    signal VN1079_in2 : std_logic_vector(1 downto 0);
    signal VN1079_in3 : std_logic_vector(1 downto 0);
    signal VN1079_in4 : std_logic_vector(1 downto 0);
    signal VN1079_in5 : std_logic_vector(1 downto 0);
    signal VN1080_in0 : std_logic_vector(1 downto 0);
    signal VN1080_in1 : std_logic_vector(1 downto 0);
    signal VN1080_in2 : std_logic_vector(1 downto 0);
    signal VN1080_in3 : std_logic_vector(1 downto 0);
    signal VN1080_in4 : std_logic_vector(1 downto 0);
    signal VN1080_in5 : std_logic_vector(1 downto 0);
    signal VN1081_in0 : std_logic_vector(1 downto 0);
    signal VN1081_in1 : std_logic_vector(1 downto 0);
    signal VN1081_in2 : std_logic_vector(1 downto 0);
    signal VN1081_in3 : std_logic_vector(1 downto 0);
    signal VN1081_in4 : std_logic_vector(1 downto 0);
    signal VN1081_in5 : std_logic_vector(1 downto 0);
    signal VN1082_in0 : std_logic_vector(1 downto 0);
    signal VN1082_in1 : std_logic_vector(1 downto 0);
    signal VN1082_in2 : std_logic_vector(1 downto 0);
    signal VN1082_in3 : std_logic_vector(1 downto 0);
    signal VN1082_in4 : std_logic_vector(1 downto 0);
    signal VN1082_in5 : std_logic_vector(1 downto 0);
    signal VN1083_in0 : std_logic_vector(1 downto 0);
    signal VN1083_in1 : std_logic_vector(1 downto 0);
    signal VN1083_in2 : std_logic_vector(1 downto 0);
    signal VN1083_in3 : std_logic_vector(1 downto 0);
    signal VN1083_in4 : std_logic_vector(1 downto 0);
    signal VN1083_in5 : std_logic_vector(1 downto 0);
    signal VN1084_in0 : std_logic_vector(1 downto 0);
    signal VN1084_in1 : std_logic_vector(1 downto 0);
    signal VN1084_in2 : std_logic_vector(1 downto 0);
    signal VN1084_in3 : std_logic_vector(1 downto 0);
    signal VN1084_in4 : std_logic_vector(1 downto 0);
    signal VN1084_in5 : std_logic_vector(1 downto 0);
    signal VN1085_in0 : std_logic_vector(1 downto 0);
    signal VN1085_in1 : std_logic_vector(1 downto 0);
    signal VN1085_in2 : std_logic_vector(1 downto 0);
    signal VN1085_in3 : std_logic_vector(1 downto 0);
    signal VN1085_in4 : std_logic_vector(1 downto 0);
    signal VN1085_in5 : std_logic_vector(1 downto 0);
    signal VN1086_in0 : std_logic_vector(1 downto 0);
    signal VN1086_in1 : std_logic_vector(1 downto 0);
    signal VN1086_in2 : std_logic_vector(1 downto 0);
    signal VN1086_in3 : std_logic_vector(1 downto 0);
    signal VN1086_in4 : std_logic_vector(1 downto 0);
    signal VN1086_in5 : std_logic_vector(1 downto 0);
    signal VN1087_in0 : std_logic_vector(1 downto 0);
    signal VN1087_in1 : std_logic_vector(1 downto 0);
    signal VN1087_in2 : std_logic_vector(1 downto 0);
    signal VN1087_in3 : std_logic_vector(1 downto 0);
    signal VN1087_in4 : std_logic_vector(1 downto 0);
    signal VN1087_in5 : std_logic_vector(1 downto 0);
    signal VN1088_in0 : std_logic_vector(1 downto 0);
    signal VN1088_in1 : std_logic_vector(1 downto 0);
    signal VN1088_in2 : std_logic_vector(1 downto 0);
    signal VN1088_in3 : std_logic_vector(1 downto 0);
    signal VN1088_in4 : std_logic_vector(1 downto 0);
    signal VN1088_in5 : std_logic_vector(1 downto 0);
    signal VN1089_in0 : std_logic_vector(1 downto 0);
    signal VN1089_in1 : std_logic_vector(1 downto 0);
    signal VN1089_in2 : std_logic_vector(1 downto 0);
    signal VN1089_in3 : std_logic_vector(1 downto 0);
    signal VN1089_in4 : std_logic_vector(1 downto 0);
    signal VN1089_in5 : std_logic_vector(1 downto 0);
    signal VN1090_in0 : std_logic_vector(1 downto 0);
    signal VN1090_in1 : std_logic_vector(1 downto 0);
    signal VN1090_in2 : std_logic_vector(1 downto 0);
    signal VN1090_in3 : std_logic_vector(1 downto 0);
    signal VN1090_in4 : std_logic_vector(1 downto 0);
    signal VN1090_in5 : std_logic_vector(1 downto 0);
    signal VN1091_in0 : std_logic_vector(1 downto 0);
    signal VN1091_in1 : std_logic_vector(1 downto 0);
    signal VN1091_in2 : std_logic_vector(1 downto 0);
    signal VN1091_in3 : std_logic_vector(1 downto 0);
    signal VN1091_in4 : std_logic_vector(1 downto 0);
    signal VN1091_in5 : std_logic_vector(1 downto 0);
    signal VN1092_in0 : std_logic_vector(1 downto 0);
    signal VN1092_in1 : std_logic_vector(1 downto 0);
    signal VN1092_in2 : std_logic_vector(1 downto 0);
    signal VN1092_in3 : std_logic_vector(1 downto 0);
    signal VN1092_in4 : std_logic_vector(1 downto 0);
    signal VN1092_in5 : std_logic_vector(1 downto 0);
    signal VN1093_in0 : std_logic_vector(1 downto 0);
    signal VN1093_in1 : std_logic_vector(1 downto 0);
    signal VN1093_in2 : std_logic_vector(1 downto 0);
    signal VN1093_in3 : std_logic_vector(1 downto 0);
    signal VN1093_in4 : std_logic_vector(1 downto 0);
    signal VN1093_in5 : std_logic_vector(1 downto 0);
    signal VN1094_in0 : std_logic_vector(1 downto 0);
    signal VN1094_in1 : std_logic_vector(1 downto 0);
    signal VN1094_in2 : std_logic_vector(1 downto 0);
    signal VN1094_in3 : std_logic_vector(1 downto 0);
    signal VN1094_in4 : std_logic_vector(1 downto 0);
    signal VN1094_in5 : std_logic_vector(1 downto 0);
    signal VN1095_in0 : std_logic_vector(1 downto 0);
    signal VN1095_in1 : std_logic_vector(1 downto 0);
    signal VN1095_in2 : std_logic_vector(1 downto 0);
    signal VN1095_in3 : std_logic_vector(1 downto 0);
    signal VN1095_in4 : std_logic_vector(1 downto 0);
    signal VN1095_in5 : std_logic_vector(1 downto 0);
    signal VN1096_in0 : std_logic_vector(1 downto 0);
    signal VN1096_in1 : std_logic_vector(1 downto 0);
    signal VN1096_in2 : std_logic_vector(1 downto 0);
    signal VN1096_in3 : std_logic_vector(1 downto 0);
    signal VN1096_in4 : std_logic_vector(1 downto 0);
    signal VN1096_in5 : std_logic_vector(1 downto 0);
    signal VN1097_in0 : std_logic_vector(1 downto 0);
    signal VN1097_in1 : std_logic_vector(1 downto 0);
    signal VN1097_in2 : std_logic_vector(1 downto 0);
    signal VN1097_in3 : std_logic_vector(1 downto 0);
    signal VN1097_in4 : std_logic_vector(1 downto 0);
    signal VN1097_in5 : std_logic_vector(1 downto 0);
    signal VN1098_in0 : std_logic_vector(1 downto 0);
    signal VN1098_in1 : std_logic_vector(1 downto 0);
    signal VN1098_in2 : std_logic_vector(1 downto 0);
    signal VN1098_in3 : std_logic_vector(1 downto 0);
    signal VN1098_in4 : std_logic_vector(1 downto 0);
    signal VN1098_in5 : std_logic_vector(1 downto 0);
    signal VN1099_in0 : std_logic_vector(1 downto 0);
    signal VN1099_in1 : std_logic_vector(1 downto 0);
    signal VN1099_in2 : std_logic_vector(1 downto 0);
    signal VN1099_in3 : std_logic_vector(1 downto 0);
    signal VN1099_in4 : std_logic_vector(1 downto 0);
    signal VN1099_in5 : std_logic_vector(1 downto 0);
    signal VN1100_in0 : std_logic_vector(1 downto 0);
    signal VN1100_in1 : std_logic_vector(1 downto 0);
    signal VN1100_in2 : std_logic_vector(1 downto 0);
    signal VN1100_in3 : std_logic_vector(1 downto 0);
    signal VN1100_in4 : std_logic_vector(1 downto 0);
    signal VN1100_in5 : std_logic_vector(1 downto 0);
    signal VN1101_in0 : std_logic_vector(1 downto 0);
    signal VN1101_in1 : std_logic_vector(1 downto 0);
    signal VN1101_in2 : std_logic_vector(1 downto 0);
    signal VN1101_in3 : std_logic_vector(1 downto 0);
    signal VN1101_in4 : std_logic_vector(1 downto 0);
    signal VN1101_in5 : std_logic_vector(1 downto 0);
    signal VN1102_in0 : std_logic_vector(1 downto 0);
    signal VN1102_in1 : std_logic_vector(1 downto 0);
    signal VN1102_in2 : std_logic_vector(1 downto 0);
    signal VN1102_in3 : std_logic_vector(1 downto 0);
    signal VN1102_in4 : std_logic_vector(1 downto 0);
    signal VN1102_in5 : std_logic_vector(1 downto 0);
    signal VN1103_in0 : std_logic_vector(1 downto 0);
    signal VN1103_in1 : std_logic_vector(1 downto 0);
    signal VN1103_in2 : std_logic_vector(1 downto 0);
    signal VN1103_in3 : std_logic_vector(1 downto 0);
    signal VN1103_in4 : std_logic_vector(1 downto 0);
    signal VN1103_in5 : std_logic_vector(1 downto 0);
    signal VN1104_in0 : std_logic_vector(1 downto 0);
    signal VN1104_in1 : std_logic_vector(1 downto 0);
    signal VN1104_in2 : std_logic_vector(1 downto 0);
    signal VN1104_in3 : std_logic_vector(1 downto 0);
    signal VN1104_in4 : std_logic_vector(1 downto 0);
    signal VN1104_in5 : std_logic_vector(1 downto 0);
    signal VN1105_in0 : std_logic_vector(1 downto 0);
    signal VN1105_in1 : std_logic_vector(1 downto 0);
    signal VN1105_in2 : std_logic_vector(1 downto 0);
    signal VN1105_in3 : std_logic_vector(1 downto 0);
    signal VN1105_in4 : std_logic_vector(1 downto 0);
    signal VN1105_in5 : std_logic_vector(1 downto 0);
    signal VN1106_in0 : std_logic_vector(1 downto 0);
    signal VN1106_in1 : std_logic_vector(1 downto 0);
    signal VN1106_in2 : std_logic_vector(1 downto 0);
    signal VN1106_in3 : std_logic_vector(1 downto 0);
    signal VN1106_in4 : std_logic_vector(1 downto 0);
    signal VN1106_in5 : std_logic_vector(1 downto 0);
    signal VN1107_in0 : std_logic_vector(1 downto 0);
    signal VN1107_in1 : std_logic_vector(1 downto 0);
    signal VN1107_in2 : std_logic_vector(1 downto 0);
    signal VN1107_in3 : std_logic_vector(1 downto 0);
    signal VN1107_in4 : std_logic_vector(1 downto 0);
    signal VN1107_in5 : std_logic_vector(1 downto 0);
    signal VN1108_in0 : std_logic_vector(1 downto 0);
    signal VN1108_in1 : std_logic_vector(1 downto 0);
    signal VN1108_in2 : std_logic_vector(1 downto 0);
    signal VN1108_in3 : std_logic_vector(1 downto 0);
    signal VN1108_in4 : std_logic_vector(1 downto 0);
    signal VN1108_in5 : std_logic_vector(1 downto 0);
    signal VN1109_in0 : std_logic_vector(1 downto 0);
    signal VN1109_in1 : std_logic_vector(1 downto 0);
    signal VN1109_in2 : std_logic_vector(1 downto 0);
    signal VN1109_in3 : std_logic_vector(1 downto 0);
    signal VN1109_in4 : std_logic_vector(1 downto 0);
    signal VN1109_in5 : std_logic_vector(1 downto 0);
    signal VN1110_in0 : std_logic_vector(1 downto 0);
    signal VN1110_in1 : std_logic_vector(1 downto 0);
    signal VN1110_in2 : std_logic_vector(1 downto 0);
    signal VN1110_in3 : std_logic_vector(1 downto 0);
    signal VN1110_in4 : std_logic_vector(1 downto 0);
    signal VN1110_in5 : std_logic_vector(1 downto 0);
    signal VN1111_in0 : std_logic_vector(1 downto 0);
    signal VN1111_in1 : std_logic_vector(1 downto 0);
    signal VN1111_in2 : std_logic_vector(1 downto 0);
    signal VN1111_in3 : std_logic_vector(1 downto 0);
    signal VN1111_in4 : std_logic_vector(1 downto 0);
    signal VN1111_in5 : std_logic_vector(1 downto 0);
    signal VN1112_in0 : std_logic_vector(1 downto 0);
    signal VN1112_in1 : std_logic_vector(1 downto 0);
    signal VN1112_in2 : std_logic_vector(1 downto 0);
    signal VN1112_in3 : std_logic_vector(1 downto 0);
    signal VN1112_in4 : std_logic_vector(1 downto 0);
    signal VN1112_in5 : std_logic_vector(1 downto 0);
    signal VN1113_in0 : std_logic_vector(1 downto 0);
    signal VN1113_in1 : std_logic_vector(1 downto 0);
    signal VN1113_in2 : std_logic_vector(1 downto 0);
    signal VN1113_in3 : std_logic_vector(1 downto 0);
    signal VN1113_in4 : std_logic_vector(1 downto 0);
    signal VN1113_in5 : std_logic_vector(1 downto 0);
    signal VN1114_in0 : std_logic_vector(1 downto 0);
    signal VN1114_in1 : std_logic_vector(1 downto 0);
    signal VN1114_in2 : std_logic_vector(1 downto 0);
    signal VN1114_in3 : std_logic_vector(1 downto 0);
    signal VN1114_in4 : std_logic_vector(1 downto 0);
    signal VN1114_in5 : std_logic_vector(1 downto 0);
    signal VN1115_in0 : std_logic_vector(1 downto 0);
    signal VN1115_in1 : std_logic_vector(1 downto 0);
    signal VN1115_in2 : std_logic_vector(1 downto 0);
    signal VN1115_in3 : std_logic_vector(1 downto 0);
    signal VN1115_in4 : std_logic_vector(1 downto 0);
    signal VN1115_in5 : std_logic_vector(1 downto 0);
    signal VN1116_in0 : std_logic_vector(1 downto 0);
    signal VN1116_in1 : std_logic_vector(1 downto 0);
    signal VN1116_in2 : std_logic_vector(1 downto 0);
    signal VN1116_in3 : std_logic_vector(1 downto 0);
    signal VN1116_in4 : std_logic_vector(1 downto 0);
    signal VN1116_in5 : std_logic_vector(1 downto 0);
    signal VN1117_in0 : std_logic_vector(1 downto 0);
    signal VN1117_in1 : std_logic_vector(1 downto 0);
    signal VN1117_in2 : std_logic_vector(1 downto 0);
    signal VN1117_in3 : std_logic_vector(1 downto 0);
    signal VN1117_in4 : std_logic_vector(1 downto 0);
    signal VN1117_in5 : std_logic_vector(1 downto 0);
    signal VN1118_in0 : std_logic_vector(1 downto 0);
    signal VN1118_in1 : std_logic_vector(1 downto 0);
    signal VN1118_in2 : std_logic_vector(1 downto 0);
    signal VN1118_in3 : std_logic_vector(1 downto 0);
    signal VN1118_in4 : std_logic_vector(1 downto 0);
    signal VN1118_in5 : std_logic_vector(1 downto 0);
    signal VN1119_in0 : std_logic_vector(1 downto 0);
    signal VN1119_in1 : std_logic_vector(1 downto 0);
    signal VN1119_in2 : std_logic_vector(1 downto 0);
    signal VN1119_in3 : std_logic_vector(1 downto 0);
    signal VN1119_in4 : std_logic_vector(1 downto 0);
    signal VN1119_in5 : std_logic_vector(1 downto 0);
    signal VN1120_in0 : std_logic_vector(1 downto 0);
    signal VN1120_in1 : std_logic_vector(1 downto 0);
    signal VN1120_in2 : std_logic_vector(1 downto 0);
    signal VN1120_in3 : std_logic_vector(1 downto 0);
    signal VN1120_in4 : std_logic_vector(1 downto 0);
    signal VN1120_in5 : std_logic_vector(1 downto 0);
    signal VN1121_in0 : std_logic_vector(1 downto 0);
    signal VN1121_in1 : std_logic_vector(1 downto 0);
    signal VN1121_in2 : std_logic_vector(1 downto 0);
    signal VN1121_in3 : std_logic_vector(1 downto 0);
    signal VN1121_in4 : std_logic_vector(1 downto 0);
    signal VN1121_in5 : std_logic_vector(1 downto 0);
    signal VN1122_in0 : std_logic_vector(1 downto 0);
    signal VN1122_in1 : std_logic_vector(1 downto 0);
    signal VN1122_in2 : std_logic_vector(1 downto 0);
    signal VN1122_in3 : std_logic_vector(1 downto 0);
    signal VN1122_in4 : std_logic_vector(1 downto 0);
    signal VN1122_in5 : std_logic_vector(1 downto 0);
    signal VN1123_in0 : std_logic_vector(1 downto 0);
    signal VN1123_in1 : std_logic_vector(1 downto 0);
    signal VN1123_in2 : std_logic_vector(1 downto 0);
    signal VN1123_in3 : std_logic_vector(1 downto 0);
    signal VN1123_in4 : std_logic_vector(1 downto 0);
    signal VN1123_in5 : std_logic_vector(1 downto 0);
    signal VN1124_in0 : std_logic_vector(1 downto 0);
    signal VN1124_in1 : std_logic_vector(1 downto 0);
    signal VN1124_in2 : std_logic_vector(1 downto 0);
    signal VN1124_in3 : std_logic_vector(1 downto 0);
    signal VN1124_in4 : std_logic_vector(1 downto 0);
    signal VN1124_in5 : std_logic_vector(1 downto 0);
    signal VN1125_in0 : std_logic_vector(1 downto 0);
    signal VN1125_in1 : std_logic_vector(1 downto 0);
    signal VN1125_in2 : std_logic_vector(1 downto 0);
    signal VN1125_in3 : std_logic_vector(1 downto 0);
    signal VN1125_in4 : std_logic_vector(1 downto 0);
    signal VN1125_in5 : std_logic_vector(1 downto 0);
    signal VN1126_in0 : std_logic_vector(1 downto 0);
    signal VN1126_in1 : std_logic_vector(1 downto 0);
    signal VN1126_in2 : std_logic_vector(1 downto 0);
    signal VN1126_in3 : std_logic_vector(1 downto 0);
    signal VN1126_in4 : std_logic_vector(1 downto 0);
    signal VN1126_in5 : std_logic_vector(1 downto 0);
    signal VN1127_in0 : std_logic_vector(1 downto 0);
    signal VN1127_in1 : std_logic_vector(1 downto 0);
    signal VN1127_in2 : std_logic_vector(1 downto 0);
    signal VN1127_in3 : std_logic_vector(1 downto 0);
    signal VN1127_in4 : std_logic_vector(1 downto 0);
    signal VN1127_in5 : std_logic_vector(1 downto 0);
    signal VN1128_in0 : std_logic_vector(1 downto 0);
    signal VN1128_in1 : std_logic_vector(1 downto 0);
    signal VN1128_in2 : std_logic_vector(1 downto 0);
    signal VN1128_in3 : std_logic_vector(1 downto 0);
    signal VN1128_in4 : std_logic_vector(1 downto 0);
    signal VN1128_in5 : std_logic_vector(1 downto 0);
    signal VN1129_in0 : std_logic_vector(1 downto 0);
    signal VN1129_in1 : std_logic_vector(1 downto 0);
    signal VN1129_in2 : std_logic_vector(1 downto 0);
    signal VN1129_in3 : std_logic_vector(1 downto 0);
    signal VN1129_in4 : std_logic_vector(1 downto 0);
    signal VN1129_in5 : std_logic_vector(1 downto 0);
    signal VN1130_in0 : std_logic_vector(1 downto 0);
    signal VN1130_in1 : std_logic_vector(1 downto 0);
    signal VN1130_in2 : std_logic_vector(1 downto 0);
    signal VN1130_in3 : std_logic_vector(1 downto 0);
    signal VN1130_in4 : std_logic_vector(1 downto 0);
    signal VN1130_in5 : std_logic_vector(1 downto 0);
    signal VN1131_in0 : std_logic_vector(1 downto 0);
    signal VN1131_in1 : std_logic_vector(1 downto 0);
    signal VN1131_in2 : std_logic_vector(1 downto 0);
    signal VN1131_in3 : std_logic_vector(1 downto 0);
    signal VN1131_in4 : std_logic_vector(1 downto 0);
    signal VN1131_in5 : std_logic_vector(1 downto 0);
    signal VN1132_in0 : std_logic_vector(1 downto 0);
    signal VN1132_in1 : std_logic_vector(1 downto 0);
    signal VN1132_in2 : std_logic_vector(1 downto 0);
    signal VN1132_in3 : std_logic_vector(1 downto 0);
    signal VN1132_in4 : std_logic_vector(1 downto 0);
    signal VN1132_in5 : std_logic_vector(1 downto 0);
    signal VN1133_in0 : std_logic_vector(1 downto 0);
    signal VN1133_in1 : std_logic_vector(1 downto 0);
    signal VN1133_in2 : std_logic_vector(1 downto 0);
    signal VN1133_in3 : std_logic_vector(1 downto 0);
    signal VN1133_in4 : std_logic_vector(1 downto 0);
    signal VN1133_in5 : std_logic_vector(1 downto 0);
    signal VN1134_in0 : std_logic_vector(1 downto 0);
    signal VN1134_in1 : std_logic_vector(1 downto 0);
    signal VN1134_in2 : std_logic_vector(1 downto 0);
    signal VN1134_in3 : std_logic_vector(1 downto 0);
    signal VN1134_in4 : std_logic_vector(1 downto 0);
    signal VN1134_in5 : std_logic_vector(1 downto 0);
    signal VN1135_in0 : std_logic_vector(1 downto 0);
    signal VN1135_in1 : std_logic_vector(1 downto 0);
    signal VN1135_in2 : std_logic_vector(1 downto 0);
    signal VN1135_in3 : std_logic_vector(1 downto 0);
    signal VN1135_in4 : std_logic_vector(1 downto 0);
    signal VN1135_in5 : std_logic_vector(1 downto 0);
    signal VN1136_in0 : std_logic_vector(1 downto 0);
    signal VN1136_in1 : std_logic_vector(1 downto 0);
    signal VN1136_in2 : std_logic_vector(1 downto 0);
    signal VN1136_in3 : std_logic_vector(1 downto 0);
    signal VN1136_in4 : std_logic_vector(1 downto 0);
    signal VN1136_in5 : std_logic_vector(1 downto 0);
    signal VN1137_in0 : std_logic_vector(1 downto 0);
    signal VN1137_in1 : std_logic_vector(1 downto 0);
    signal VN1137_in2 : std_logic_vector(1 downto 0);
    signal VN1137_in3 : std_logic_vector(1 downto 0);
    signal VN1137_in4 : std_logic_vector(1 downto 0);
    signal VN1137_in5 : std_logic_vector(1 downto 0);
    signal VN1138_in0 : std_logic_vector(1 downto 0);
    signal VN1138_in1 : std_logic_vector(1 downto 0);
    signal VN1138_in2 : std_logic_vector(1 downto 0);
    signal VN1138_in3 : std_logic_vector(1 downto 0);
    signal VN1138_in4 : std_logic_vector(1 downto 0);
    signal VN1138_in5 : std_logic_vector(1 downto 0);
    signal VN1139_in0 : std_logic_vector(1 downto 0);
    signal VN1139_in1 : std_logic_vector(1 downto 0);
    signal VN1139_in2 : std_logic_vector(1 downto 0);
    signal VN1139_in3 : std_logic_vector(1 downto 0);
    signal VN1139_in4 : std_logic_vector(1 downto 0);
    signal VN1139_in5 : std_logic_vector(1 downto 0);
    signal VN1140_in0 : std_logic_vector(1 downto 0);
    signal VN1140_in1 : std_logic_vector(1 downto 0);
    signal VN1140_in2 : std_logic_vector(1 downto 0);
    signal VN1140_in3 : std_logic_vector(1 downto 0);
    signal VN1140_in4 : std_logic_vector(1 downto 0);
    signal VN1140_in5 : std_logic_vector(1 downto 0);
    signal VN1141_in0 : std_logic_vector(1 downto 0);
    signal VN1141_in1 : std_logic_vector(1 downto 0);
    signal VN1141_in2 : std_logic_vector(1 downto 0);
    signal VN1141_in3 : std_logic_vector(1 downto 0);
    signal VN1141_in4 : std_logic_vector(1 downto 0);
    signal VN1141_in5 : std_logic_vector(1 downto 0);
    signal VN1142_in0 : std_logic_vector(1 downto 0);
    signal VN1142_in1 : std_logic_vector(1 downto 0);
    signal VN1142_in2 : std_logic_vector(1 downto 0);
    signal VN1142_in3 : std_logic_vector(1 downto 0);
    signal VN1142_in4 : std_logic_vector(1 downto 0);
    signal VN1142_in5 : std_logic_vector(1 downto 0);
    signal VN1143_in0 : std_logic_vector(1 downto 0);
    signal VN1143_in1 : std_logic_vector(1 downto 0);
    signal VN1143_in2 : std_logic_vector(1 downto 0);
    signal VN1143_in3 : std_logic_vector(1 downto 0);
    signal VN1143_in4 : std_logic_vector(1 downto 0);
    signal VN1143_in5 : std_logic_vector(1 downto 0);
    signal VN1144_in0 : std_logic_vector(1 downto 0);
    signal VN1144_in1 : std_logic_vector(1 downto 0);
    signal VN1144_in2 : std_logic_vector(1 downto 0);
    signal VN1144_in3 : std_logic_vector(1 downto 0);
    signal VN1144_in4 : std_logic_vector(1 downto 0);
    signal VN1144_in5 : std_logic_vector(1 downto 0);
    signal VN1145_in0 : std_logic_vector(1 downto 0);
    signal VN1145_in1 : std_logic_vector(1 downto 0);
    signal VN1145_in2 : std_logic_vector(1 downto 0);
    signal VN1145_in3 : std_logic_vector(1 downto 0);
    signal VN1145_in4 : std_logic_vector(1 downto 0);
    signal VN1145_in5 : std_logic_vector(1 downto 0);
    signal VN1146_in0 : std_logic_vector(1 downto 0);
    signal VN1146_in1 : std_logic_vector(1 downto 0);
    signal VN1146_in2 : std_logic_vector(1 downto 0);
    signal VN1146_in3 : std_logic_vector(1 downto 0);
    signal VN1146_in4 : std_logic_vector(1 downto 0);
    signal VN1146_in5 : std_logic_vector(1 downto 0);
    signal VN1147_in0 : std_logic_vector(1 downto 0);
    signal VN1147_in1 : std_logic_vector(1 downto 0);
    signal VN1147_in2 : std_logic_vector(1 downto 0);
    signal VN1147_in3 : std_logic_vector(1 downto 0);
    signal VN1147_in4 : std_logic_vector(1 downto 0);
    signal VN1147_in5 : std_logic_vector(1 downto 0);
    signal VN1148_in0 : std_logic_vector(1 downto 0);
    signal VN1148_in1 : std_logic_vector(1 downto 0);
    signal VN1148_in2 : std_logic_vector(1 downto 0);
    signal VN1148_in3 : std_logic_vector(1 downto 0);
    signal VN1148_in4 : std_logic_vector(1 downto 0);
    signal VN1148_in5 : std_logic_vector(1 downto 0);
    signal VN1149_in0 : std_logic_vector(1 downto 0);
    signal VN1149_in1 : std_logic_vector(1 downto 0);
    signal VN1149_in2 : std_logic_vector(1 downto 0);
    signal VN1149_in3 : std_logic_vector(1 downto 0);
    signal VN1149_in4 : std_logic_vector(1 downto 0);
    signal VN1149_in5 : std_logic_vector(1 downto 0);
    signal VN1150_in0 : std_logic_vector(1 downto 0);
    signal VN1150_in1 : std_logic_vector(1 downto 0);
    signal VN1150_in2 : std_logic_vector(1 downto 0);
    signal VN1150_in3 : std_logic_vector(1 downto 0);
    signal VN1150_in4 : std_logic_vector(1 downto 0);
    signal VN1150_in5 : std_logic_vector(1 downto 0);
    signal VN1151_in0 : std_logic_vector(1 downto 0);
    signal VN1151_in1 : std_logic_vector(1 downto 0);
    signal VN1151_in2 : std_logic_vector(1 downto 0);
    signal VN1151_in3 : std_logic_vector(1 downto 0);
    signal VN1151_in4 : std_logic_vector(1 downto 0);
    signal VN1151_in5 : std_logic_vector(1 downto 0);
    signal VN1152_in0 : std_logic_vector(1 downto 0);
    signal VN1152_in1 : std_logic_vector(1 downto 0);
    signal VN1152_in2 : std_logic_vector(1 downto 0);
    signal VN1152_in3 : std_logic_vector(1 downto 0);
    signal VN1152_in4 : std_logic_vector(1 downto 0);
    signal VN1152_in5 : std_logic_vector(1 downto 0);
    signal VN1153_in0 : std_logic_vector(1 downto 0);
    signal VN1153_in1 : std_logic_vector(1 downto 0);
    signal VN1153_in2 : std_logic_vector(1 downto 0);
    signal VN1153_in3 : std_logic_vector(1 downto 0);
    signal VN1153_in4 : std_logic_vector(1 downto 0);
    signal VN1153_in5 : std_logic_vector(1 downto 0);
    signal VN1154_in0 : std_logic_vector(1 downto 0);
    signal VN1154_in1 : std_logic_vector(1 downto 0);
    signal VN1154_in2 : std_logic_vector(1 downto 0);
    signal VN1154_in3 : std_logic_vector(1 downto 0);
    signal VN1154_in4 : std_logic_vector(1 downto 0);
    signal VN1154_in5 : std_logic_vector(1 downto 0);
    signal VN1155_in0 : std_logic_vector(1 downto 0);
    signal VN1155_in1 : std_logic_vector(1 downto 0);
    signal VN1155_in2 : std_logic_vector(1 downto 0);
    signal VN1155_in3 : std_logic_vector(1 downto 0);
    signal VN1155_in4 : std_logic_vector(1 downto 0);
    signal VN1155_in5 : std_logic_vector(1 downto 0);
    signal VN1156_in0 : std_logic_vector(1 downto 0);
    signal VN1156_in1 : std_logic_vector(1 downto 0);
    signal VN1156_in2 : std_logic_vector(1 downto 0);
    signal VN1156_in3 : std_logic_vector(1 downto 0);
    signal VN1156_in4 : std_logic_vector(1 downto 0);
    signal VN1156_in5 : std_logic_vector(1 downto 0);
    signal VN1157_in0 : std_logic_vector(1 downto 0);
    signal VN1157_in1 : std_logic_vector(1 downto 0);
    signal VN1157_in2 : std_logic_vector(1 downto 0);
    signal VN1157_in3 : std_logic_vector(1 downto 0);
    signal VN1157_in4 : std_logic_vector(1 downto 0);
    signal VN1157_in5 : std_logic_vector(1 downto 0);
    signal VN1158_in0 : std_logic_vector(1 downto 0);
    signal VN1158_in1 : std_logic_vector(1 downto 0);
    signal VN1158_in2 : std_logic_vector(1 downto 0);
    signal VN1158_in3 : std_logic_vector(1 downto 0);
    signal VN1158_in4 : std_logic_vector(1 downto 0);
    signal VN1158_in5 : std_logic_vector(1 downto 0);
    signal VN1159_in0 : std_logic_vector(1 downto 0);
    signal VN1159_in1 : std_logic_vector(1 downto 0);
    signal VN1159_in2 : std_logic_vector(1 downto 0);
    signal VN1159_in3 : std_logic_vector(1 downto 0);
    signal VN1159_in4 : std_logic_vector(1 downto 0);
    signal VN1159_in5 : std_logic_vector(1 downto 0);
    signal VN1160_in0 : std_logic_vector(1 downto 0);
    signal VN1160_in1 : std_logic_vector(1 downto 0);
    signal VN1160_in2 : std_logic_vector(1 downto 0);
    signal VN1160_in3 : std_logic_vector(1 downto 0);
    signal VN1160_in4 : std_logic_vector(1 downto 0);
    signal VN1160_in5 : std_logic_vector(1 downto 0);
    signal VN1161_in0 : std_logic_vector(1 downto 0);
    signal VN1161_in1 : std_logic_vector(1 downto 0);
    signal VN1161_in2 : std_logic_vector(1 downto 0);
    signal VN1161_in3 : std_logic_vector(1 downto 0);
    signal VN1161_in4 : std_logic_vector(1 downto 0);
    signal VN1161_in5 : std_logic_vector(1 downto 0);
    signal VN1162_in0 : std_logic_vector(1 downto 0);
    signal VN1162_in1 : std_logic_vector(1 downto 0);
    signal VN1162_in2 : std_logic_vector(1 downto 0);
    signal VN1162_in3 : std_logic_vector(1 downto 0);
    signal VN1162_in4 : std_logic_vector(1 downto 0);
    signal VN1162_in5 : std_logic_vector(1 downto 0);
    signal VN1163_in0 : std_logic_vector(1 downto 0);
    signal VN1163_in1 : std_logic_vector(1 downto 0);
    signal VN1163_in2 : std_logic_vector(1 downto 0);
    signal VN1163_in3 : std_logic_vector(1 downto 0);
    signal VN1163_in4 : std_logic_vector(1 downto 0);
    signal VN1163_in5 : std_logic_vector(1 downto 0);
    signal VN1164_in0 : std_logic_vector(1 downto 0);
    signal VN1164_in1 : std_logic_vector(1 downto 0);
    signal VN1164_in2 : std_logic_vector(1 downto 0);
    signal VN1164_in3 : std_logic_vector(1 downto 0);
    signal VN1164_in4 : std_logic_vector(1 downto 0);
    signal VN1164_in5 : std_logic_vector(1 downto 0);
    signal VN1165_in0 : std_logic_vector(1 downto 0);
    signal VN1165_in1 : std_logic_vector(1 downto 0);
    signal VN1165_in2 : std_logic_vector(1 downto 0);
    signal VN1165_in3 : std_logic_vector(1 downto 0);
    signal VN1165_in4 : std_logic_vector(1 downto 0);
    signal VN1165_in5 : std_logic_vector(1 downto 0);
    signal VN1166_in0 : std_logic_vector(1 downto 0);
    signal VN1166_in1 : std_logic_vector(1 downto 0);
    signal VN1166_in2 : std_logic_vector(1 downto 0);
    signal VN1166_in3 : std_logic_vector(1 downto 0);
    signal VN1166_in4 : std_logic_vector(1 downto 0);
    signal VN1166_in5 : std_logic_vector(1 downto 0);
    signal VN1167_in0 : std_logic_vector(1 downto 0);
    signal VN1167_in1 : std_logic_vector(1 downto 0);
    signal VN1167_in2 : std_logic_vector(1 downto 0);
    signal VN1167_in3 : std_logic_vector(1 downto 0);
    signal VN1167_in4 : std_logic_vector(1 downto 0);
    signal VN1167_in5 : std_logic_vector(1 downto 0);
    signal VN1168_in0 : std_logic_vector(1 downto 0);
    signal VN1168_in1 : std_logic_vector(1 downto 0);
    signal VN1168_in2 : std_logic_vector(1 downto 0);
    signal VN1168_in3 : std_logic_vector(1 downto 0);
    signal VN1168_in4 : std_logic_vector(1 downto 0);
    signal VN1168_in5 : std_logic_vector(1 downto 0);
    signal VN1169_in0 : std_logic_vector(1 downto 0);
    signal VN1169_in1 : std_logic_vector(1 downto 0);
    signal VN1169_in2 : std_logic_vector(1 downto 0);
    signal VN1169_in3 : std_logic_vector(1 downto 0);
    signal VN1169_in4 : std_logic_vector(1 downto 0);
    signal VN1169_in5 : std_logic_vector(1 downto 0);
    signal VN1170_in0 : std_logic_vector(1 downto 0);
    signal VN1170_in1 : std_logic_vector(1 downto 0);
    signal VN1170_in2 : std_logic_vector(1 downto 0);
    signal VN1170_in3 : std_logic_vector(1 downto 0);
    signal VN1170_in4 : std_logic_vector(1 downto 0);
    signal VN1170_in5 : std_logic_vector(1 downto 0);
    signal VN1171_in0 : std_logic_vector(1 downto 0);
    signal VN1171_in1 : std_logic_vector(1 downto 0);
    signal VN1171_in2 : std_logic_vector(1 downto 0);
    signal VN1171_in3 : std_logic_vector(1 downto 0);
    signal VN1171_in4 : std_logic_vector(1 downto 0);
    signal VN1171_in5 : std_logic_vector(1 downto 0);
    signal VN1172_in0 : std_logic_vector(1 downto 0);
    signal VN1172_in1 : std_logic_vector(1 downto 0);
    signal VN1172_in2 : std_logic_vector(1 downto 0);
    signal VN1172_in3 : std_logic_vector(1 downto 0);
    signal VN1172_in4 : std_logic_vector(1 downto 0);
    signal VN1172_in5 : std_logic_vector(1 downto 0);
    signal VN1173_in0 : std_logic_vector(1 downto 0);
    signal VN1173_in1 : std_logic_vector(1 downto 0);
    signal VN1173_in2 : std_logic_vector(1 downto 0);
    signal VN1173_in3 : std_logic_vector(1 downto 0);
    signal VN1173_in4 : std_logic_vector(1 downto 0);
    signal VN1173_in5 : std_logic_vector(1 downto 0);
    signal VN1174_in0 : std_logic_vector(1 downto 0);
    signal VN1174_in1 : std_logic_vector(1 downto 0);
    signal VN1174_in2 : std_logic_vector(1 downto 0);
    signal VN1174_in3 : std_logic_vector(1 downto 0);
    signal VN1174_in4 : std_logic_vector(1 downto 0);
    signal VN1174_in5 : std_logic_vector(1 downto 0);
    signal VN1175_in0 : std_logic_vector(1 downto 0);
    signal VN1175_in1 : std_logic_vector(1 downto 0);
    signal VN1175_in2 : std_logic_vector(1 downto 0);
    signal VN1175_in3 : std_logic_vector(1 downto 0);
    signal VN1175_in4 : std_logic_vector(1 downto 0);
    signal VN1175_in5 : std_logic_vector(1 downto 0);
    signal VN1176_in0 : std_logic_vector(1 downto 0);
    signal VN1176_in1 : std_logic_vector(1 downto 0);
    signal VN1176_in2 : std_logic_vector(1 downto 0);
    signal VN1176_in3 : std_logic_vector(1 downto 0);
    signal VN1176_in4 : std_logic_vector(1 downto 0);
    signal VN1176_in5 : std_logic_vector(1 downto 0);
    signal VN1177_in0 : std_logic_vector(1 downto 0);
    signal VN1177_in1 : std_logic_vector(1 downto 0);
    signal VN1177_in2 : std_logic_vector(1 downto 0);
    signal VN1177_in3 : std_logic_vector(1 downto 0);
    signal VN1177_in4 : std_logic_vector(1 downto 0);
    signal VN1177_in5 : std_logic_vector(1 downto 0);
    signal VN1178_in0 : std_logic_vector(1 downto 0);
    signal VN1178_in1 : std_logic_vector(1 downto 0);
    signal VN1178_in2 : std_logic_vector(1 downto 0);
    signal VN1178_in3 : std_logic_vector(1 downto 0);
    signal VN1178_in4 : std_logic_vector(1 downto 0);
    signal VN1178_in5 : std_logic_vector(1 downto 0);
    signal VN1179_in0 : std_logic_vector(1 downto 0);
    signal VN1179_in1 : std_logic_vector(1 downto 0);
    signal VN1179_in2 : std_logic_vector(1 downto 0);
    signal VN1179_in3 : std_logic_vector(1 downto 0);
    signal VN1179_in4 : std_logic_vector(1 downto 0);
    signal VN1179_in5 : std_logic_vector(1 downto 0);
    signal VN1180_in0 : std_logic_vector(1 downto 0);
    signal VN1180_in1 : std_logic_vector(1 downto 0);
    signal VN1180_in2 : std_logic_vector(1 downto 0);
    signal VN1180_in3 : std_logic_vector(1 downto 0);
    signal VN1180_in4 : std_logic_vector(1 downto 0);
    signal VN1180_in5 : std_logic_vector(1 downto 0);
    signal VN1181_in0 : std_logic_vector(1 downto 0);
    signal VN1181_in1 : std_logic_vector(1 downto 0);
    signal VN1181_in2 : std_logic_vector(1 downto 0);
    signal VN1181_in3 : std_logic_vector(1 downto 0);
    signal VN1181_in4 : std_logic_vector(1 downto 0);
    signal VN1181_in5 : std_logic_vector(1 downto 0);
    signal VN1182_in0 : std_logic_vector(1 downto 0);
    signal VN1182_in1 : std_logic_vector(1 downto 0);
    signal VN1182_in2 : std_logic_vector(1 downto 0);
    signal VN1182_in3 : std_logic_vector(1 downto 0);
    signal VN1182_in4 : std_logic_vector(1 downto 0);
    signal VN1182_in5 : std_logic_vector(1 downto 0);
    signal VN1183_in0 : std_logic_vector(1 downto 0);
    signal VN1183_in1 : std_logic_vector(1 downto 0);
    signal VN1183_in2 : std_logic_vector(1 downto 0);
    signal VN1183_in3 : std_logic_vector(1 downto 0);
    signal VN1183_in4 : std_logic_vector(1 downto 0);
    signal VN1183_in5 : std_logic_vector(1 downto 0);
    signal VN1184_in0 : std_logic_vector(1 downto 0);
    signal VN1184_in1 : std_logic_vector(1 downto 0);
    signal VN1184_in2 : std_logic_vector(1 downto 0);
    signal VN1184_in3 : std_logic_vector(1 downto 0);
    signal VN1184_in4 : std_logic_vector(1 downto 0);
    signal VN1184_in5 : std_logic_vector(1 downto 0);
    signal VN1185_in0 : std_logic_vector(1 downto 0);
    signal VN1185_in1 : std_logic_vector(1 downto 0);
    signal VN1185_in2 : std_logic_vector(1 downto 0);
    signal VN1185_in3 : std_logic_vector(1 downto 0);
    signal VN1185_in4 : std_logic_vector(1 downto 0);
    signal VN1185_in5 : std_logic_vector(1 downto 0);
    signal VN1186_in0 : std_logic_vector(1 downto 0);
    signal VN1186_in1 : std_logic_vector(1 downto 0);
    signal VN1186_in2 : std_logic_vector(1 downto 0);
    signal VN1186_in3 : std_logic_vector(1 downto 0);
    signal VN1186_in4 : std_logic_vector(1 downto 0);
    signal VN1186_in5 : std_logic_vector(1 downto 0);
    signal VN1187_in0 : std_logic_vector(1 downto 0);
    signal VN1187_in1 : std_logic_vector(1 downto 0);
    signal VN1187_in2 : std_logic_vector(1 downto 0);
    signal VN1187_in3 : std_logic_vector(1 downto 0);
    signal VN1187_in4 : std_logic_vector(1 downto 0);
    signal VN1187_in5 : std_logic_vector(1 downto 0);
    signal VN1188_in0 : std_logic_vector(1 downto 0);
    signal VN1188_in1 : std_logic_vector(1 downto 0);
    signal VN1188_in2 : std_logic_vector(1 downto 0);
    signal VN1188_in3 : std_logic_vector(1 downto 0);
    signal VN1188_in4 : std_logic_vector(1 downto 0);
    signal VN1188_in5 : std_logic_vector(1 downto 0);
    signal VN1189_in0 : std_logic_vector(1 downto 0);
    signal VN1189_in1 : std_logic_vector(1 downto 0);
    signal VN1189_in2 : std_logic_vector(1 downto 0);
    signal VN1189_in3 : std_logic_vector(1 downto 0);
    signal VN1189_in4 : std_logic_vector(1 downto 0);
    signal VN1189_in5 : std_logic_vector(1 downto 0);
    signal VN1190_in0 : std_logic_vector(1 downto 0);
    signal VN1190_in1 : std_logic_vector(1 downto 0);
    signal VN1190_in2 : std_logic_vector(1 downto 0);
    signal VN1190_in3 : std_logic_vector(1 downto 0);
    signal VN1190_in4 : std_logic_vector(1 downto 0);
    signal VN1190_in5 : std_logic_vector(1 downto 0);
    signal VN1191_in0 : std_logic_vector(1 downto 0);
    signal VN1191_in1 : std_logic_vector(1 downto 0);
    signal VN1191_in2 : std_logic_vector(1 downto 0);
    signal VN1191_in3 : std_logic_vector(1 downto 0);
    signal VN1191_in4 : std_logic_vector(1 downto 0);
    signal VN1191_in5 : std_logic_vector(1 downto 0);
    signal VN1192_in0 : std_logic_vector(1 downto 0);
    signal VN1192_in1 : std_logic_vector(1 downto 0);
    signal VN1192_in2 : std_logic_vector(1 downto 0);
    signal VN1192_in3 : std_logic_vector(1 downto 0);
    signal VN1192_in4 : std_logic_vector(1 downto 0);
    signal VN1192_in5 : std_logic_vector(1 downto 0);
    signal VN1193_in0 : std_logic_vector(1 downto 0);
    signal VN1193_in1 : std_logic_vector(1 downto 0);
    signal VN1193_in2 : std_logic_vector(1 downto 0);
    signal VN1193_in3 : std_logic_vector(1 downto 0);
    signal VN1193_in4 : std_logic_vector(1 downto 0);
    signal VN1193_in5 : std_logic_vector(1 downto 0);
    signal VN1194_in0 : std_logic_vector(1 downto 0);
    signal VN1194_in1 : std_logic_vector(1 downto 0);
    signal VN1194_in2 : std_logic_vector(1 downto 0);
    signal VN1194_in3 : std_logic_vector(1 downto 0);
    signal VN1194_in4 : std_logic_vector(1 downto 0);
    signal VN1194_in5 : std_logic_vector(1 downto 0);
    signal VN1195_in0 : std_logic_vector(1 downto 0);
    signal VN1195_in1 : std_logic_vector(1 downto 0);
    signal VN1195_in2 : std_logic_vector(1 downto 0);
    signal VN1195_in3 : std_logic_vector(1 downto 0);
    signal VN1195_in4 : std_logic_vector(1 downto 0);
    signal VN1195_in5 : std_logic_vector(1 downto 0);
    signal VN1196_in0 : std_logic_vector(1 downto 0);
    signal VN1196_in1 : std_logic_vector(1 downto 0);
    signal VN1196_in2 : std_logic_vector(1 downto 0);
    signal VN1196_in3 : std_logic_vector(1 downto 0);
    signal VN1196_in4 : std_logic_vector(1 downto 0);
    signal VN1196_in5 : std_logic_vector(1 downto 0);
    signal VN1197_in0 : std_logic_vector(1 downto 0);
    signal VN1197_in1 : std_logic_vector(1 downto 0);
    signal VN1197_in2 : std_logic_vector(1 downto 0);
    signal VN1197_in3 : std_logic_vector(1 downto 0);
    signal VN1197_in4 : std_logic_vector(1 downto 0);
    signal VN1197_in5 : std_logic_vector(1 downto 0);
    signal VN1198_in0 : std_logic_vector(1 downto 0);
    signal VN1198_in1 : std_logic_vector(1 downto 0);
    signal VN1198_in2 : std_logic_vector(1 downto 0);
    signal VN1198_in3 : std_logic_vector(1 downto 0);
    signal VN1198_in4 : std_logic_vector(1 downto 0);
    signal VN1198_in5 : std_logic_vector(1 downto 0);
    signal VN1199_in0 : std_logic_vector(1 downto 0);
    signal VN1199_in1 : std_logic_vector(1 downto 0);
    signal VN1199_in2 : std_logic_vector(1 downto 0);
    signal VN1199_in3 : std_logic_vector(1 downto 0);
    signal VN1199_in4 : std_logic_vector(1 downto 0);
    signal VN1199_in5 : std_logic_vector(1 downto 0);
    signal VN1200_in0 : std_logic_vector(1 downto 0);
    signal VN1200_in1 : std_logic_vector(1 downto 0);
    signal VN1200_in2 : std_logic_vector(1 downto 0);
    signal VN1200_in3 : std_logic_vector(1 downto 0);
    signal VN1200_in4 : std_logic_vector(1 downto 0);
    signal VN1200_in5 : std_logic_vector(1 downto 0);
    signal VN1201_in0 : std_logic_vector(1 downto 0);
    signal VN1201_in1 : std_logic_vector(1 downto 0);
    signal VN1201_in2 : std_logic_vector(1 downto 0);
    signal VN1201_in3 : std_logic_vector(1 downto 0);
    signal VN1201_in4 : std_logic_vector(1 downto 0);
    signal VN1201_in5 : std_logic_vector(1 downto 0);
    signal VN1202_in0 : std_logic_vector(1 downto 0);
    signal VN1202_in1 : std_logic_vector(1 downto 0);
    signal VN1202_in2 : std_logic_vector(1 downto 0);
    signal VN1202_in3 : std_logic_vector(1 downto 0);
    signal VN1202_in4 : std_logic_vector(1 downto 0);
    signal VN1202_in5 : std_logic_vector(1 downto 0);
    signal VN1203_in0 : std_logic_vector(1 downto 0);
    signal VN1203_in1 : std_logic_vector(1 downto 0);
    signal VN1203_in2 : std_logic_vector(1 downto 0);
    signal VN1203_in3 : std_logic_vector(1 downto 0);
    signal VN1203_in4 : std_logic_vector(1 downto 0);
    signal VN1203_in5 : std_logic_vector(1 downto 0);
    signal VN1204_in0 : std_logic_vector(1 downto 0);
    signal VN1204_in1 : std_logic_vector(1 downto 0);
    signal VN1204_in2 : std_logic_vector(1 downto 0);
    signal VN1204_in3 : std_logic_vector(1 downto 0);
    signal VN1204_in4 : std_logic_vector(1 downto 0);
    signal VN1204_in5 : std_logic_vector(1 downto 0);
    signal VN1205_in0 : std_logic_vector(1 downto 0);
    signal VN1205_in1 : std_logic_vector(1 downto 0);
    signal VN1205_in2 : std_logic_vector(1 downto 0);
    signal VN1205_in3 : std_logic_vector(1 downto 0);
    signal VN1205_in4 : std_logic_vector(1 downto 0);
    signal VN1205_in5 : std_logic_vector(1 downto 0);
    signal VN1206_in0 : std_logic_vector(1 downto 0);
    signal VN1206_in1 : std_logic_vector(1 downto 0);
    signal VN1206_in2 : std_logic_vector(1 downto 0);
    signal VN1206_in3 : std_logic_vector(1 downto 0);
    signal VN1206_in4 : std_logic_vector(1 downto 0);
    signal VN1206_in5 : std_logic_vector(1 downto 0);
    signal VN1207_in0 : std_logic_vector(1 downto 0);
    signal VN1207_in1 : std_logic_vector(1 downto 0);
    signal VN1207_in2 : std_logic_vector(1 downto 0);
    signal VN1207_in3 : std_logic_vector(1 downto 0);
    signal VN1207_in4 : std_logic_vector(1 downto 0);
    signal VN1207_in5 : std_logic_vector(1 downto 0);
    signal VN1208_in0 : std_logic_vector(1 downto 0);
    signal VN1208_in1 : std_logic_vector(1 downto 0);
    signal VN1208_in2 : std_logic_vector(1 downto 0);
    signal VN1208_in3 : std_logic_vector(1 downto 0);
    signal VN1208_in4 : std_logic_vector(1 downto 0);
    signal VN1208_in5 : std_logic_vector(1 downto 0);
    signal VN1209_in0 : std_logic_vector(1 downto 0);
    signal VN1209_in1 : std_logic_vector(1 downto 0);
    signal VN1209_in2 : std_logic_vector(1 downto 0);
    signal VN1209_in3 : std_logic_vector(1 downto 0);
    signal VN1209_in4 : std_logic_vector(1 downto 0);
    signal VN1209_in5 : std_logic_vector(1 downto 0);
    signal VN1210_in0 : std_logic_vector(1 downto 0);
    signal VN1210_in1 : std_logic_vector(1 downto 0);
    signal VN1210_in2 : std_logic_vector(1 downto 0);
    signal VN1210_in3 : std_logic_vector(1 downto 0);
    signal VN1210_in4 : std_logic_vector(1 downto 0);
    signal VN1210_in5 : std_logic_vector(1 downto 0);
    signal VN1211_in0 : std_logic_vector(1 downto 0);
    signal VN1211_in1 : std_logic_vector(1 downto 0);
    signal VN1211_in2 : std_logic_vector(1 downto 0);
    signal VN1211_in3 : std_logic_vector(1 downto 0);
    signal VN1211_in4 : std_logic_vector(1 downto 0);
    signal VN1211_in5 : std_logic_vector(1 downto 0);
    signal VN1212_in0 : std_logic_vector(1 downto 0);
    signal VN1212_in1 : std_logic_vector(1 downto 0);
    signal VN1212_in2 : std_logic_vector(1 downto 0);
    signal VN1212_in3 : std_logic_vector(1 downto 0);
    signal VN1212_in4 : std_logic_vector(1 downto 0);
    signal VN1212_in5 : std_logic_vector(1 downto 0);
    signal VN1213_in0 : std_logic_vector(1 downto 0);
    signal VN1213_in1 : std_logic_vector(1 downto 0);
    signal VN1213_in2 : std_logic_vector(1 downto 0);
    signal VN1213_in3 : std_logic_vector(1 downto 0);
    signal VN1213_in4 : std_logic_vector(1 downto 0);
    signal VN1213_in5 : std_logic_vector(1 downto 0);
    signal VN1214_in0 : std_logic_vector(1 downto 0);
    signal VN1214_in1 : std_logic_vector(1 downto 0);
    signal VN1214_in2 : std_logic_vector(1 downto 0);
    signal VN1214_in3 : std_logic_vector(1 downto 0);
    signal VN1214_in4 : std_logic_vector(1 downto 0);
    signal VN1214_in5 : std_logic_vector(1 downto 0);
    signal VN1215_in0 : std_logic_vector(1 downto 0);
    signal VN1215_in1 : std_logic_vector(1 downto 0);
    signal VN1215_in2 : std_logic_vector(1 downto 0);
    signal VN1215_in3 : std_logic_vector(1 downto 0);
    signal VN1215_in4 : std_logic_vector(1 downto 0);
    signal VN1215_in5 : std_logic_vector(1 downto 0);
    signal VN1216_in0 : std_logic_vector(1 downto 0);
    signal VN1216_in1 : std_logic_vector(1 downto 0);
    signal VN1216_in2 : std_logic_vector(1 downto 0);
    signal VN1216_in3 : std_logic_vector(1 downto 0);
    signal VN1216_in4 : std_logic_vector(1 downto 0);
    signal VN1216_in5 : std_logic_vector(1 downto 0);
    signal VN1217_in0 : std_logic_vector(1 downto 0);
    signal VN1217_in1 : std_logic_vector(1 downto 0);
    signal VN1217_in2 : std_logic_vector(1 downto 0);
    signal VN1217_in3 : std_logic_vector(1 downto 0);
    signal VN1217_in4 : std_logic_vector(1 downto 0);
    signal VN1217_in5 : std_logic_vector(1 downto 0);
    signal VN1218_in0 : std_logic_vector(1 downto 0);
    signal VN1218_in1 : std_logic_vector(1 downto 0);
    signal VN1218_in2 : std_logic_vector(1 downto 0);
    signal VN1218_in3 : std_logic_vector(1 downto 0);
    signal VN1218_in4 : std_logic_vector(1 downto 0);
    signal VN1218_in5 : std_logic_vector(1 downto 0);
    signal VN1219_in0 : std_logic_vector(1 downto 0);
    signal VN1219_in1 : std_logic_vector(1 downto 0);
    signal VN1219_in2 : std_logic_vector(1 downto 0);
    signal VN1219_in3 : std_logic_vector(1 downto 0);
    signal VN1219_in4 : std_logic_vector(1 downto 0);
    signal VN1219_in5 : std_logic_vector(1 downto 0);
    signal VN1220_in0 : std_logic_vector(1 downto 0);
    signal VN1220_in1 : std_logic_vector(1 downto 0);
    signal VN1220_in2 : std_logic_vector(1 downto 0);
    signal VN1220_in3 : std_logic_vector(1 downto 0);
    signal VN1220_in4 : std_logic_vector(1 downto 0);
    signal VN1220_in5 : std_logic_vector(1 downto 0);
    signal VN1221_in0 : std_logic_vector(1 downto 0);
    signal VN1221_in1 : std_logic_vector(1 downto 0);
    signal VN1221_in2 : std_logic_vector(1 downto 0);
    signal VN1221_in3 : std_logic_vector(1 downto 0);
    signal VN1221_in4 : std_logic_vector(1 downto 0);
    signal VN1221_in5 : std_logic_vector(1 downto 0);
    signal VN1222_in0 : std_logic_vector(1 downto 0);
    signal VN1222_in1 : std_logic_vector(1 downto 0);
    signal VN1222_in2 : std_logic_vector(1 downto 0);
    signal VN1222_in3 : std_logic_vector(1 downto 0);
    signal VN1222_in4 : std_logic_vector(1 downto 0);
    signal VN1222_in5 : std_logic_vector(1 downto 0);
    signal VN1223_in0 : std_logic_vector(1 downto 0);
    signal VN1223_in1 : std_logic_vector(1 downto 0);
    signal VN1223_in2 : std_logic_vector(1 downto 0);
    signal VN1223_in3 : std_logic_vector(1 downto 0);
    signal VN1223_in4 : std_logic_vector(1 downto 0);
    signal VN1223_in5 : std_logic_vector(1 downto 0);
    signal VN1224_in0 : std_logic_vector(1 downto 0);
    signal VN1224_in1 : std_logic_vector(1 downto 0);
    signal VN1224_in2 : std_logic_vector(1 downto 0);
    signal VN1224_in3 : std_logic_vector(1 downto 0);
    signal VN1224_in4 : std_logic_vector(1 downto 0);
    signal VN1224_in5 : std_logic_vector(1 downto 0);
    signal VN1225_in0 : std_logic_vector(1 downto 0);
    signal VN1225_in1 : std_logic_vector(1 downto 0);
    signal VN1225_in2 : std_logic_vector(1 downto 0);
    signal VN1225_in3 : std_logic_vector(1 downto 0);
    signal VN1225_in4 : std_logic_vector(1 downto 0);
    signal VN1225_in5 : std_logic_vector(1 downto 0);
    signal VN1226_in0 : std_logic_vector(1 downto 0);
    signal VN1226_in1 : std_logic_vector(1 downto 0);
    signal VN1226_in2 : std_logic_vector(1 downto 0);
    signal VN1226_in3 : std_logic_vector(1 downto 0);
    signal VN1226_in4 : std_logic_vector(1 downto 0);
    signal VN1226_in5 : std_logic_vector(1 downto 0);
    signal VN1227_in0 : std_logic_vector(1 downto 0);
    signal VN1227_in1 : std_logic_vector(1 downto 0);
    signal VN1227_in2 : std_logic_vector(1 downto 0);
    signal VN1227_in3 : std_logic_vector(1 downto 0);
    signal VN1227_in4 : std_logic_vector(1 downto 0);
    signal VN1227_in5 : std_logic_vector(1 downto 0);
    signal VN1228_in0 : std_logic_vector(1 downto 0);
    signal VN1228_in1 : std_logic_vector(1 downto 0);
    signal VN1228_in2 : std_logic_vector(1 downto 0);
    signal VN1228_in3 : std_logic_vector(1 downto 0);
    signal VN1228_in4 : std_logic_vector(1 downto 0);
    signal VN1228_in5 : std_logic_vector(1 downto 0);
    signal VN1229_in0 : std_logic_vector(1 downto 0);
    signal VN1229_in1 : std_logic_vector(1 downto 0);
    signal VN1229_in2 : std_logic_vector(1 downto 0);
    signal VN1229_in3 : std_logic_vector(1 downto 0);
    signal VN1229_in4 : std_logic_vector(1 downto 0);
    signal VN1229_in5 : std_logic_vector(1 downto 0);
    signal VN1230_in0 : std_logic_vector(1 downto 0);
    signal VN1230_in1 : std_logic_vector(1 downto 0);
    signal VN1230_in2 : std_logic_vector(1 downto 0);
    signal VN1230_in3 : std_logic_vector(1 downto 0);
    signal VN1230_in4 : std_logic_vector(1 downto 0);
    signal VN1230_in5 : std_logic_vector(1 downto 0);
    signal VN1231_in0 : std_logic_vector(1 downto 0);
    signal VN1231_in1 : std_logic_vector(1 downto 0);
    signal VN1231_in2 : std_logic_vector(1 downto 0);
    signal VN1231_in3 : std_logic_vector(1 downto 0);
    signal VN1231_in4 : std_logic_vector(1 downto 0);
    signal VN1231_in5 : std_logic_vector(1 downto 0);
    signal VN1232_in0 : std_logic_vector(1 downto 0);
    signal VN1232_in1 : std_logic_vector(1 downto 0);
    signal VN1232_in2 : std_logic_vector(1 downto 0);
    signal VN1232_in3 : std_logic_vector(1 downto 0);
    signal VN1232_in4 : std_logic_vector(1 downto 0);
    signal VN1232_in5 : std_logic_vector(1 downto 0);
    signal VN1233_in0 : std_logic_vector(1 downto 0);
    signal VN1233_in1 : std_logic_vector(1 downto 0);
    signal VN1233_in2 : std_logic_vector(1 downto 0);
    signal VN1233_in3 : std_logic_vector(1 downto 0);
    signal VN1233_in4 : std_logic_vector(1 downto 0);
    signal VN1233_in5 : std_logic_vector(1 downto 0);
    signal VN1234_in0 : std_logic_vector(1 downto 0);
    signal VN1234_in1 : std_logic_vector(1 downto 0);
    signal VN1234_in2 : std_logic_vector(1 downto 0);
    signal VN1234_in3 : std_logic_vector(1 downto 0);
    signal VN1234_in4 : std_logic_vector(1 downto 0);
    signal VN1234_in5 : std_logic_vector(1 downto 0);
    signal VN1235_in0 : std_logic_vector(1 downto 0);
    signal VN1235_in1 : std_logic_vector(1 downto 0);
    signal VN1235_in2 : std_logic_vector(1 downto 0);
    signal VN1235_in3 : std_logic_vector(1 downto 0);
    signal VN1235_in4 : std_logic_vector(1 downto 0);
    signal VN1235_in5 : std_logic_vector(1 downto 0);
    signal VN1236_in0 : std_logic_vector(1 downto 0);
    signal VN1236_in1 : std_logic_vector(1 downto 0);
    signal VN1236_in2 : std_logic_vector(1 downto 0);
    signal VN1236_in3 : std_logic_vector(1 downto 0);
    signal VN1236_in4 : std_logic_vector(1 downto 0);
    signal VN1236_in5 : std_logic_vector(1 downto 0);
    signal VN1237_in0 : std_logic_vector(1 downto 0);
    signal VN1237_in1 : std_logic_vector(1 downto 0);
    signal VN1237_in2 : std_logic_vector(1 downto 0);
    signal VN1237_in3 : std_logic_vector(1 downto 0);
    signal VN1237_in4 : std_logic_vector(1 downto 0);
    signal VN1237_in5 : std_logic_vector(1 downto 0);
    signal VN1238_in0 : std_logic_vector(1 downto 0);
    signal VN1238_in1 : std_logic_vector(1 downto 0);
    signal VN1238_in2 : std_logic_vector(1 downto 0);
    signal VN1238_in3 : std_logic_vector(1 downto 0);
    signal VN1238_in4 : std_logic_vector(1 downto 0);
    signal VN1238_in5 : std_logic_vector(1 downto 0);
    signal VN1239_in0 : std_logic_vector(1 downto 0);
    signal VN1239_in1 : std_logic_vector(1 downto 0);
    signal VN1239_in2 : std_logic_vector(1 downto 0);
    signal VN1239_in3 : std_logic_vector(1 downto 0);
    signal VN1239_in4 : std_logic_vector(1 downto 0);
    signal VN1239_in5 : std_logic_vector(1 downto 0);
    signal VN1240_in0 : std_logic_vector(1 downto 0);
    signal VN1240_in1 : std_logic_vector(1 downto 0);
    signal VN1240_in2 : std_logic_vector(1 downto 0);
    signal VN1240_in3 : std_logic_vector(1 downto 0);
    signal VN1240_in4 : std_logic_vector(1 downto 0);
    signal VN1240_in5 : std_logic_vector(1 downto 0);
    signal VN1241_in0 : std_logic_vector(1 downto 0);
    signal VN1241_in1 : std_logic_vector(1 downto 0);
    signal VN1241_in2 : std_logic_vector(1 downto 0);
    signal VN1241_in3 : std_logic_vector(1 downto 0);
    signal VN1241_in4 : std_logic_vector(1 downto 0);
    signal VN1241_in5 : std_logic_vector(1 downto 0);
    signal VN1242_in0 : std_logic_vector(1 downto 0);
    signal VN1242_in1 : std_logic_vector(1 downto 0);
    signal VN1242_in2 : std_logic_vector(1 downto 0);
    signal VN1242_in3 : std_logic_vector(1 downto 0);
    signal VN1242_in4 : std_logic_vector(1 downto 0);
    signal VN1242_in5 : std_logic_vector(1 downto 0);
    signal VN1243_in0 : std_logic_vector(1 downto 0);
    signal VN1243_in1 : std_logic_vector(1 downto 0);
    signal VN1243_in2 : std_logic_vector(1 downto 0);
    signal VN1243_in3 : std_logic_vector(1 downto 0);
    signal VN1243_in4 : std_logic_vector(1 downto 0);
    signal VN1243_in5 : std_logic_vector(1 downto 0);
    signal VN1244_in0 : std_logic_vector(1 downto 0);
    signal VN1244_in1 : std_logic_vector(1 downto 0);
    signal VN1244_in2 : std_logic_vector(1 downto 0);
    signal VN1244_in3 : std_logic_vector(1 downto 0);
    signal VN1244_in4 : std_logic_vector(1 downto 0);
    signal VN1244_in5 : std_logic_vector(1 downto 0);
    signal VN1245_in0 : std_logic_vector(1 downto 0);
    signal VN1245_in1 : std_logic_vector(1 downto 0);
    signal VN1245_in2 : std_logic_vector(1 downto 0);
    signal VN1245_in3 : std_logic_vector(1 downto 0);
    signal VN1245_in4 : std_logic_vector(1 downto 0);
    signal VN1245_in5 : std_logic_vector(1 downto 0);
    signal VN1246_in0 : std_logic_vector(1 downto 0);
    signal VN1246_in1 : std_logic_vector(1 downto 0);
    signal VN1246_in2 : std_logic_vector(1 downto 0);
    signal VN1246_in3 : std_logic_vector(1 downto 0);
    signal VN1246_in4 : std_logic_vector(1 downto 0);
    signal VN1246_in5 : std_logic_vector(1 downto 0);
    signal VN1247_in0 : std_logic_vector(1 downto 0);
    signal VN1247_in1 : std_logic_vector(1 downto 0);
    signal VN1247_in2 : std_logic_vector(1 downto 0);
    signal VN1247_in3 : std_logic_vector(1 downto 0);
    signal VN1247_in4 : std_logic_vector(1 downto 0);
    signal VN1247_in5 : std_logic_vector(1 downto 0);
    signal VN1248_in0 : std_logic_vector(1 downto 0);
    signal VN1248_in1 : std_logic_vector(1 downto 0);
    signal VN1248_in2 : std_logic_vector(1 downto 0);
    signal VN1248_in3 : std_logic_vector(1 downto 0);
    signal VN1248_in4 : std_logic_vector(1 downto 0);
    signal VN1248_in5 : std_logic_vector(1 downto 0);
    signal VN1249_in0 : std_logic_vector(1 downto 0);
    signal VN1249_in1 : std_logic_vector(1 downto 0);
    signal VN1249_in2 : std_logic_vector(1 downto 0);
    signal VN1249_in3 : std_logic_vector(1 downto 0);
    signal VN1249_in4 : std_logic_vector(1 downto 0);
    signal VN1249_in5 : std_logic_vector(1 downto 0);
    signal VN1250_in0 : std_logic_vector(1 downto 0);
    signal VN1250_in1 : std_logic_vector(1 downto 0);
    signal VN1250_in2 : std_logic_vector(1 downto 0);
    signal VN1250_in3 : std_logic_vector(1 downto 0);
    signal VN1250_in4 : std_logic_vector(1 downto 0);
    signal VN1250_in5 : std_logic_vector(1 downto 0);
    signal VN1251_in0 : std_logic_vector(1 downto 0);
    signal VN1251_in1 : std_logic_vector(1 downto 0);
    signal VN1251_in2 : std_logic_vector(1 downto 0);
    signal VN1251_in3 : std_logic_vector(1 downto 0);
    signal VN1251_in4 : std_logic_vector(1 downto 0);
    signal VN1251_in5 : std_logic_vector(1 downto 0);
    signal VN1252_in0 : std_logic_vector(1 downto 0);
    signal VN1252_in1 : std_logic_vector(1 downto 0);
    signal VN1252_in2 : std_logic_vector(1 downto 0);
    signal VN1252_in3 : std_logic_vector(1 downto 0);
    signal VN1252_in4 : std_logic_vector(1 downto 0);
    signal VN1252_in5 : std_logic_vector(1 downto 0);
    signal VN1253_in0 : std_logic_vector(1 downto 0);
    signal VN1253_in1 : std_logic_vector(1 downto 0);
    signal VN1253_in2 : std_logic_vector(1 downto 0);
    signal VN1253_in3 : std_logic_vector(1 downto 0);
    signal VN1253_in4 : std_logic_vector(1 downto 0);
    signal VN1253_in5 : std_logic_vector(1 downto 0);
    signal VN1254_in0 : std_logic_vector(1 downto 0);
    signal VN1254_in1 : std_logic_vector(1 downto 0);
    signal VN1254_in2 : std_logic_vector(1 downto 0);
    signal VN1254_in3 : std_logic_vector(1 downto 0);
    signal VN1254_in4 : std_logic_vector(1 downto 0);
    signal VN1254_in5 : std_logic_vector(1 downto 0);
    signal VN1255_in0 : std_logic_vector(1 downto 0);
    signal VN1255_in1 : std_logic_vector(1 downto 0);
    signal VN1255_in2 : std_logic_vector(1 downto 0);
    signal VN1255_in3 : std_logic_vector(1 downto 0);
    signal VN1255_in4 : std_logic_vector(1 downto 0);
    signal VN1255_in5 : std_logic_vector(1 downto 0);
    signal VN1256_in0 : std_logic_vector(1 downto 0);
    signal VN1256_in1 : std_logic_vector(1 downto 0);
    signal VN1256_in2 : std_logic_vector(1 downto 0);
    signal VN1256_in3 : std_logic_vector(1 downto 0);
    signal VN1256_in4 : std_logic_vector(1 downto 0);
    signal VN1256_in5 : std_logic_vector(1 downto 0);
    signal VN1257_in0 : std_logic_vector(1 downto 0);
    signal VN1257_in1 : std_logic_vector(1 downto 0);
    signal VN1257_in2 : std_logic_vector(1 downto 0);
    signal VN1257_in3 : std_logic_vector(1 downto 0);
    signal VN1257_in4 : std_logic_vector(1 downto 0);
    signal VN1257_in5 : std_logic_vector(1 downto 0);
    signal VN1258_in0 : std_logic_vector(1 downto 0);
    signal VN1258_in1 : std_logic_vector(1 downto 0);
    signal VN1258_in2 : std_logic_vector(1 downto 0);
    signal VN1258_in3 : std_logic_vector(1 downto 0);
    signal VN1258_in4 : std_logic_vector(1 downto 0);
    signal VN1258_in5 : std_logic_vector(1 downto 0);
    signal VN1259_in0 : std_logic_vector(1 downto 0);
    signal VN1259_in1 : std_logic_vector(1 downto 0);
    signal VN1259_in2 : std_logic_vector(1 downto 0);
    signal VN1259_in3 : std_logic_vector(1 downto 0);
    signal VN1259_in4 : std_logic_vector(1 downto 0);
    signal VN1259_in5 : std_logic_vector(1 downto 0);
    signal VN1260_in0 : std_logic_vector(1 downto 0);
    signal VN1260_in1 : std_logic_vector(1 downto 0);
    signal VN1260_in2 : std_logic_vector(1 downto 0);
    signal VN1260_in3 : std_logic_vector(1 downto 0);
    signal VN1260_in4 : std_logic_vector(1 downto 0);
    signal VN1260_in5 : std_logic_vector(1 downto 0);
    signal VN1261_in0 : std_logic_vector(1 downto 0);
    signal VN1261_in1 : std_logic_vector(1 downto 0);
    signal VN1261_in2 : std_logic_vector(1 downto 0);
    signal VN1261_in3 : std_logic_vector(1 downto 0);
    signal VN1261_in4 : std_logic_vector(1 downto 0);
    signal VN1261_in5 : std_logic_vector(1 downto 0);
    signal VN1262_in0 : std_logic_vector(1 downto 0);
    signal VN1262_in1 : std_logic_vector(1 downto 0);
    signal VN1262_in2 : std_logic_vector(1 downto 0);
    signal VN1262_in3 : std_logic_vector(1 downto 0);
    signal VN1262_in4 : std_logic_vector(1 downto 0);
    signal VN1262_in5 : std_logic_vector(1 downto 0);
    signal VN1263_in0 : std_logic_vector(1 downto 0);
    signal VN1263_in1 : std_logic_vector(1 downto 0);
    signal VN1263_in2 : std_logic_vector(1 downto 0);
    signal VN1263_in3 : std_logic_vector(1 downto 0);
    signal VN1263_in4 : std_logic_vector(1 downto 0);
    signal VN1263_in5 : std_logic_vector(1 downto 0);
    signal VN1264_in0 : std_logic_vector(1 downto 0);
    signal VN1264_in1 : std_logic_vector(1 downto 0);
    signal VN1264_in2 : std_logic_vector(1 downto 0);
    signal VN1264_in3 : std_logic_vector(1 downto 0);
    signal VN1264_in4 : std_logic_vector(1 downto 0);
    signal VN1264_in5 : std_logic_vector(1 downto 0);
    signal VN1265_in0 : std_logic_vector(1 downto 0);
    signal VN1265_in1 : std_logic_vector(1 downto 0);
    signal VN1265_in2 : std_logic_vector(1 downto 0);
    signal VN1265_in3 : std_logic_vector(1 downto 0);
    signal VN1265_in4 : std_logic_vector(1 downto 0);
    signal VN1265_in5 : std_logic_vector(1 downto 0);
    signal VN1266_in0 : std_logic_vector(1 downto 0);
    signal VN1266_in1 : std_logic_vector(1 downto 0);
    signal VN1266_in2 : std_logic_vector(1 downto 0);
    signal VN1266_in3 : std_logic_vector(1 downto 0);
    signal VN1266_in4 : std_logic_vector(1 downto 0);
    signal VN1266_in5 : std_logic_vector(1 downto 0);
    signal VN1267_in0 : std_logic_vector(1 downto 0);
    signal VN1267_in1 : std_logic_vector(1 downto 0);
    signal VN1267_in2 : std_logic_vector(1 downto 0);
    signal VN1267_in3 : std_logic_vector(1 downto 0);
    signal VN1267_in4 : std_logic_vector(1 downto 0);
    signal VN1267_in5 : std_logic_vector(1 downto 0);
    signal VN1268_in0 : std_logic_vector(1 downto 0);
    signal VN1268_in1 : std_logic_vector(1 downto 0);
    signal VN1268_in2 : std_logic_vector(1 downto 0);
    signal VN1268_in3 : std_logic_vector(1 downto 0);
    signal VN1268_in4 : std_logic_vector(1 downto 0);
    signal VN1268_in5 : std_logic_vector(1 downto 0);
    signal VN1269_in0 : std_logic_vector(1 downto 0);
    signal VN1269_in1 : std_logic_vector(1 downto 0);
    signal VN1269_in2 : std_logic_vector(1 downto 0);
    signal VN1269_in3 : std_logic_vector(1 downto 0);
    signal VN1269_in4 : std_logic_vector(1 downto 0);
    signal VN1269_in5 : std_logic_vector(1 downto 0);
    signal VN1270_in0 : std_logic_vector(1 downto 0);
    signal VN1270_in1 : std_logic_vector(1 downto 0);
    signal VN1270_in2 : std_logic_vector(1 downto 0);
    signal VN1270_in3 : std_logic_vector(1 downto 0);
    signal VN1270_in4 : std_logic_vector(1 downto 0);
    signal VN1270_in5 : std_logic_vector(1 downto 0);
    signal VN1271_in0 : std_logic_vector(1 downto 0);
    signal VN1271_in1 : std_logic_vector(1 downto 0);
    signal VN1271_in2 : std_logic_vector(1 downto 0);
    signal VN1271_in3 : std_logic_vector(1 downto 0);
    signal VN1271_in4 : std_logic_vector(1 downto 0);
    signal VN1271_in5 : std_logic_vector(1 downto 0);
    signal VN1272_in0 : std_logic_vector(1 downto 0);
    signal VN1272_in1 : std_logic_vector(1 downto 0);
    signal VN1272_in2 : std_logic_vector(1 downto 0);
    signal VN1272_in3 : std_logic_vector(1 downto 0);
    signal VN1272_in4 : std_logic_vector(1 downto 0);
    signal VN1272_in5 : std_logic_vector(1 downto 0);
    signal VN1273_in0 : std_logic_vector(1 downto 0);
    signal VN1273_in1 : std_logic_vector(1 downto 0);
    signal VN1273_in2 : std_logic_vector(1 downto 0);
    signal VN1273_in3 : std_logic_vector(1 downto 0);
    signal VN1273_in4 : std_logic_vector(1 downto 0);
    signal VN1273_in5 : std_logic_vector(1 downto 0);
    signal VN1274_in0 : std_logic_vector(1 downto 0);
    signal VN1274_in1 : std_logic_vector(1 downto 0);
    signal VN1274_in2 : std_logic_vector(1 downto 0);
    signal VN1274_in3 : std_logic_vector(1 downto 0);
    signal VN1274_in4 : std_logic_vector(1 downto 0);
    signal VN1274_in5 : std_logic_vector(1 downto 0);
    signal VN1275_in0 : std_logic_vector(1 downto 0);
    signal VN1275_in1 : std_logic_vector(1 downto 0);
    signal VN1275_in2 : std_logic_vector(1 downto 0);
    signal VN1275_in3 : std_logic_vector(1 downto 0);
    signal VN1275_in4 : std_logic_vector(1 downto 0);
    signal VN1275_in5 : std_logic_vector(1 downto 0);
    signal VN1276_in0 : std_logic_vector(1 downto 0);
    signal VN1276_in1 : std_logic_vector(1 downto 0);
    signal VN1276_in2 : std_logic_vector(1 downto 0);
    signal VN1276_in3 : std_logic_vector(1 downto 0);
    signal VN1276_in4 : std_logic_vector(1 downto 0);
    signal VN1276_in5 : std_logic_vector(1 downto 0);
    signal VN1277_in0 : std_logic_vector(1 downto 0);
    signal VN1277_in1 : std_logic_vector(1 downto 0);
    signal VN1277_in2 : std_logic_vector(1 downto 0);
    signal VN1277_in3 : std_logic_vector(1 downto 0);
    signal VN1277_in4 : std_logic_vector(1 downto 0);
    signal VN1277_in5 : std_logic_vector(1 downto 0);
    signal VN1278_in0 : std_logic_vector(1 downto 0);
    signal VN1278_in1 : std_logic_vector(1 downto 0);
    signal VN1278_in2 : std_logic_vector(1 downto 0);
    signal VN1278_in3 : std_logic_vector(1 downto 0);
    signal VN1278_in4 : std_logic_vector(1 downto 0);
    signal VN1278_in5 : std_logic_vector(1 downto 0);
    signal VN1279_in0 : std_logic_vector(1 downto 0);
    signal VN1279_in1 : std_logic_vector(1 downto 0);
    signal VN1279_in2 : std_logic_vector(1 downto 0);
    signal VN1279_in3 : std_logic_vector(1 downto 0);
    signal VN1279_in4 : std_logic_vector(1 downto 0);
    signal VN1279_in5 : std_logic_vector(1 downto 0);
    signal VN1280_in0 : std_logic_vector(1 downto 0);
    signal VN1280_in1 : std_logic_vector(1 downto 0);
    signal VN1280_in2 : std_logic_vector(1 downto 0);
    signal VN1280_in3 : std_logic_vector(1 downto 0);
    signal VN1280_in4 : std_logic_vector(1 downto 0);
    signal VN1280_in5 : std_logic_vector(1 downto 0);
    signal VN1281_in0 : std_logic_vector(1 downto 0);
    signal VN1281_in1 : std_logic_vector(1 downto 0);
    signal VN1281_in2 : std_logic_vector(1 downto 0);
    signal VN1281_in3 : std_logic_vector(1 downto 0);
    signal VN1281_in4 : std_logic_vector(1 downto 0);
    signal VN1281_in5 : std_logic_vector(1 downto 0);
    signal VN1282_in0 : std_logic_vector(1 downto 0);
    signal VN1282_in1 : std_logic_vector(1 downto 0);
    signal VN1282_in2 : std_logic_vector(1 downto 0);
    signal VN1282_in3 : std_logic_vector(1 downto 0);
    signal VN1282_in4 : std_logic_vector(1 downto 0);
    signal VN1282_in5 : std_logic_vector(1 downto 0);
    signal VN1283_in0 : std_logic_vector(1 downto 0);
    signal VN1283_in1 : std_logic_vector(1 downto 0);
    signal VN1283_in2 : std_logic_vector(1 downto 0);
    signal VN1283_in3 : std_logic_vector(1 downto 0);
    signal VN1283_in4 : std_logic_vector(1 downto 0);
    signal VN1283_in5 : std_logic_vector(1 downto 0);
    signal VN1284_in0 : std_logic_vector(1 downto 0);
    signal VN1284_in1 : std_logic_vector(1 downto 0);
    signal VN1284_in2 : std_logic_vector(1 downto 0);
    signal VN1284_in3 : std_logic_vector(1 downto 0);
    signal VN1284_in4 : std_logic_vector(1 downto 0);
    signal VN1284_in5 : std_logic_vector(1 downto 0);
    signal VN1285_in0 : std_logic_vector(1 downto 0);
    signal VN1285_in1 : std_logic_vector(1 downto 0);
    signal VN1285_in2 : std_logic_vector(1 downto 0);
    signal VN1285_in3 : std_logic_vector(1 downto 0);
    signal VN1285_in4 : std_logic_vector(1 downto 0);
    signal VN1285_in5 : std_logic_vector(1 downto 0);
    signal VN1286_in0 : std_logic_vector(1 downto 0);
    signal VN1286_in1 : std_logic_vector(1 downto 0);
    signal VN1286_in2 : std_logic_vector(1 downto 0);
    signal VN1286_in3 : std_logic_vector(1 downto 0);
    signal VN1286_in4 : std_logic_vector(1 downto 0);
    signal VN1286_in5 : std_logic_vector(1 downto 0);
    signal VN1287_in0 : std_logic_vector(1 downto 0);
    signal VN1287_in1 : std_logic_vector(1 downto 0);
    signal VN1287_in2 : std_logic_vector(1 downto 0);
    signal VN1287_in3 : std_logic_vector(1 downto 0);
    signal VN1287_in4 : std_logic_vector(1 downto 0);
    signal VN1287_in5 : std_logic_vector(1 downto 0);
    signal VN1288_in0 : std_logic_vector(1 downto 0);
    signal VN1288_in1 : std_logic_vector(1 downto 0);
    signal VN1288_in2 : std_logic_vector(1 downto 0);
    signal VN1288_in3 : std_logic_vector(1 downto 0);
    signal VN1288_in4 : std_logic_vector(1 downto 0);
    signal VN1288_in5 : std_logic_vector(1 downto 0);
    signal VN1289_in0 : std_logic_vector(1 downto 0);
    signal VN1289_in1 : std_logic_vector(1 downto 0);
    signal VN1289_in2 : std_logic_vector(1 downto 0);
    signal VN1289_in3 : std_logic_vector(1 downto 0);
    signal VN1289_in4 : std_logic_vector(1 downto 0);
    signal VN1289_in5 : std_logic_vector(1 downto 0);
    signal VN1290_in0 : std_logic_vector(1 downto 0);
    signal VN1290_in1 : std_logic_vector(1 downto 0);
    signal VN1290_in2 : std_logic_vector(1 downto 0);
    signal VN1290_in3 : std_logic_vector(1 downto 0);
    signal VN1290_in4 : std_logic_vector(1 downto 0);
    signal VN1290_in5 : std_logic_vector(1 downto 0);
    signal VN1291_in0 : std_logic_vector(1 downto 0);
    signal VN1291_in1 : std_logic_vector(1 downto 0);
    signal VN1291_in2 : std_logic_vector(1 downto 0);
    signal VN1291_in3 : std_logic_vector(1 downto 0);
    signal VN1291_in4 : std_logic_vector(1 downto 0);
    signal VN1291_in5 : std_logic_vector(1 downto 0);
    signal VN1292_in0 : std_logic_vector(1 downto 0);
    signal VN1292_in1 : std_logic_vector(1 downto 0);
    signal VN1292_in2 : std_logic_vector(1 downto 0);
    signal VN1292_in3 : std_logic_vector(1 downto 0);
    signal VN1292_in4 : std_logic_vector(1 downto 0);
    signal VN1292_in5 : std_logic_vector(1 downto 0);
    signal VN1293_in0 : std_logic_vector(1 downto 0);
    signal VN1293_in1 : std_logic_vector(1 downto 0);
    signal VN1293_in2 : std_logic_vector(1 downto 0);
    signal VN1293_in3 : std_logic_vector(1 downto 0);
    signal VN1293_in4 : std_logic_vector(1 downto 0);
    signal VN1293_in5 : std_logic_vector(1 downto 0);
    signal VN1294_in0 : std_logic_vector(1 downto 0);
    signal VN1294_in1 : std_logic_vector(1 downto 0);
    signal VN1294_in2 : std_logic_vector(1 downto 0);
    signal VN1294_in3 : std_logic_vector(1 downto 0);
    signal VN1294_in4 : std_logic_vector(1 downto 0);
    signal VN1294_in5 : std_logic_vector(1 downto 0);
    signal VN1295_in0 : std_logic_vector(1 downto 0);
    signal VN1295_in1 : std_logic_vector(1 downto 0);
    signal VN1295_in2 : std_logic_vector(1 downto 0);
    signal VN1295_in3 : std_logic_vector(1 downto 0);
    signal VN1295_in4 : std_logic_vector(1 downto 0);
    signal VN1295_in5 : std_logic_vector(1 downto 0);
    signal VN1296_in0 : std_logic_vector(1 downto 0);
    signal VN1296_in1 : std_logic_vector(1 downto 0);
    signal VN1296_in2 : std_logic_vector(1 downto 0);
    signal VN1296_in3 : std_logic_vector(1 downto 0);
    signal VN1296_in4 : std_logic_vector(1 downto 0);
    signal VN1296_in5 : std_logic_vector(1 downto 0);
    signal VN1297_in0 : std_logic_vector(1 downto 0);
    signal VN1297_in1 : std_logic_vector(1 downto 0);
    signal VN1297_in2 : std_logic_vector(1 downto 0);
    signal VN1297_in3 : std_logic_vector(1 downto 0);
    signal VN1297_in4 : std_logic_vector(1 downto 0);
    signal VN1297_in5 : std_logic_vector(1 downto 0);
    signal VN1298_in0 : std_logic_vector(1 downto 0);
    signal VN1298_in1 : std_logic_vector(1 downto 0);
    signal VN1298_in2 : std_logic_vector(1 downto 0);
    signal VN1298_in3 : std_logic_vector(1 downto 0);
    signal VN1298_in4 : std_logic_vector(1 downto 0);
    signal VN1298_in5 : std_logic_vector(1 downto 0);
    signal VN1299_in0 : std_logic_vector(1 downto 0);
    signal VN1299_in1 : std_logic_vector(1 downto 0);
    signal VN1299_in2 : std_logic_vector(1 downto 0);
    signal VN1299_in3 : std_logic_vector(1 downto 0);
    signal VN1299_in4 : std_logic_vector(1 downto 0);
    signal VN1299_in5 : std_logic_vector(1 downto 0);
    signal VN1300_in0 : std_logic_vector(1 downto 0);
    signal VN1300_in1 : std_logic_vector(1 downto 0);
    signal VN1300_in2 : std_logic_vector(1 downto 0);
    signal VN1300_in3 : std_logic_vector(1 downto 0);
    signal VN1300_in4 : std_logic_vector(1 downto 0);
    signal VN1300_in5 : std_logic_vector(1 downto 0);
    signal VN1301_in0 : std_logic_vector(1 downto 0);
    signal VN1301_in1 : std_logic_vector(1 downto 0);
    signal VN1301_in2 : std_logic_vector(1 downto 0);
    signal VN1301_in3 : std_logic_vector(1 downto 0);
    signal VN1301_in4 : std_logic_vector(1 downto 0);
    signal VN1301_in5 : std_logic_vector(1 downto 0);
    signal VN1302_in0 : std_logic_vector(1 downto 0);
    signal VN1302_in1 : std_logic_vector(1 downto 0);
    signal VN1302_in2 : std_logic_vector(1 downto 0);
    signal VN1302_in3 : std_logic_vector(1 downto 0);
    signal VN1302_in4 : std_logic_vector(1 downto 0);
    signal VN1302_in5 : std_logic_vector(1 downto 0);
    signal VN1303_in0 : std_logic_vector(1 downto 0);
    signal VN1303_in1 : std_logic_vector(1 downto 0);
    signal VN1303_in2 : std_logic_vector(1 downto 0);
    signal VN1303_in3 : std_logic_vector(1 downto 0);
    signal VN1303_in4 : std_logic_vector(1 downto 0);
    signal VN1303_in5 : std_logic_vector(1 downto 0);
    signal VN1304_in0 : std_logic_vector(1 downto 0);
    signal VN1304_in1 : std_logic_vector(1 downto 0);
    signal VN1304_in2 : std_logic_vector(1 downto 0);
    signal VN1304_in3 : std_logic_vector(1 downto 0);
    signal VN1304_in4 : std_logic_vector(1 downto 0);
    signal VN1304_in5 : std_logic_vector(1 downto 0);
    signal VN1305_in0 : std_logic_vector(1 downto 0);
    signal VN1305_in1 : std_logic_vector(1 downto 0);
    signal VN1305_in2 : std_logic_vector(1 downto 0);
    signal VN1305_in3 : std_logic_vector(1 downto 0);
    signal VN1305_in4 : std_logic_vector(1 downto 0);
    signal VN1305_in5 : std_logic_vector(1 downto 0);
    signal VN1306_in0 : std_logic_vector(1 downto 0);
    signal VN1306_in1 : std_logic_vector(1 downto 0);
    signal VN1306_in2 : std_logic_vector(1 downto 0);
    signal VN1306_in3 : std_logic_vector(1 downto 0);
    signal VN1306_in4 : std_logic_vector(1 downto 0);
    signal VN1306_in5 : std_logic_vector(1 downto 0);
    signal VN1307_in0 : std_logic_vector(1 downto 0);
    signal VN1307_in1 : std_logic_vector(1 downto 0);
    signal VN1307_in2 : std_logic_vector(1 downto 0);
    signal VN1307_in3 : std_logic_vector(1 downto 0);
    signal VN1307_in4 : std_logic_vector(1 downto 0);
    signal VN1307_in5 : std_logic_vector(1 downto 0);
    signal VN1308_in0 : std_logic_vector(1 downto 0);
    signal VN1308_in1 : std_logic_vector(1 downto 0);
    signal VN1308_in2 : std_logic_vector(1 downto 0);
    signal VN1308_in3 : std_logic_vector(1 downto 0);
    signal VN1308_in4 : std_logic_vector(1 downto 0);
    signal VN1308_in5 : std_logic_vector(1 downto 0);
    signal VN1309_in0 : std_logic_vector(1 downto 0);
    signal VN1309_in1 : std_logic_vector(1 downto 0);
    signal VN1309_in2 : std_logic_vector(1 downto 0);
    signal VN1309_in3 : std_logic_vector(1 downto 0);
    signal VN1309_in4 : std_logic_vector(1 downto 0);
    signal VN1309_in5 : std_logic_vector(1 downto 0);
    signal VN1310_in0 : std_logic_vector(1 downto 0);
    signal VN1310_in1 : std_logic_vector(1 downto 0);
    signal VN1310_in2 : std_logic_vector(1 downto 0);
    signal VN1310_in3 : std_logic_vector(1 downto 0);
    signal VN1310_in4 : std_logic_vector(1 downto 0);
    signal VN1310_in5 : std_logic_vector(1 downto 0);
    signal VN1311_in0 : std_logic_vector(1 downto 0);
    signal VN1311_in1 : std_logic_vector(1 downto 0);
    signal VN1311_in2 : std_logic_vector(1 downto 0);
    signal VN1311_in3 : std_logic_vector(1 downto 0);
    signal VN1311_in4 : std_logic_vector(1 downto 0);
    signal VN1311_in5 : std_logic_vector(1 downto 0);
    signal VN1312_in0 : std_logic_vector(1 downto 0);
    signal VN1312_in1 : std_logic_vector(1 downto 0);
    signal VN1312_in2 : std_logic_vector(1 downto 0);
    signal VN1312_in3 : std_logic_vector(1 downto 0);
    signal VN1312_in4 : std_logic_vector(1 downto 0);
    signal VN1312_in5 : std_logic_vector(1 downto 0);
    signal VN1313_in0 : std_logic_vector(1 downto 0);
    signal VN1313_in1 : std_logic_vector(1 downto 0);
    signal VN1313_in2 : std_logic_vector(1 downto 0);
    signal VN1313_in3 : std_logic_vector(1 downto 0);
    signal VN1313_in4 : std_logic_vector(1 downto 0);
    signal VN1313_in5 : std_logic_vector(1 downto 0);
    signal VN1314_in0 : std_logic_vector(1 downto 0);
    signal VN1314_in1 : std_logic_vector(1 downto 0);
    signal VN1314_in2 : std_logic_vector(1 downto 0);
    signal VN1314_in3 : std_logic_vector(1 downto 0);
    signal VN1314_in4 : std_logic_vector(1 downto 0);
    signal VN1314_in5 : std_logic_vector(1 downto 0);
    signal VN1315_in0 : std_logic_vector(1 downto 0);
    signal VN1315_in1 : std_logic_vector(1 downto 0);
    signal VN1315_in2 : std_logic_vector(1 downto 0);
    signal VN1315_in3 : std_logic_vector(1 downto 0);
    signal VN1315_in4 : std_logic_vector(1 downto 0);
    signal VN1315_in5 : std_logic_vector(1 downto 0);
    signal VN1316_in0 : std_logic_vector(1 downto 0);
    signal VN1316_in1 : std_logic_vector(1 downto 0);
    signal VN1316_in2 : std_logic_vector(1 downto 0);
    signal VN1316_in3 : std_logic_vector(1 downto 0);
    signal VN1316_in4 : std_logic_vector(1 downto 0);
    signal VN1316_in5 : std_logic_vector(1 downto 0);
    signal VN1317_in0 : std_logic_vector(1 downto 0);
    signal VN1317_in1 : std_logic_vector(1 downto 0);
    signal VN1317_in2 : std_logic_vector(1 downto 0);
    signal VN1317_in3 : std_logic_vector(1 downto 0);
    signal VN1317_in4 : std_logic_vector(1 downto 0);
    signal VN1317_in5 : std_logic_vector(1 downto 0);
    signal VN1318_in0 : std_logic_vector(1 downto 0);
    signal VN1318_in1 : std_logic_vector(1 downto 0);
    signal VN1318_in2 : std_logic_vector(1 downto 0);
    signal VN1318_in3 : std_logic_vector(1 downto 0);
    signal VN1318_in4 : std_logic_vector(1 downto 0);
    signal VN1318_in5 : std_logic_vector(1 downto 0);
    signal VN1319_in0 : std_logic_vector(1 downto 0);
    signal VN1319_in1 : std_logic_vector(1 downto 0);
    signal VN1319_in2 : std_logic_vector(1 downto 0);
    signal VN1319_in3 : std_logic_vector(1 downto 0);
    signal VN1319_in4 : std_logic_vector(1 downto 0);
    signal VN1319_in5 : std_logic_vector(1 downto 0);
    signal VN1320_in0 : std_logic_vector(1 downto 0);
    signal VN1320_in1 : std_logic_vector(1 downto 0);
    signal VN1320_in2 : std_logic_vector(1 downto 0);
    signal VN1320_in3 : std_logic_vector(1 downto 0);
    signal VN1320_in4 : std_logic_vector(1 downto 0);
    signal VN1320_in5 : std_logic_vector(1 downto 0);
    signal VN1321_in0 : std_logic_vector(1 downto 0);
    signal VN1321_in1 : std_logic_vector(1 downto 0);
    signal VN1321_in2 : std_logic_vector(1 downto 0);
    signal VN1321_in3 : std_logic_vector(1 downto 0);
    signal VN1321_in4 : std_logic_vector(1 downto 0);
    signal VN1321_in5 : std_logic_vector(1 downto 0);
    signal VN1322_in0 : std_logic_vector(1 downto 0);
    signal VN1322_in1 : std_logic_vector(1 downto 0);
    signal VN1322_in2 : std_logic_vector(1 downto 0);
    signal VN1322_in3 : std_logic_vector(1 downto 0);
    signal VN1322_in4 : std_logic_vector(1 downto 0);
    signal VN1322_in5 : std_logic_vector(1 downto 0);
    signal VN1323_in0 : std_logic_vector(1 downto 0);
    signal VN1323_in1 : std_logic_vector(1 downto 0);
    signal VN1323_in2 : std_logic_vector(1 downto 0);
    signal VN1323_in3 : std_logic_vector(1 downto 0);
    signal VN1323_in4 : std_logic_vector(1 downto 0);
    signal VN1323_in5 : std_logic_vector(1 downto 0);
    signal VN1324_in0 : std_logic_vector(1 downto 0);
    signal VN1324_in1 : std_logic_vector(1 downto 0);
    signal VN1324_in2 : std_logic_vector(1 downto 0);
    signal VN1324_in3 : std_logic_vector(1 downto 0);
    signal VN1324_in4 : std_logic_vector(1 downto 0);
    signal VN1324_in5 : std_logic_vector(1 downto 0);
    signal VN1325_in0 : std_logic_vector(1 downto 0);
    signal VN1325_in1 : std_logic_vector(1 downto 0);
    signal VN1325_in2 : std_logic_vector(1 downto 0);
    signal VN1325_in3 : std_logic_vector(1 downto 0);
    signal VN1325_in4 : std_logic_vector(1 downto 0);
    signal VN1325_in5 : std_logic_vector(1 downto 0);
    signal VN1326_in0 : std_logic_vector(1 downto 0);
    signal VN1326_in1 : std_logic_vector(1 downto 0);
    signal VN1326_in2 : std_logic_vector(1 downto 0);
    signal VN1326_in3 : std_logic_vector(1 downto 0);
    signal VN1326_in4 : std_logic_vector(1 downto 0);
    signal VN1326_in5 : std_logic_vector(1 downto 0);
    signal VN1327_in0 : std_logic_vector(1 downto 0);
    signal VN1327_in1 : std_logic_vector(1 downto 0);
    signal VN1327_in2 : std_logic_vector(1 downto 0);
    signal VN1327_in3 : std_logic_vector(1 downto 0);
    signal VN1327_in4 : std_logic_vector(1 downto 0);
    signal VN1327_in5 : std_logic_vector(1 downto 0);
    signal VN1328_in0 : std_logic_vector(1 downto 0);
    signal VN1328_in1 : std_logic_vector(1 downto 0);
    signal VN1328_in2 : std_logic_vector(1 downto 0);
    signal VN1328_in3 : std_logic_vector(1 downto 0);
    signal VN1328_in4 : std_logic_vector(1 downto 0);
    signal VN1328_in5 : std_logic_vector(1 downto 0);
    signal VN1329_in0 : std_logic_vector(1 downto 0);
    signal VN1329_in1 : std_logic_vector(1 downto 0);
    signal VN1329_in2 : std_logic_vector(1 downto 0);
    signal VN1329_in3 : std_logic_vector(1 downto 0);
    signal VN1329_in4 : std_logic_vector(1 downto 0);
    signal VN1329_in5 : std_logic_vector(1 downto 0);
    signal VN1330_in0 : std_logic_vector(1 downto 0);
    signal VN1330_in1 : std_logic_vector(1 downto 0);
    signal VN1330_in2 : std_logic_vector(1 downto 0);
    signal VN1330_in3 : std_logic_vector(1 downto 0);
    signal VN1330_in4 : std_logic_vector(1 downto 0);
    signal VN1330_in5 : std_logic_vector(1 downto 0);
    signal VN1331_in0 : std_logic_vector(1 downto 0);
    signal VN1331_in1 : std_logic_vector(1 downto 0);
    signal VN1331_in2 : std_logic_vector(1 downto 0);
    signal VN1331_in3 : std_logic_vector(1 downto 0);
    signal VN1331_in4 : std_logic_vector(1 downto 0);
    signal VN1331_in5 : std_logic_vector(1 downto 0);
    signal VN1332_in0 : std_logic_vector(1 downto 0);
    signal VN1332_in1 : std_logic_vector(1 downto 0);
    signal VN1332_in2 : std_logic_vector(1 downto 0);
    signal VN1332_in3 : std_logic_vector(1 downto 0);
    signal VN1332_in4 : std_logic_vector(1 downto 0);
    signal VN1332_in5 : std_logic_vector(1 downto 0);
    signal VN1333_in0 : std_logic_vector(1 downto 0);
    signal VN1333_in1 : std_logic_vector(1 downto 0);
    signal VN1333_in2 : std_logic_vector(1 downto 0);
    signal VN1333_in3 : std_logic_vector(1 downto 0);
    signal VN1333_in4 : std_logic_vector(1 downto 0);
    signal VN1333_in5 : std_logic_vector(1 downto 0);
    signal VN1334_in0 : std_logic_vector(1 downto 0);
    signal VN1334_in1 : std_logic_vector(1 downto 0);
    signal VN1334_in2 : std_logic_vector(1 downto 0);
    signal VN1334_in3 : std_logic_vector(1 downto 0);
    signal VN1334_in4 : std_logic_vector(1 downto 0);
    signal VN1334_in5 : std_logic_vector(1 downto 0);
    signal VN1335_in0 : std_logic_vector(1 downto 0);
    signal VN1335_in1 : std_logic_vector(1 downto 0);
    signal VN1335_in2 : std_logic_vector(1 downto 0);
    signal VN1335_in3 : std_logic_vector(1 downto 0);
    signal VN1335_in4 : std_logic_vector(1 downto 0);
    signal VN1335_in5 : std_logic_vector(1 downto 0);
    signal VN1336_in0 : std_logic_vector(1 downto 0);
    signal VN1336_in1 : std_logic_vector(1 downto 0);
    signal VN1336_in2 : std_logic_vector(1 downto 0);
    signal VN1336_in3 : std_logic_vector(1 downto 0);
    signal VN1336_in4 : std_logic_vector(1 downto 0);
    signal VN1336_in5 : std_logic_vector(1 downto 0);
    signal VN1337_in0 : std_logic_vector(1 downto 0);
    signal VN1337_in1 : std_logic_vector(1 downto 0);
    signal VN1337_in2 : std_logic_vector(1 downto 0);
    signal VN1337_in3 : std_logic_vector(1 downto 0);
    signal VN1337_in4 : std_logic_vector(1 downto 0);
    signal VN1337_in5 : std_logic_vector(1 downto 0);
    signal VN1338_in0 : std_logic_vector(1 downto 0);
    signal VN1338_in1 : std_logic_vector(1 downto 0);
    signal VN1338_in2 : std_logic_vector(1 downto 0);
    signal VN1338_in3 : std_logic_vector(1 downto 0);
    signal VN1338_in4 : std_logic_vector(1 downto 0);
    signal VN1338_in5 : std_logic_vector(1 downto 0);
    signal VN1339_in0 : std_logic_vector(1 downto 0);
    signal VN1339_in1 : std_logic_vector(1 downto 0);
    signal VN1339_in2 : std_logic_vector(1 downto 0);
    signal VN1339_in3 : std_logic_vector(1 downto 0);
    signal VN1339_in4 : std_logic_vector(1 downto 0);
    signal VN1339_in5 : std_logic_vector(1 downto 0);
    signal VN1340_in0 : std_logic_vector(1 downto 0);
    signal VN1340_in1 : std_logic_vector(1 downto 0);
    signal VN1340_in2 : std_logic_vector(1 downto 0);
    signal VN1340_in3 : std_logic_vector(1 downto 0);
    signal VN1340_in4 : std_logic_vector(1 downto 0);
    signal VN1340_in5 : std_logic_vector(1 downto 0);
    signal VN1341_in0 : std_logic_vector(1 downto 0);
    signal VN1341_in1 : std_logic_vector(1 downto 0);
    signal VN1341_in2 : std_logic_vector(1 downto 0);
    signal VN1341_in3 : std_logic_vector(1 downto 0);
    signal VN1341_in4 : std_logic_vector(1 downto 0);
    signal VN1341_in5 : std_logic_vector(1 downto 0);
    signal VN1342_in0 : std_logic_vector(1 downto 0);
    signal VN1342_in1 : std_logic_vector(1 downto 0);
    signal VN1342_in2 : std_logic_vector(1 downto 0);
    signal VN1342_in3 : std_logic_vector(1 downto 0);
    signal VN1342_in4 : std_logic_vector(1 downto 0);
    signal VN1342_in5 : std_logic_vector(1 downto 0);
    signal VN1343_in0 : std_logic_vector(1 downto 0);
    signal VN1343_in1 : std_logic_vector(1 downto 0);
    signal VN1343_in2 : std_logic_vector(1 downto 0);
    signal VN1343_in3 : std_logic_vector(1 downto 0);
    signal VN1343_in4 : std_logic_vector(1 downto 0);
    signal VN1343_in5 : std_logic_vector(1 downto 0);
    signal VN1344_in0 : std_logic_vector(1 downto 0);
    signal VN1344_in1 : std_logic_vector(1 downto 0);
    signal VN1344_in2 : std_logic_vector(1 downto 0);
    signal VN1344_in3 : std_logic_vector(1 downto 0);
    signal VN1344_in4 : std_logic_vector(1 downto 0);
    signal VN1344_in5 : std_logic_vector(1 downto 0);
    signal VN1345_in0 : std_logic_vector(1 downto 0);
    signal VN1345_in1 : std_logic_vector(1 downto 0);
    signal VN1345_in2 : std_logic_vector(1 downto 0);
    signal VN1345_in3 : std_logic_vector(1 downto 0);
    signal VN1345_in4 : std_logic_vector(1 downto 0);
    signal VN1345_in5 : std_logic_vector(1 downto 0);
    signal VN1346_in0 : std_logic_vector(1 downto 0);
    signal VN1346_in1 : std_logic_vector(1 downto 0);
    signal VN1346_in2 : std_logic_vector(1 downto 0);
    signal VN1346_in3 : std_logic_vector(1 downto 0);
    signal VN1346_in4 : std_logic_vector(1 downto 0);
    signal VN1346_in5 : std_logic_vector(1 downto 0);
    signal VN1347_in0 : std_logic_vector(1 downto 0);
    signal VN1347_in1 : std_logic_vector(1 downto 0);
    signal VN1347_in2 : std_logic_vector(1 downto 0);
    signal VN1347_in3 : std_logic_vector(1 downto 0);
    signal VN1347_in4 : std_logic_vector(1 downto 0);
    signal VN1347_in5 : std_logic_vector(1 downto 0);
    signal VN1348_in0 : std_logic_vector(1 downto 0);
    signal VN1348_in1 : std_logic_vector(1 downto 0);
    signal VN1348_in2 : std_logic_vector(1 downto 0);
    signal VN1348_in3 : std_logic_vector(1 downto 0);
    signal VN1348_in4 : std_logic_vector(1 downto 0);
    signal VN1348_in5 : std_logic_vector(1 downto 0);
    signal VN1349_in0 : std_logic_vector(1 downto 0);
    signal VN1349_in1 : std_logic_vector(1 downto 0);
    signal VN1349_in2 : std_logic_vector(1 downto 0);
    signal VN1349_in3 : std_logic_vector(1 downto 0);
    signal VN1349_in4 : std_logic_vector(1 downto 0);
    signal VN1349_in5 : std_logic_vector(1 downto 0);
    signal VN1350_in0 : std_logic_vector(1 downto 0);
    signal VN1350_in1 : std_logic_vector(1 downto 0);
    signal VN1350_in2 : std_logic_vector(1 downto 0);
    signal VN1350_in3 : std_logic_vector(1 downto 0);
    signal VN1350_in4 : std_logic_vector(1 downto 0);
    signal VN1350_in5 : std_logic_vector(1 downto 0);
    signal VN1351_in0 : std_logic_vector(1 downto 0);
    signal VN1351_in1 : std_logic_vector(1 downto 0);
    signal VN1351_in2 : std_logic_vector(1 downto 0);
    signal VN1351_in3 : std_logic_vector(1 downto 0);
    signal VN1351_in4 : std_logic_vector(1 downto 0);
    signal VN1351_in5 : std_logic_vector(1 downto 0);
    signal VN1352_in0 : std_logic_vector(1 downto 0);
    signal VN1352_in1 : std_logic_vector(1 downto 0);
    signal VN1352_in2 : std_logic_vector(1 downto 0);
    signal VN1352_in3 : std_logic_vector(1 downto 0);
    signal VN1352_in4 : std_logic_vector(1 downto 0);
    signal VN1352_in5 : std_logic_vector(1 downto 0);
    signal VN1353_in0 : std_logic_vector(1 downto 0);
    signal VN1353_in1 : std_logic_vector(1 downto 0);
    signal VN1353_in2 : std_logic_vector(1 downto 0);
    signal VN1353_in3 : std_logic_vector(1 downto 0);
    signal VN1353_in4 : std_logic_vector(1 downto 0);
    signal VN1353_in5 : std_logic_vector(1 downto 0);
    signal VN1354_in0 : std_logic_vector(1 downto 0);
    signal VN1354_in1 : std_logic_vector(1 downto 0);
    signal VN1354_in2 : std_logic_vector(1 downto 0);
    signal VN1354_in3 : std_logic_vector(1 downto 0);
    signal VN1354_in4 : std_logic_vector(1 downto 0);
    signal VN1354_in5 : std_logic_vector(1 downto 0);
    signal VN1355_in0 : std_logic_vector(1 downto 0);
    signal VN1355_in1 : std_logic_vector(1 downto 0);
    signal VN1355_in2 : std_logic_vector(1 downto 0);
    signal VN1355_in3 : std_logic_vector(1 downto 0);
    signal VN1355_in4 : std_logic_vector(1 downto 0);
    signal VN1355_in5 : std_logic_vector(1 downto 0);
    signal VN1356_in0 : std_logic_vector(1 downto 0);
    signal VN1356_in1 : std_logic_vector(1 downto 0);
    signal VN1356_in2 : std_logic_vector(1 downto 0);
    signal VN1356_in3 : std_logic_vector(1 downto 0);
    signal VN1356_in4 : std_logic_vector(1 downto 0);
    signal VN1356_in5 : std_logic_vector(1 downto 0);
    signal VN1357_in0 : std_logic_vector(1 downto 0);
    signal VN1357_in1 : std_logic_vector(1 downto 0);
    signal VN1357_in2 : std_logic_vector(1 downto 0);
    signal VN1357_in3 : std_logic_vector(1 downto 0);
    signal VN1357_in4 : std_logic_vector(1 downto 0);
    signal VN1357_in5 : std_logic_vector(1 downto 0);
    signal VN1358_in0 : std_logic_vector(1 downto 0);
    signal VN1358_in1 : std_logic_vector(1 downto 0);
    signal VN1358_in2 : std_logic_vector(1 downto 0);
    signal VN1358_in3 : std_logic_vector(1 downto 0);
    signal VN1358_in4 : std_logic_vector(1 downto 0);
    signal VN1358_in5 : std_logic_vector(1 downto 0);
    signal VN1359_in0 : std_logic_vector(1 downto 0);
    signal VN1359_in1 : std_logic_vector(1 downto 0);
    signal VN1359_in2 : std_logic_vector(1 downto 0);
    signal VN1359_in3 : std_logic_vector(1 downto 0);
    signal VN1359_in4 : std_logic_vector(1 downto 0);
    signal VN1359_in5 : std_logic_vector(1 downto 0);
    signal VN1360_in0 : std_logic_vector(1 downto 0);
    signal VN1360_in1 : std_logic_vector(1 downto 0);
    signal VN1360_in2 : std_logic_vector(1 downto 0);
    signal VN1360_in3 : std_logic_vector(1 downto 0);
    signal VN1360_in4 : std_logic_vector(1 downto 0);
    signal VN1360_in5 : std_logic_vector(1 downto 0);
    signal VN1361_in0 : std_logic_vector(1 downto 0);
    signal VN1361_in1 : std_logic_vector(1 downto 0);
    signal VN1361_in2 : std_logic_vector(1 downto 0);
    signal VN1361_in3 : std_logic_vector(1 downto 0);
    signal VN1361_in4 : std_logic_vector(1 downto 0);
    signal VN1361_in5 : std_logic_vector(1 downto 0);
    signal VN1362_in0 : std_logic_vector(1 downto 0);
    signal VN1362_in1 : std_logic_vector(1 downto 0);
    signal VN1362_in2 : std_logic_vector(1 downto 0);
    signal VN1362_in3 : std_logic_vector(1 downto 0);
    signal VN1362_in4 : std_logic_vector(1 downto 0);
    signal VN1362_in5 : std_logic_vector(1 downto 0);
    signal VN1363_in0 : std_logic_vector(1 downto 0);
    signal VN1363_in1 : std_logic_vector(1 downto 0);
    signal VN1363_in2 : std_logic_vector(1 downto 0);
    signal VN1363_in3 : std_logic_vector(1 downto 0);
    signal VN1363_in4 : std_logic_vector(1 downto 0);
    signal VN1363_in5 : std_logic_vector(1 downto 0);
    signal VN1364_in0 : std_logic_vector(1 downto 0);
    signal VN1364_in1 : std_logic_vector(1 downto 0);
    signal VN1364_in2 : std_logic_vector(1 downto 0);
    signal VN1364_in3 : std_logic_vector(1 downto 0);
    signal VN1364_in4 : std_logic_vector(1 downto 0);
    signal VN1364_in5 : std_logic_vector(1 downto 0);
    signal VN1365_in0 : std_logic_vector(1 downto 0);
    signal VN1365_in1 : std_logic_vector(1 downto 0);
    signal VN1365_in2 : std_logic_vector(1 downto 0);
    signal VN1365_in3 : std_logic_vector(1 downto 0);
    signal VN1365_in4 : std_logic_vector(1 downto 0);
    signal VN1365_in5 : std_logic_vector(1 downto 0);
    signal VN1366_in0 : std_logic_vector(1 downto 0);
    signal VN1366_in1 : std_logic_vector(1 downto 0);
    signal VN1366_in2 : std_logic_vector(1 downto 0);
    signal VN1366_in3 : std_logic_vector(1 downto 0);
    signal VN1366_in4 : std_logic_vector(1 downto 0);
    signal VN1366_in5 : std_logic_vector(1 downto 0);
    signal VN1367_in0 : std_logic_vector(1 downto 0);
    signal VN1367_in1 : std_logic_vector(1 downto 0);
    signal VN1367_in2 : std_logic_vector(1 downto 0);
    signal VN1367_in3 : std_logic_vector(1 downto 0);
    signal VN1367_in4 : std_logic_vector(1 downto 0);
    signal VN1367_in5 : std_logic_vector(1 downto 0);
    signal VN1368_in0 : std_logic_vector(1 downto 0);
    signal VN1368_in1 : std_logic_vector(1 downto 0);
    signal VN1368_in2 : std_logic_vector(1 downto 0);
    signal VN1368_in3 : std_logic_vector(1 downto 0);
    signal VN1368_in4 : std_logic_vector(1 downto 0);
    signal VN1368_in5 : std_logic_vector(1 downto 0);
    signal VN1369_in0 : std_logic_vector(1 downto 0);
    signal VN1369_in1 : std_logic_vector(1 downto 0);
    signal VN1369_in2 : std_logic_vector(1 downto 0);
    signal VN1369_in3 : std_logic_vector(1 downto 0);
    signal VN1369_in4 : std_logic_vector(1 downto 0);
    signal VN1369_in5 : std_logic_vector(1 downto 0);
    signal VN1370_in0 : std_logic_vector(1 downto 0);
    signal VN1370_in1 : std_logic_vector(1 downto 0);
    signal VN1370_in2 : std_logic_vector(1 downto 0);
    signal VN1370_in3 : std_logic_vector(1 downto 0);
    signal VN1370_in4 : std_logic_vector(1 downto 0);
    signal VN1370_in5 : std_logic_vector(1 downto 0);
    signal VN1371_in0 : std_logic_vector(1 downto 0);
    signal VN1371_in1 : std_logic_vector(1 downto 0);
    signal VN1371_in2 : std_logic_vector(1 downto 0);
    signal VN1371_in3 : std_logic_vector(1 downto 0);
    signal VN1371_in4 : std_logic_vector(1 downto 0);
    signal VN1371_in5 : std_logic_vector(1 downto 0);
    signal VN1372_in0 : std_logic_vector(1 downto 0);
    signal VN1372_in1 : std_logic_vector(1 downto 0);
    signal VN1372_in2 : std_logic_vector(1 downto 0);
    signal VN1372_in3 : std_logic_vector(1 downto 0);
    signal VN1372_in4 : std_logic_vector(1 downto 0);
    signal VN1372_in5 : std_logic_vector(1 downto 0);
    signal VN1373_in0 : std_logic_vector(1 downto 0);
    signal VN1373_in1 : std_logic_vector(1 downto 0);
    signal VN1373_in2 : std_logic_vector(1 downto 0);
    signal VN1373_in3 : std_logic_vector(1 downto 0);
    signal VN1373_in4 : std_logic_vector(1 downto 0);
    signal VN1373_in5 : std_logic_vector(1 downto 0);
    signal VN1374_in0 : std_logic_vector(1 downto 0);
    signal VN1374_in1 : std_logic_vector(1 downto 0);
    signal VN1374_in2 : std_logic_vector(1 downto 0);
    signal VN1374_in3 : std_logic_vector(1 downto 0);
    signal VN1374_in4 : std_logic_vector(1 downto 0);
    signal VN1374_in5 : std_logic_vector(1 downto 0);
    signal VN1375_in0 : std_logic_vector(1 downto 0);
    signal VN1375_in1 : std_logic_vector(1 downto 0);
    signal VN1375_in2 : std_logic_vector(1 downto 0);
    signal VN1375_in3 : std_logic_vector(1 downto 0);
    signal VN1375_in4 : std_logic_vector(1 downto 0);
    signal VN1375_in5 : std_logic_vector(1 downto 0);
    signal VN1376_in0 : std_logic_vector(1 downto 0);
    signal VN1376_in1 : std_logic_vector(1 downto 0);
    signal VN1376_in2 : std_logic_vector(1 downto 0);
    signal VN1376_in3 : std_logic_vector(1 downto 0);
    signal VN1376_in4 : std_logic_vector(1 downto 0);
    signal VN1376_in5 : std_logic_vector(1 downto 0);
    signal VN1377_in0 : std_logic_vector(1 downto 0);
    signal VN1377_in1 : std_logic_vector(1 downto 0);
    signal VN1377_in2 : std_logic_vector(1 downto 0);
    signal VN1377_in3 : std_logic_vector(1 downto 0);
    signal VN1377_in4 : std_logic_vector(1 downto 0);
    signal VN1377_in5 : std_logic_vector(1 downto 0);
    signal VN1378_in0 : std_logic_vector(1 downto 0);
    signal VN1378_in1 : std_logic_vector(1 downto 0);
    signal VN1378_in2 : std_logic_vector(1 downto 0);
    signal VN1378_in3 : std_logic_vector(1 downto 0);
    signal VN1378_in4 : std_logic_vector(1 downto 0);
    signal VN1378_in5 : std_logic_vector(1 downto 0);
    signal VN1379_in0 : std_logic_vector(1 downto 0);
    signal VN1379_in1 : std_logic_vector(1 downto 0);
    signal VN1379_in2 : std_logic_vector(1 downto 0);
    signal VN1379_in3 : std_logic_vector(1 downto 0);
    signal VN1379_in4 : std_logic_vector(1 downto 0);
    signal VN1379_in5 : std_logic_vector(1 downto 0);
    signal VN1380_in0 : std_logic_vector(1 downto 0);
    signal VN1380_in1 : std_logic_vector(1 downto 0);
    signal VN1380_in2 : std_logic_vector(1 downto 0);
    signal VN1380_in3 : std_logic_vector(1 downto 0);
    signal VN1380_in4 : std_logic_vector(1 downto 0);
    signal VN1380_in5 : std_logic_vector(1 downto 0);
    signal VN1381_in0 : std_logic_vector(1 downto 0);
    signal VN1381_in1 : std_logic_vector(1 downto 0);
    signal VN1381_in2 : std_logic_vector(1 downto 0);
    signal VN1381_in3 : std_logic_vector(1 downto 0);
    signal VN1381_in4 : std_logic_vector(1 downto 0);
    signal VN1381_in5 : std_logic_vector(1 downto 0);
    signal VN1382_in0 : std_logic_vector(1 downto 0);
    signal VN1382_in1 : std_logic_vector(1 downto 0);
    signal VN1382_in2 : std_logic_vector(1 downto 0);
    signal VN1382_in3 : std_logic_vector(1 downto 0);
    signal VN1382_in4 : std_logic_vector(1 downto 0);
    signal VN1382_in5 : std_logic_vector(1 downto 0);
    signal VN1383_in0 : std_logic_vector(1 downto 0);
    signal VN1383_in1 : std_logic_vector(1 downto 0);
    signal VN1383_in2 : std_logic_vector(1 downto 0);
    signal VN1383_in3 : std_logic_vector(1 downto 0);
    signal VN1383_in4 : std_logic_vector(1 downto 0);
    signal VN1383_in5 : std_logic_vector(1 downto 0);
    signal VN1384_in0 : std_logic_vector(1 downto 0);
    signal VN1384_in1 : std_logic_vector(1 downto 0);
    signal VN1384_in2 : std_logic_vector(1 downto 0);
    signal VN1384_in3 : std_logic_vector(1 downto 0);
    signal VN1384_in4 : std_logic_vector(1 downto 0);
    signal VN1384_in5 : std_logic_vector(1 downto 0);
    signal VN1385_in0 : std_logic_vector(1 downto 0);
    signal VN1385_in1 : std_logic_vector(1 downto 0);
    signal VN1385_in2 : std_logic_vector(1 downto 0);
    signal VN1385_in3 : std_logic_vector(1 downto 0);
    signal VN1385_in4 : std_logic_vector(1 downto 0);
    signal VN1385_in5 : std_logic_vector(1 downto 0);
    signal VN1386_in0 : std_logic_vector(1 downto 0);
    signal VN1386_in1 : std_logic_vector(1 downto 0);
    signal VN1386_in2 : std_logic_vector(1 downto 0);
    signal VN1386_in3 : std_logic_vector(1 downto 0);
    signal VN1386_in4 : std_logic_vector(1 downto 0);
    signal VN1386_in5 : std_logic_vector(1 downto 0);
    signal VN1387_in0 : std_logic_vector(1 downto 0);
    signal VN1387_in1 : std_logic_vector(1 downto 0);
    signal VN1387_in2 : std_logic_vector(1 downto 0);
    signal VN1387_in3 : std_logic_vector(1 downto 0);
    signal VN1387_in4 : std_logic_vector(1 downto 0);
    signal VN1387_in5 : std_logic_vector(1 downto 0);
    signal VN1388_in0 : std_logic_vector(1 downto 0);
    signal VN1388_in1 : std_logic_vector(1 downto 0);
    signal VN1388_in2 : std_logic_vector(1 downto 0);
    signal VN1388_in3 : std_logic_vector(1 downto 0);
    signal VN1388_in4 : std_logic_vector(1 downto 0);
    signal VN1388_in5 : std_logic_vector(1 downto 0);
    signal VN1389_in0 : std_logic_vector(1 downto 0);
    signal VN1389_in1 : std_logic_vector(1 downto 0);
    signal VN1389_in2 : std_logic_vector(1 downto 0);
    signal VN1389_in3 : std_logic_vector(1 downto 0);
    signal VN1389_in4 : std_logic_vector(1 downto 0);
    signal VN1389_in5 : std_logic_vector(1 downto 0);
    signal VN1390_in0 : std_logic_vector(1 downto 0);
    signal VN1390_in1 : std_logic_vector(1 downto 0);
    signal VN1390_in2 : std_logic_vector(1 downto 0);
    signal VN1390_in3 : std_logic_vector(1 downto 0);
    signal VN1390_in4 : std_logic_vector(1 downto 0);
    signal VN1390_in5 : std_logic_vector(1 downto 0);
    signal VN1391_in0 : std_logic_vector(1 downto 0);
    signal VN1391_in1 : std_logic_vector(1 downto 0);
    signal VN1391_in2 : std_logic_vector(1 downto 0);
    signal VN1391_in3 : std_logic_vector(1 downto 0);
    signal VN1391_in4 : std_logic_vector(1 downto 0);
    signal VN1391_in5 : std_logic_vector(1 downto 0);
    signal VN1392_in0 : std_logic_vector(1 downto 0);
    signal VN1392_in1 : std_logic_vector(1 downto 0);
    signal VN1392_in2 : std_logic_vector(1 downto 0);
    signal VN1392_in3 : std_logic_vector(1 downto 0);
    signal VN1392_in4 : std_logic_vector(1 downto 0);
    signal VN1392_in5 : std_logic_vector(1 downto 0);
    signal VN1393_in0 : std_logic_vector(1 downto 0);
    signal VN1393_in1 : std_logic_vector(1 downto 0);
    signal VN1393_in2 : std_logic_vector(1 downto 0);
    signal VN1393_in3 : std_logic_vector(1 downto 0);
    signal VN1393_in4 : std_logic_vector(1 downto 0);
    signal VN1393_in5 : std_logic_vector(1 downto 0);
    signal VN1394_in0 : std_logic_vector(1 downto 0);
    signal VN1394_in1 : std_logic_vector(1 downto 0);
    signal VN1394_in2 : std_logic_vector(1 downto 0);
    signal VN1394_in3 : std_logic_vector(1 downto 0);
    signal VN1394_in4 : std_logic_vector(1 downto 0);
    signal VN1394_in5 : std_logic_vector(1 downto 0);
    signal VN1395_in0 : std_logic_vector(1 downto 0);
    signal VN1395_in1 : std_logic_vector(1 downto 0);
    signal VN1395_in2 : std_logic_vector(1 downto 0);
    signal VN1395_in3 : std_logic_vector(1 downto 0);
    signal VN1395_in4 : std_logic_vector(1 downto 0);
    signal VN1395_in5 : std_logic_vector(1 downto 0);
    signal VN1396_in0 : std_logic_vector(1 downto 0);
    signal VN1396_in1 : std_logic_vector(1 downto 0);
    signal VN1396_in2 : std_logic_vector(1 downto 0);
    signal VN1396_in3 : std_logic_vector(1 downto 0);
    signal VN1396_in4 : std_logic_vector(1 downto 0);
    signal VN1396_in5 : std_logic_vector(1 downto 0);
    signal VN1397_in0 : std_logic_vector(1 downto 0);
    signal VN1397_in1 : std_logic_vector(1 downto 0);
    signal VN1397_in2 : std_logic_vector(1 downto 0);
    signal VN1397_in3 : std_logic_vector(1 downto 0);
    signal VN1397_in4 : std_logic_vector(1 downto 0);
    signal VN1397_in5 : std_logic_vector(1 downto 0);
    signal VN1398_in0 : std_logic_vector(1 downto 0);
    signal VN1398_in1 : std_logic_vector(1 downto 0);
    signal VN1398_in2 : std_logic_vector(1 downto 0);
    signal VN1398_in3 : std_logic_vector(1 downto 0);
    signal VN1398_in4 : std_logic_vector(1 downto 0);
    signal VN1398_in5 : std_logic_vector(1 downto 0);
    signal VN1399_in0 : std_logic_vector(1 downto 0);
    signal VN1399_in1 : std_logic_vector(1 downto 0);
    signal VN1399_in2 : std_logic_vector(1 downto 0);
    signal VN1399_in3 : std_logic_vector(1 downto 0);
    signal VN1399_in4 : std_logic_vector(1 downto 0);
    signal VN1399_in5 : std_logic_vector(1 downto 0);
    signal VN1400_in0 : std_logic_vector(1 downto 0);
    signal VN1400_in1 : std_logic_vector(1 downto 0);
    signal VN1400_in2 : std_logic_vector(1 downto 0);
    signal VN1400_in3 : std_logic_vector(1 downto 0);
    signal VN1400_in4 : std_logic_vector(1 downto 0);
    signal VN1400_in5 : std_logic_vector(1 downto 0);
    signal VN1401_in0 : std_logic_vector(1 downto 0);
    signal VN1401_in1 : std_logic_vector(1 downto 0);
    signal VN1401_in2 : std_logic_vector(1 downto 0);
    signal VN1401_in3 : std_logic_vector(1 downto 0);
    signal VN1401_in4 : std_logic_vector(1 downto 0);
    signal VN1401_in5 : std_logic_vector(1 downto 0);
    signal VN1402_in0 : std_logic_vector(1 downto 0);
    signal VN1402_in1 : std_logic_vector(1 downto 0);
    signal VN1402_in2 : std_logic_vector(1 downto 0);
    signal VN1402_in3 : std_logic_vector(1 downto 0);
    signal VN1402_in4 : std_logic_vector(1 downto 0);
    signal VN1402_in5 : std_logic_vector(1 downto 0);
    signal VN1403_in0 : std_logic_vector(1 downto 0);
    signal VN1403_in1 : std_logic_vector(1 downto 0);
    signal VN1403_in2 : std_logic_vector(1 downto 0);
    signal VN1403_in3 : std_logic_vector(1 downto 0);
    signal VN1403_in4 : std_logic_vector(1 downto 0);
    signal VN1403_in5 : std_logic_vector(1 downto 0);
    signal VN1404_in0 : std_logic_vector(1 downto 0);
    signal VN1404_in1 : std_logic_vector(1 downto 0);
    signal VN1404_in2 : std_logic_vector(1 downto 0);
    signal VN1404_in3 : std_logic_vector(1 downto 0);
    signal VN1404_in4 : std_logic_vector(1 downto 0);
    signal VN1404_in5 : std_logic_vector(1 downto 0);
    signal VN1405_in0 : std_logic_vector(1 downto 0);
    signal VN1405_in1 : std_logic_vector(1 downto 0);
    signal VN1405_in2 : std_logic_vector(1 downto 0);
    signal VN1405_in3 : std_logic_vector(1 downto 0);
    signal VN1405_in4 : std_logic_vector(1 downto 0);
    signal VN1405_in5 : std_logic_vector(1 downto 0);
    signal VN1406_in0 : std_logic_vector(1 downto 0);
    signal VN1406_in1 : std_logic_vector(1 downto 0);
    signal VN1406_in2 : std_logic_vector(1 downto 0);
    signal VN1406_in3 : std_logic_vector(1 downto 0);
    signal VN1406_in4 : std_logic_vector(1 downto 0);
    signal VN1406_in5 : std_logic_vector(1 downto 0);
    signal VN1407_in0 : std_logic_vector(1 downto 0);
    signal VN1407_in1 : std_logic_vector(1 downto 0);
    signal VN1407_in2 : std_logic_vector(1 downto 0);
    signal VN1407_in3 : std_logic_vector(1 downto 0);
    signal VN1407_in4 : std_logic_vector(1 downto 0);
    signal VN1407_in5 : std_logic_vector(1 downto 0);
    signal VN1408_in0 : std_logic_vector(1 downto 0);
    signal VN1408_in1 : std_logic_vector(1 downto 0);
    signal VN1408_in2 : std_logic_vector(1 downto 0);
    signal VN1408_in3 : std_logic_vector(1 downto 0);
    signal VN1408_in4 : std_logic_vector(1 downto 0);
    signal VN1408_in5 : std_logic_vector(1 downto 0);
    signal VN1409_in0 : std_logic_vector(1 downto 0);
    signal VN1409_in1 : std_logic_vector(1 downto 0);
    signal VN1409_in2 : std_logic_vector(1 downto 0);
    signal VN1409_in3 : std_logic_vector(1 downto 0);
    signal VN1409_in4 : std_logic_vector(1 downto 0);
    signal VN1409_in5 : std_logic_vector(1 downto 0);
    signal VN1410_in0 : std_logic_vector(1 downto 0);
    signal VN1410_in1 : std_logic_vector(1 downto 0);
    signal VN1410_in2 : std_logic_vector(1 downto 0);
    signal VN1410_in3 : std_logic_vector(1 downto 0);
    signal VN1410_in4 : std_logic_vector(1 downto 0);
    signal VN1410_in5 : std_logic_vector(1 downto 0);
    signal VN1411_in0 : std_logic_vector(1 downto 0);
    signal VN1411_in1 : std_logic_vector(1 downto 0);
    signal VN1411_in2 : std_logic_vector(1 downto 0);
    signal VN1411_in3 : std_logic_vector(1 downto 0);
    signal VN1411_in4 : std_logic_vector(1 downto 0);
    signal VN1411_in5 : std_logic_vector(1 downto 0);
    signal VN1412_in0 : std_logic_vector(1 downto 0);
    signal VN1412_in1 : std_logic_vector(1 downto 0);
    signal VN1412_in2 : std_logic_vector(1 downto 0);
    signal VN1412_in3 : std_logic_vector(1 downto 0);
    signal VN1412_in4 : std_logic_vector(1 downto 0);
    signal VN1412_in5 : std_logic_vector(1 downto 0);
    signal VN1413_in0 : std_logic_vector(1 downto 0);
    signal VN1413_in1 : std_logic_vector(1 downto 0);
    signal VN1413_in2 : std_logic_vector(1 downto 0);
    signal VN1413_in3 : std_logic_vector(1 downto 0);
    signal VN1413_in4 : std_logic_vector(1 downto 0);
    signal VN1413_in5 : std_logic_vector(1 downto 0);
    signal VN1414_in0 : std_logic_vector(1 downto 0);
    signal VN1414_in1 : std_logic_vector(1 downto 0);
    signal VN1414_in2 : std_logic_vector(1 downto 0);
    signal VN1414_in3 : std_logic_vector(1 downto 0);
    signal VN1414_in4 : std_logic_vector(1 downto 0);
    signal VN1414_in5 : std_logic_vector(1 downto 0);
    signal VN1415_in0 : std_logic_vector(1 downto 0);
    signal VN1415_in1 : std_logic_vector(1 downto 0);
    signal VN1415_in2 : std_logic_vector(1 downto 0);
    signal VN1415_in3 : std_logic_vector(1 downto 0);
    signal VN1415_in4 : std_logic_vector(1 downto 0);
    signal VN1415_in5 : std_logic_vector(1 downto 0);
    signal VN1416_in0 : std_logic_vector(1 downto 0);
    signal VN1416_in1 : std_logic_vector(1 downto 0);
    signal VN1416_in2 : std_logic_vector(1 downto 0);
    signal VN1416_in3 : std_logic_vector(1 downto 0);
    signal VN1416_in4 : std_logic_vector(1 downto 0);
    signal VN1416_in5 : std_logic_vector(1 downto 0);
    signal VN1417_in0 : std_logic_vector(1 downto 0);
    signal VN1417_in1 : std_logic_vector(1 downto 0);
    signal VN1417_in2 : std_logic_vector(1 downto 0);
    signal VN1417_in3 : std_logic_vector(1 downto 0);
    signal VN1417_in4 : std_logic_vector(1 downto 0);
    signal VN1417_in5 : std_logic_vector(1 downto 0);
    signal VN1418_in0 : std_logic_vector(1 downto 0);
    signal VN1418_in1 : std_logic_vector(1 downto 0);
    signal VN1418_in2 : std_logic_vector(1 downto 0);
    signal VN1418_in3 : std_logic_vector(1 downto 0);
    signal VN1418_in4 : std_logic_vector(1 downto 0);
    signal VN1418_in5 : std_logic_vector(1 downto 0);
    signal VN1419_in0 : std_logic_vector(1 downto 0);
    signal VN1419_in1 : std_logic_vector(1 downto 0);
    signal VN1419_in2 : std_logic_vector(1 downto 0);
    signal VN1419_in3 : std_logic_vector(1 downto 0);
    signal VN1419_in4 : std_logic_vector(1 downto 0);
    signal VN1419_in5 : std_logic_vector(1 downto 0);
    signal VN1420_in0 : std_logic_vector(1 downto 0);
    signal VN1420_in1 : std_logic_vector(1 downto 0);
    signal VN1420_in2 : std_logic_vector(1 downto 0);
    signal VN1420_in3 : std_logic_vector(1 downto 0);
    signal VN1420_in4 : std_logic_vector(1 downto 0);
    signal VN1420_in5 : std_logic_vector(1 downto 0);
    signal VN1421_in0 : std_logic_vector(1 downto 0);
    signal VN1421_in1 : std_logic_vector(1 downto 0);
    signal VN1421_in2 : std_logic_vector(1 downto 0);
    signal VN1421_in3 : std_logic_vector(1 downto 0);
    signal VN1421_in4 : std_logic_vector(1 downto 0);
    signal VN1421_in5 : std_logic_vector(1 downto 0);
    signal VN1422_in0 : std_logic_vector(1 downto 0);
    signal VN1422_in1 : std_logic_vector(1 downto 0);
    signal VN1422_in2 : std_logic_vector(1 downto 0);
    signal VN1422_in3 : std_logic_vector(1 downto 0);
    signal VN1422_in4 : std_logic_vector(1 downto 0);
    signal VN1422_in5 : std_logic_vector(1 downto 0);
    signal VN1423_in0 : std_logic_vector(1 downto 0);
    signal VN1423_in1 : std_logic_vector(1 downto 0);
    signal VN1423_in2 : std_logic_vector(1 downto 0);
    signal VN1423_in3 : std_logic_vector(1 downto 0);
    signal VN1423_in4 : std_logic_vector(1 downto 0);
    signal VN1423_in5 : std_logic_vector(1 downto 0);
    signal VN1424_in0 : std_logic_vector(1 downto 0);
    signal VN1424_in1 : std_logic_vector(1 downto 0);
    signal VN1424_in2 : std_logic_vector(1 downto 0);
    signal VN1424_in3 : std_logic_vector(1 downto 0);
    signal VN1424_in4 : std_logic_vector(1 downto 0);
    signal VN1424_in5 : std_logic_vector(1 downto 0);
    signal VN1425_in0 : std_logic_vector(1 downto 0);
    signal VN1425_in1 : std_logic_vector(1 downto 0);
    signal VN1425_in2 : std_logic_vector(1 downto 0);
    signal VN1425_in3 : std_logic_vector(1 downto 0);
    signal VN1425_in4 : std_logic_vector(1 downto 0);
    signal VN1425_in5 : std_logic_vector(1 downto 0);
    signal VN1426_in0 : std_logic_vector(1 downto 0);
    signal VN1426_in1 : std_logic_vector(1 downto 0);
    signal VN1426_in2 : std_logic_vector(1 downto 0);
    signal VN1426_in3 : std_logic_vector(1 downto 0);
    signal VN1426_in4 : std_logic_vector(1 downto 0);
    signal VN1426_in5 : std_logic_vector(1 downto 0);
    signal VN1427_in0 : std_logic_vector(1 downto 0);
    signal VN1427_in1 : std_logic_vector(1 downto 0);
    signal VN1427_in2 : std_logic_vector(1 downto 0);
    signal VN1427_in3 : std_logic_vector(1 downto 0);
    signal VN1427_in4 : std_logic_vector(1 downto 0);
    signal VN1427_in5 : std_logic_vector(1 downto 0);
    signal VN1428_in0 : std_logic_vector(1 downto 0);
    signal VN1428_in1 : std_logic_vector(1 downto 0);
    signal VN1428_in2 : std_logic_vector(1 downto 0);
    signal VN1428_in3 : std_logic_vector(1 downto 0);
    signal VN1428_in4 : std_logic_vector(1 downto 0);
    signal VN1428_in5 : std_logic_vector(1 downto 0);
    signal VN1429_in0 : std_logic_vector(1 downto 0);
    signal VN1429_in1 : std_logic_vector(1 downto 0);
    signal VN1429_in2 : std_logic_vector(1 downto 0);
    signal VN1429_in3 : std_logic_vector(1 downto 0);
    signal VN1429_in4 : std_logic_vector(1 downto 0);
    signal VN1429_in5 : std_logic_vector(1 downto 0);
    signal VN1430_in0 : std_logic_vector(1 downto 0);
    signal VN1430_in1 : std_logic_vector(1 downto 0);
    signal VN1430_in2 : std_logic_vector(1 downto 0);
    signal VN1430_in3 : std_logic_vector(1 downto 0);
    signal VN1430_in4 : std_logic_vector(1 downto 0);
    signal VN1430_in5 : std_logic_vector(1 downto 0);
    signal VN1431_in0 : std_logic_vector(1 downto 0);
    signal VN1431_in1 : std_logic_vector(1 downto 0);
    signal VN1431_in2 : std_logic_vector(1 downto 0);
    signal VN1431_in3 : std_logic_vector(1 downto 0);
    signal VN1431_in4 : std_logic_vector(1 downto 0);
    signal VN1431_in5 : std_logic_vector(1 downto 0);
    signal VN1432_in0 : std_logic_vector(1 downto 0);
    signal VN1432_in1 : std_logic_vector(1 downto 0);
    signal VN1432_in2 : std_logic_vector(1 downto 0);
    signal VN1432_in3 : std_logic_vector(1 downto 0);
    signal VN1432_in4 : std_logic_vector(1 downto 0);
    signal VN1432_in5 : std_logic_vector(1 downto 0);
    signal VN1433_in0 : std_logic_vector(1 downto 0);
    signal VN1433_in1 : std_logic_vector(1 downto 0);
    signal VN1433_in2 : std_logic_vector(1 downto 0);
    signal VN1433_in3 : std_logic_vector(1 downto 0);
    signal VN1433_in4 : std_logic_vector(1 downto 0);
    signal VN1433_in5 : std_logic_vector(1 downto 0);
    signal VN1434_in0 : std_logic_vector(1 downto 0);
    signal VN1434_in1 : std_logic_vector(1 downto 0);
    signal VN1434_in2 : std_logic_vector(1 downto 0);
    signal VN1434_in3 : std_logic_vector(1 downto 0);
    signal VN1434_in4 : std_logic_vector(1 downto 0);
    signal VN1434_in5 : std_logic_vector(1 downto 0);
    signal VN1435_in0 : std_logic_vector(1 downto 0);
    signal VN1435_in1 : std_logic_vector(1 downto 0);
    signal VN1435_in2 : std_logic_vector(1 downto 0);
    signal VN1435_in3 : std_logic_vector(1 downto 0);
    signal VN1435_in4 : std_logic_vector(1 downto 0);
    signal VN1435_in5 : std_logic_vector(1 downto 0);
    signal VN1436_in0 : std_logic_vector(1 downto 0);
    signal VN1436_in1 : std_logic_vector(1 downto 0);
    signal VN1436_in2 : std_logic_vector(1 downto 0);
    signal VN1436_in3 : std_logic_vector(1 downto 0);
    signal VN1436_in4 : std_logic_vector(1 downto 0);
    signal VN1436_in5 : std_logic_vector(1 downto 0);
    signal VN1437_in0 : std_logic_vector(1 downto 0);
    signal VN1437_in1 : std_logic_vector(1 downto 0);
    signal VN1437_in2 : std_logic_vector(1 downto 0);
    signal VN1437_in3 : std_logic_vector(1 downto 0);
    signal VN1437_in4 : std_logic_vector(1 downto 0);
    signal VN1437_in5 : std_logic_vector(1 downto 0);
    signal VN1438_in0 : std_logic_vector(1 downto 0);
    signal VN1438_in1 : std_logic_vector(1 downto 0);
    signal VN1438_in2 : std_logic_vector(1 downto 0);
    signal VN1438_in3 : std_logic_vector(1 downto 0);
    signal VN1438_in4 : std_logic_vector(1 downto 0);
    signal VN1438_in5 : std_logic_vector(1 downto 0);
    signal VN1439_in0 : std_logic_vector(1 downto 0);
    signal VN1439_in1 : std_logic_vector(1 downto 0);
    signal VN1439_in2 : std_logic_vector(1 downto 0);
    signal VN1439_in3 : std_logic_vector(1 downto 0);
    signal VN1439_in4 : std_logic_vector(1 downto 0);
    signal VN1439_in5 : std_logic_vector(1 downto 0);
    signal VN1440_in0 : std_logic_vector(1 downto 0);
    signal VN1440_in1 : std_logic_vector(1 downto 0);
    signal VN1440_in2 : std_logic_vector(1 downto 0);
    signal VN1440_in3 : std_logic_vector(1 downto 0);
    signal VN1440_in4 : std_logic_vector(1 downto 0);
    signal VN1440_in5 : std_logic_vector(1 downto 0);
    signal VN1441_in0 : std_logic_vector(1 downto 0);
    signal VN1441_in1 : std_logic_vector(1 downto 0);
    signal VN1441_in2 : std_logic_vector(1 downto 0);
    signal VN1441_in3 : std_logic_vector(1 downto 0);
    signal VN1441_in4 : std_logic_vector(1 downto 0);
    signal VN1441_in5 : std_logic_vector(1 downto 0);
    signal VN1442_in0 : std_logic_vector(1 downto 0);
    signal VN1442_in1 : std_logic_vector(1 downto 0);
    signal VN1442_in2 : std_logic_vector(1 downto 0);
    signal VN1442_in3 : std_logic_vector(1 downto 0);
    signal VN1442_in4 : std_logic_vector(1 downto 0);
    signal VN1442_in5 : std_logic_vector(1 downto 0);
    signal VN1443_in0 : std_logic_vector(1 downto 0);
    signal VN1443_in1 : std_logic_vector(1 downto 0);
    signal VN1443_in2 : std_logic_vector(1 downto 0);
    signal VN1443_in3 : std_logic_vector(1 downto 0);
    signal VN1443_in4 : std_logic_vector(1 downto 0);
    signal VN1443_in5 : std_logic_vector(1 downto 0);
    signal VN1444_in0 : std_logic_vector(1 downto 0);
    signal VN1444_in1 : std_logic_vector(1 downto 0);
    signal VN1444_in2 : std_logic_vector(1 downto 0);
    signal VN1444_in3 : std_logic_vector(1 downto 0);
    signal VN1444_in4 : std_logic_vector(1 downto 0);
    signal VN1444_in5 : std_logic_vector(1 downto 0);
    signal VN1445_in0 : std_logic_vector(1 downto 0);
    signal VN1445_in1 : std_logic_vector(1 downto 0);
    signal VN1445_in2 : std_logic_vector(1 downto 0);
    signal VN1445_in3 : std_logic_vector(1 downto 0);
    signal VN1445_in4 : std_logic_vector(1 downto 0);
    signal VN1445_in5 : std_logic_vector(1 downto 0);
    signal VN1446_in0 : std_logic_vector(1 downto 0);
    signal VN1446_in1 : std_logic_vector(1 downto 0);
    signal VN1446_in2 : std_logic_vector(1 downto 0);
    signal VN1446_in3 : std_logic_vector(1 downto 0);
    signal VN1446_in4 : std_logic_vector(1 downto 0);
    signal VN1446_in5 : std_logic_vector(1 downto 0);
    signal VN1447_in0 : std_logic_vector(1 downto 0);
    signal VN1447_in1 : std_logic_vector(1 downto 0);
    signal VN1447_in2 : std_logic_vector(1 downto 0);
    signal VN1447_in3 : std_logic_vector(1 downto 0);
    signal VN1447_in4 : std_logic_vector(1 downto 0);
    signal VN1447_in5 : std_logic_vector(1 downto 0);
    signal VN1448_in0 : std_logic_vector(1 downto 0);
    signal VN1448_in1 : std_logic_vector(1 downto 0);
    signal VN1448_in2 : std_logic_vector(1 downto 0);
    signal VN1448_in3 : std_logic_vector(1 downto 0);
    signal VN1448_in4 : std_logic_vector(1 downto 0);
    signal VN1448_in5 : std_logic_vector(1 downto 0);
    signal VN1449_in0 : std_logic_vector(1 downto 0);
    signal VN1449_in1 : std_logic_vector(1 downto 0);
    signal VN1449_in2 : std_logic_vector(1 downto 0);
    signal VN1449_in3 : std_logic_vector(1 downto 0);
    signal VN1449_in4 : std_logic_vector(1 downto 0);
    signal VN1449_in5 : std_logic_vector(1 downto 0);
    signal VN1450_in0 : std_logic_vector(1 downto 0);
    signal VN1450_in1 : std_logic_vector(1 downto 0);
    signal VN1450_in2 : std_logic_vector(1 downto 0);
    signal VN1450_in3 : std_logic_vector(1 downto 0);
    signal VN1450_in4 : std_logic_vector(1 downto 0);
    signal VN1450_in5 : std_logic_vector(1 downto 0);
    signal VN1451_in0 : std_logic_vector(1 downto 0);
    signal VN1451_in1 : std_logic_vector(1 downto 0);
    signal VN1451_in2 : std_logic_vector(1 downto 0);
    signal VN1451_in3 : std_logic_vector(1 downto 0);
    signal VN1451_in4 : std_logic_vector(1 downto 0);
    signal VN1451_in5 : std_logic_vector(1 downto 0);
    signal VN1452_in0 : std_logic_vector(1 downto 0);
    signal VN1452_in1 : std_logic_vector(1 downto 0);
    signal VN1452_in2 : std_logic_vector(1 downto 0);
    signal VN1452_in3 : std_logic_vector(1 downto 0);
    signal VN1452_in4 : std_logic_vector(1 downto 0);
    signal VN1452_in5 : std_logic_vector(1 downto 0);
    signal VN1453_in0 : std_logic_vector(1 downto 0);
    signal VN1453_in1 : std_logic_vector(1 downto 0);
    signal VN1453_in2 : std_logic_vector(1 downto 0);
    signal VN1453_in3 : std_logic_vector(1 downto 0);
    signal VN1453_in4 : std_logic_vector(1 downto 0);
    signal VN1453_in5 : std_logic_vector(1 downto 0);
    signal VN1454_in0 : std_logic_vector(1 downto 0);
    signal VN1454_in1 : std_logic_vector(1 downto 0);
    signal VN1454_in2 : std_logic_vector(1 downto 0);
    signal VN1454_in3 : std_logic_vector(1 downto 0);
    signal VN1454_in4 : std_logic_vector(1 downto 0);
    signal VN1454_in5 : std_logic_vector(1 downto 0);
    signal VN1455_in0 : std_logic_vector(1 downto 0);
    signal VN1455_in1 : std_logic_vector(1 downto 0);
    signal VN1455_in2 : std_logic_vector(1 downto 0);
    signal VN1455_in3 : std_logic_vector(1 downto 0);
    signal VN1455_in4 : std_logic_vector(1 downto 0);
    signal VN1455_in5 : std_logic_vector(1 downto 0);
    signal VN1456_in0 : std_logic_vector(1 downto 0);
    signal VN1456_in1 : std_logic_vector(1 downto 0);
    signal VN1456_in2 : std_logic_vector(1 downto 0);
    signal VN1456_in3 : std_logic_vector(1 downto 0);
    signal VN1456_in4 : std_logic_vector(1 downto 0);
    signal VN1456_in5 : std_logic_vector(1 downto 0);
    signal VN1457_in0 : std_logic_vector(1 downto 0);
    signal VN1457_in1 : std_logic_vector(1 downto 0);
    signal VN1457_in2 : std_logic_vector(1 downto 0);
    signal VN1457_in3 : std_logic_vector(1 downto 0);
    signal VN1457_in4 : std_logic_vector(1 downto 0);
    signal VN1457_in5 : std_logic_vector(1 downto 0);
    signal VN1458_in0 : std_logic_vector(1 downto 0);
    signal VN1458_in1 : std_logic_vector(1 downto 0);
    signal VN1458_in2 : std_logic_vector(1 downto 0);
    signal VN1458_in3 : std_logic_vector(1 downto 0);
    signal VN1458_in4 : std_logic_vector(1 downto 0);
    signal VN1458_in5 : std_logic_vector(1 downto 0);
    signal VN1459_in0 : std_logic_vector(1 downto 0);
    signal VN1459_in1 : std_logic_vector(1 downto 0);
    signal VN1459_in2 : std_logic_vector(1 downto 0);
    signal VN1459_in3 : std_logic_vector(1 downto 0);
    signal VN1459_in4 : std_logic_vector(1 downto 0);
    signal VN1459_in5 : std_logic_vector(1 downto 0);
    signal VN1460_in0 : std_logic_vector(1 downto 0);
    signal VN1460_in1 : std_logic_vector(1 downto 0);
    signal VN1460_in2 : std_logic_vector(1 downto 0);
    signal VN1460_in3 : std_logic_vector(1 downto 0);
    signal VN1460_in4 : std_logic_vector(1 downto 0);
    signal VN1460_in5 : std_logic_vector(1 downto 0);
    signal VN1461_in0 : std_logic_vector(1 downto 0);
    signal VN1461_in1 : std_logic_vector(1 downto 0);
    signal VN1461_in2 : std_logic_vector(1 downto 0);
    signal VN1461_in3 : std_logic_vector(1 downto 0);
    signal VN1461_in4 : std_logic_vector(1 downto 0);
    signal VN1461_in5 : std_logic_vector(1 downto 0);
    signal VN1462_in0 : std_logic_vector(1 downto 0);
    signal VN1462_in1 : std_logic_vector(1 downto 0);
    signal VN1462_in2 : std_logic_vector(1 downto 0);
    signal VN1462_in3 : std_logic_vector(1 downto 0);
    signal VN1462_in4 : std_logic_vector(1 downto 0);
    signal VN1462_in5 : std_logic_vector(1 downto 0);
    signal VN1463_in0 : std_logic_vector(1 downto 0);
    signal VN1463_in1 : std_logic_vector(1 downto 0);
    signal VN1463_in2 : std_logic_vector(1 downto 0);
    signal VN1463_in3 : std_logic_vector(1 downto 0);
    signal VN1463_in4 : std_logic_vector(1 downto 0);
    signal VN1463_in5 : std_logic_vector(1 downto 0);
    signal VN1464_in0 : std_logic_vector(1 downto 0);
    signal VN1464_in1 : std_logic_vector(1 downto 0);
    signal VN1464_in2 : std_logic_vector(1 downto 0);
    signal VN1464_in3 : std_logic_vector(1 downto 0);
    signal VN1464_in4 : std_logic_vector(1 downto 0);
    signal VN1464_in5 : std_logic_vector(1 downto 0);
    signal VN1465_in0 : std_logic_vector(1 downto 0);
    signal VN1465_in1 : std_logic_vector(1 downto 0);
    signal VN1465_in2 : std_logic_vector(1 downto 0);
    signal VN1465_in3 : std_logic_vector(1 downto 0);
    signal VN1465_in4 : std_logic_vector(1 downto 0);
    signal VN1465_in5 : std_logic_vector(1 downto 0);
    signal VN1466_in0 : std_logic_vector(1 downto 0);
    signal VN1466_in1 : std_logic_vector(1 downto 0);
    signal VN1466_in2 : std_logic_vector(1 downto 0);
    signal VN1466_in3 : std_logic_vector(1 downto 0);
    signal VN1466_in4 : std_logic_vector(1 downto 0);
    signal VN1466_in5 : std_logic_vector(1 downto 0);
    signal VN1467_in0 : std_logic_vector(1 downto 0);
    signal VN1467_in1 : std_logic_vector(1 downto 0);
    signal VN1467_in2 : std_logic_vector(1 downto 0);
    signal VN1467_in3 : std_logic_vector(1 downto 0);
    signal VN1467_in4 : std_logic_vector(1 downto 0);
    signal VN1467_in5 : std_logic_vector(1 downto 0);
    signal VN1468_in0 : std_logic_vector(1 downto 0);
    signal VN1468_in1 : std_logic_vector(1 downto 0);
    signal VN1468_in2 : std_logic_vector(1 downto 0);
    signal VN1468_in3 : std_logic_vector(1 downto 0);
    signal VN1468_in4 : std_logic_vector(1 downto 0);
    signal VN1468_in5 : std_logic_vector(1 downto 0);
    signal VN1469_in0 : std_logic_vector(1 downto 0);
    signal VN1469_in1 : std_logic_vector(1 downto 0);
    signal VN1469_in2 : std_logic_vector(1 downto 0);
    signal VN1469_in3 : std_logic_vector(1 downto 0);
    signal VN1469_in4 : std_logic_vector(1 downto 0);
    signal VN1469_in5 : std_logic_vector(1 downto 0);
    signal VN1470_in0 : std_logic_vector(1 downto 0);
    signal VN1470_in1 : std_logic_vector(1 downto 0);
    signal VN1470_in2 : std_logic_vector(1 downto 0);
    signal VN1470_in3 : std_logic_vector(1 downto 0);
    signal VN1470_in4 : std_logic_vector(1 downto 0);
    signal VN1470_in5 : std_logic_vector(1 downto 0);
    signal VN1471_in0 : std_logic_vector(1 downto 0);
    signal VN1471_in1 : std_logic_vector(1 downto 0);
    signal VN1471_in2 : std_logic_vector(1 downto 0);
    signal VN1471_in3 : std_logic_vector(1 downto 0);
    signal VN1471_in4 : std_logic_vector(1 downto 0);
    signal VN1471_in5 : std_logic_vector(1 downto 0);
    signal VN1472_in0 : std_logic_vector(1 downto 0);
    signal VN1472_in1 : std_logic_vector(1 downto 0);
    signal VN1472_in2 : std_logic_vector(1 downto 0);
    signal VN1472_in3 : std_logic_vector(1 downto 0);
    signal VN1472_in4 : std_logic_vector(1 downto 0);
    signal VN1472_in5 : std_logic_vector(1 downto 0);
    signal VN1473_in0 : std_logic_vector(1 downto 0);
    signal VN1473_in1 : std_logic_vector(1 downto 0);
    signal VN1473_in2 : std_logic_vector(1 downto 0);
    signal VN1473_in3 : std_logic_vector(1 downto 0);
    signal VN1473_in4 : std_logic_vector(1 downto 0);
    signal VN1473_in5 : std_logic_vector(1 downto 0);
    signal VN1474_in0 : std_logic_vector(1 downto 0);
    signal VN1474_in1 : std_logic_vector(1 downto 0);
    signal VN1474_in2 : std_logic_vector(1 downto 0);
    signal VN1474_in3 : std_logic_vector(1 downto 0);
    signal VN1474_in4 : std_logic_vector(1 downto 0);
    signal VN1474_in5 : std_logic_vector(1 downto 0);
    signal VN1475_in0 : std_logic_vector(1 downto 0);
    signal VN1475_in1 : std_logic_vector(1 downto 0);
    signal VN1475_in2 : std_logic_vector(1 downto 0);
    signal VN1475_in3 : std_logic_vector(1 downto 0);
    signal VN1475_in4 : std_logic_vector(1 downto 0);
    signal VN1475_in5 : std_logic_vector(1 downto 0);
    signal VN1476_in0 : std_logic_vector(1 downto 0);
    signal VN1476_in1 : std_logic_vector(1 downto 0);
    signal VN1476_in2 : std_logic_vector(1 downto 0);
    signal VN1476_in3 : std_logic_vector(1 downto 0);
    signal VN1476_in4 : std_logic_vector(1 downto 0);
    signal VN1476_in5 : std_logic_vector(1 downto 0);
    signal VN1477_in0 : std_logic_vector(1 downto 0);
    signal VN1477_in1 : std_logic_vector(1 downto 0);
    signal VN1477_in2 : std_logic_vector(1 downto 0);
    signal VN1477_in3 : std_logic_vector(1 downto 0);
    signal VN1477_in4 : std_logic_vector(1 downto 0);
    signal VN1477_in5 : std_logic_vector(1 downto 0);
    signal VN1478_in0 : std_logic_vector(1 downto 0);
    signal VN1478_in1 : std_logic_vector(1 downto 0);
    signal VN1478_in2 : std_logic_vector(1 downto 0);
    signal VN1478_in3 : std_logic_vector(1 downto 0);
    signal VN1478_in4 : std_logic_vector(1 downto 0);
    signal VN1478_in5 : std_logic_vector(1 downto 0);
    signal VN1479_in0 : std_logic_vector(1 downto 0);
    signal VN1479_in1 : std_logic_vector(1 downto 0);
    signal VN1479_in2 : std_logic_vector(1 downto 0);
    signal VN1479_in3 : std_logic_vector(1 downto 0);
    signal VN1479_in4 : std_logic_vector(1 downto 0);
    signal VN1479_in5 : std_logic_vector(1 downto 0);
    signal VN1480_in0 : std_logic_vector(1 downto 0);
    signal VN1480_in1 : std_logic_vector(1 downto 0);
    signal VN1480_in2 : std_logic_vector(1 downto 0);
    signal VN1480_in3 : std_logic_vector(1 downto 0);
    signal VN1480_in4 : std_logic_vector(1 downto 0);
    signal VN1480_in5 : std_logic_vector(1 downto 0);
    signal VN1481_in0 : std_logic_vector(1 downto 0);
    signal VN1481_in1 : std_logic_vector(1 downto 0);
    signal VN1481_in2 : std_logic_vector(1 downto 0);
    signal VN1481_in3 : std_logic_vector(1 downto 0);
    signal VN1481_in4 : std_logic_vector(1 downto 0);
    signal VN1481_in5 : std_logic_vector(1 downto 0);
    signal VN1482_in0 : std_logic_vector(1 downto 0);
    signal VN1482_in1 : std_logic_vector(1 downto 0);
    signal VN1482_in2 : std_logic_vector(1 downto 0);
    signal VN1482_in3 : std_logic_vector(1 downto 0);
    signal VN1482_in4 : std_logic_vector(1 downto 0);
    signal VN1482_in5 : std_logic_vector(1 downto 0);
    signal VN1483_in0 : std_logic_vector(1 downto 0);
    signal VN1483_in1 : std_logic_vector(1 downto 0);
    signal VN1483_in2 : std_logic_vector(1 downto 0);
    signal VN1483_in3 : std_logic_vector(1 downto 0);
    signal VN1483_in4 : std_logic_vector(1 downto 0);
    signal VN1483_in5 : std_logic_vector(1 downto 0);
    signal VN1484_in0 : std_logic_vector(1 downto 0);
    signal VN1484_in1 : std_logic_vector(1 downto 0);
    signal VN1484_in2 : std_logic_vector(1 downto 0);
    signal VN1484_in3 : std_logic_vector(1 downto 0);
    signal VN1484_in4 : std_logic_vector(1 downto 0);
    signal VN1484_in5 : std_logic_vector(1 downto 0);
    signal VN1485_in0 : std_logic_vector(1 downto 0);
    signal VN1485_in1 : std_logic_vector(1 downto 0);
    signal VN1485_in2 : std_logic_vector(1 downto 0);
    signal VN1485_in3 : std_logic_vector(1 downto 0);
    signal VN1485_in4 : std_logic_vector(1 downto 0);
    signal VN1485_in5 : std_logic_vector(1 downto 0);
    signal VN1486_in0 : std_logic_vector(1 downto 0);
    signal VN1486_in1 : std_logic_vector(1 downto 0);
    signal VN1486_in2 : std_logic_vector(1 downto 0);
    signal VN1486_in3 : std_logic_vector(1 downto 0);
    signal VN1486_in4 : std_logic_vector(1 downto 0);
    signal VN1486_in5 : std_logic_vector(1 downto 0);
    signal VN1487_in0 : std_logic_vector(1 downto 0);
    signal VN1487_in1 : std_logic_vector(1 downto 0);
    signal VN1487_in2 : std_logic_vector(1 downto 0);
    signal VN1487_in3 : std_logic_vector(1 downto 0);
    signal VN1487_in4 : std_logic_vector(1 downto 0);
    signal VN1487_in5 : std_logic_vector(1 downto 0);
    signal VN1488_in0 : std_logic_vector(1 downto 0);
    signal VN1488_in1 : std_logic_vector(1 downto 0);
    signal VN1488_in2 : std_logic_vector(1 downto 0);
    signal VN1488_in3 : std_logic_vector(1 downto 0);
    signal VN1488_in4 : std_logic_vector(1 downto 0);
    signal VN1488_in5 : std_logic_vector(1 downto 0);
    signal VN1489_in0 : std_logic_vector(1 downto 0);
    signal VN1489_in1 : std_logic_vector(1 downto 0);
    signal VN1489_in2 : std_logic_vector(1 downto 0);
    signal VN1489_in3 : std_logic_vector(1 downto 0);
    signal VN1489_in4 : std_logic_vector(1 downto 0);
    signal VN1489_in5 : std_logic_vector(1 downto 0);
    signal VN1490_in0 : std_logic_vector(1 downto 0);
    signal VN1490_in1 : std_logic_vector(1 downto 0);
    signal VN1490_in2 : std_logic_vector(1 downto 0);
    signal VN1490_in3 : std_logic_vector(1 downto 0);
    signal VN1490_in4 : std_logic_vector(1 downto 0);
    signal VN1490_in5 : std_logic_vector(1 downto 0);
    signal VN1491_in0 : std_logic_vector(1 downto 0);
    signal VN1491_in1 : std_logic_vector(1 downto 0);
    signal VN1491_in2 : std_logic_vector(1 downto 0);
    signal VN1491_in3 : std_logic_vector(1 downto 0);
    signal VN1491_in4 : std_logic_vector(1 downto 0);
    signal VN1491_in5 : std_logic_vector(1 downto 0);
    signal VN1492_in0 : std_logic_vector(1 downto 0);
    signal VN1492_in1 : std_logic_vector(1 downto 0);
    signal VN1492_in2 : std_logic_vector(1 downto 0);
    signal VN1492_in3 : std_logic_vector(1 downto 0);
    signal VN1492_in4 : std_logic_vector(1 downto 0);
    signal VN1492_in5 : std_logic_vector(1 downto 0);
    signal VN1493_in0 : std_logic_vector(1 downto 0);
    signal VN1493_in1 : std_logic_vector(1 downto 0);
    signal VN1493_in2 : std_logic_vector(1 downto 0);
    signal VN1493_in3 : std_logic_vector(1 downto 0);
    signal VN1493_in4 : std_logic_vector(1 downto 0);
    signal VN1493_in5 : std_logic_vector(1 downto 0);
    signal VN1494_in0 : std_logic_vector(1 downto 0);
    signal VN1494_in1 : std_logic_vector(1 downto 0);
    signal VN1494_in2 : std_logic_vector(1 downto 0);
    signal VN1494_in3 : std_logic_vector(1 downto 0);
    signal VN1494_in4 : std_logic_vector(1 downto 0);
    signal VN1494_in5 : std_logic_vector(1 downto 0);
    signal VN1495_in0 : std_logic_vector(1 downto 0);
    signal VN1495_in1 : std_logic_vector(1 downto 0);
    signal VN1495_in2 : std_logic_vector(1 downto 0);
    signal VN1495_in3 : std_logic_vector(1 downto 0);
    signal VN1495_in4 : std_logic_vector(1 downto 0);
    signal VN1495_in5 : std_logic_vector(1 downto 0);
    signal VN1496_in0 : std_logic_vector(1 downto 0);
    signal VN1496_in1 : std_logic_vector(1 downto 0);
    signal VN1496_in2 : std_logic_vector(1 downto 0);
    signal VN1496_in3 : std_logic_vector(1 downto 0);
    signal VN1496_in4 : std_logic_vector(1 downto 0);
    signal VN1496_in5 : std_logic_vector(1 downto 0);
    signal VN1497_in0 : std_logic_vector(1 downto 0);
    signal VN1497_in1 : std_logic_vector(1 downto 0);
    signal VN1497_in2 : std_logic_vector(1 downto 0);
    signal VN1497_in3 : std_logic_vector(1 downto 0);
    signal VN1497_in4 : std_logic_vector(1 downto 0);
    signal VN1497_in5 : std_logic_vector(1 downto 0);
    signal VN1498_in0 : std_logic_vector(1 downto 0);
    signal VN1498_in1 : std_logic_vector(1 downto 0);
    signal VN1498_in2 : std_logic_vector(1 downto 0);
    signal VN1498_in3 : std_logic_vector(1 downto 0);
    signal VN1498_in4 : std_logic_vector(1 downto 0);
    signal VN1498_in5 : std_logic_vector(1 downto 0);
    signal VN1499_in0 : std_logic_vector(1 downto 0);
    signal VN1499_in1 : std_logic_vector(1 downto 0);
    signal VN1499_in2 : std_logic_vector(1 downto 0);
    signal VN1499_in3 : std_logic_vector(1 downto 0);
    signal VN1499_in4 : std_logic_vector(1 downto 0);
    signal VN1499_in5 : std_logic_vector(1 downto 0);
    signal VN1500_in0 : std_logic_vector(1 downto 0);
    signal VN1500_in1 : std_logic_vector(1 downto 0);
    signal VN1500_in2 : std_logic_vector(1 downto 0);
    signal VN1500_in3 : std_logic_vector(1 downto 0);
    signal VN1500_in4 : std_logic_vector(1 downto 0);
    signal VN1500_in5 : std_logic_vector(1 downto 0);
    signal VN1501_in0 : std_logic_vector(1 downto 0);
    signal VN1501_in1 : std_logic_vector(1 downto 0);
    signal VN1501_in2 : std_logic_vector(1 downto 0);
    signal VN1501_in3 : std_logic_vector(1 downto 0);
    signal VN1501_in4 : std_logic_vector(1 downto 0);
    signal VN1501_in5 : std_logic_vector(1 downto 0);
    signal VN1502_in0 : std_logic_vector(1 downto 0);
    signal VN1502_in1 : std_logic_vector(1 downto 0);
    signal VN1502_in2 : std_logic_vector(1 downto 0);
    signal VN1502_in3 : std_logic_vector(1 downto 0);
    signal VN1502_in4 : std_logic_vector(1 downto 0);
    signal VN1502_in5 : std_logic_vector(1 downto 0);
    signal VN1503_in0 : std_logic_vector(1 downto 0);
    signal VN1503_in1 : std_logic_vector(1 downto 0);
    signal VN1503_in2 : std_logic_vector(1 downto 0);
    signal VN1503_in3 : std_logic_vector(1 downto 0);
    signal VN1503_in4 : std_logic_vector(1 downto 0);
    signal VN1503_in5 : std_logic_vector(1 downto 0);
    signal VN1504_in0 : std_logic_vector(1 downto 0);
    signal VN1504_in1 : std_logic_vector(1 downto 0);
    signal VN1504_in2 : std_logic_vector(1 downto 0);
    signal VN1504_in3 : std_logic_vector(1 downto 0);
    signal VN1504_in4 : std_logic_vector(1 downto 0);
    signal VN1504_in5 : std_logic_vector(1 downto 0);
    signal VN1505_in0 : std_logic_vector(1 downto 0);
    signal VN1505_in1 : std_logic_vector(1 downto 0);
    signal VN1505_in2 : std_logic_vector(1 downto 0);
    signal VN1505_in3 : std_logic_vector(1 downto 0);
    signal VN1505_in4 : std_logic_vector(1 downto 0);
    signal VN1505_in5 : std_logic_vector(1 downto 0);
    signal VN1506_in0 : std_logic_vector(1 downto 0);
    signal VN1506_in1 : std_logic_vector(1 downto 0);
    signal VN1506_in2 : std_logic_vector(1 downto 0);
    signal VN1506_in3 : std_logic_vector(1 downto 0);
    signal VN1506_in4 : std_logic_vector(1 downto 0);
    signal VN1506_in5 : std_logic_vector(1 downto 0);
    signal VN1507_in0 : std_logic_vector(1 downto 0);
    signal VN1507_in1 : std_logic_vector(1 downto 0);
    signal VN1507_in2 : std_logic_vector(1 downto 0);
    signal VN1507_in3 : std_logic_vector(1 downto 0);
    signal VN1507_in4 : std_logic_vector(1 downto 0);
    signal VN1507_in5 : std_logic_vector(1 downto 0);
    signal VN1508_in0 : std_logic_vector(1 downto 0);
    signal VN1508_in1 : std_logic_vector(1 downto 0);
    signal VN1508_in2 : std_logic_vector(1 downto 0);
    signal VN1508_in3 : std_logic_vector(1 downto 0);
    signal VN1508_in4 : std_logic_vector(1 downto 0);
    signal VN1508_in5 : std_logic_vector(1 downto 0);
    signal VN1509_in0 : std_logic_vector(1 downto 0);
    signal VN1509_in1 : std_logic_vector(1 downto 0);
    signal VN1509_in2 : std_logic_vector(1 downto 0);
    signal VN1509_in3 : std_logic_vector(1 downto 0);
    signal VN1509_in4 : std_logic_vector(1 downto 0);
    signal VN1509_in5 : std_logic_vector(1 downto 0);
    signal VN1510_in0 : std_logic_vector(1 downto 0);
    signal VN1510_in1 : std_logic_vector(1 downto 0);
    signal VN1510_in2 : std_logic_vector(1 downto 0);
    signal VN1510_in3 : std_logic_vector(1 downto 0);
    signal VN1510_in4 : std_logic_vector(1 downto 0);
    signal VN1510_in5 : std_logic_vector(1 downto 0);
    signal VN1511_in0 : std_logic_vector(1 downto 0);
    signal VN1511_in1 : std_logic_vector(1 downto 0);
    signal VN1511_in2 : std_logic_vector(1 downto 0);
    signal VN1511_in3 : std_logic_vector(1 downto 0);
    signal VN1511_in4 : std_logic_vector(1 downto 0);
    signal VN1511_in5 : std_logic_vector(1 downto 0);
    signal VN1512_in0 : std_logic_vector(1 downto 0);
    signal VN1512_in1 : std_logic_vector(1 downto 0);
    signal VN1512_in2 : std_logic_vector(1 downto 0);
    signal VN1512_in3 : std_logic_vector(1 downto 0);
    signal VN1512_in4 : std_logic_vector(1 downto 0);
    signal VN1512_in5 : std_logic_vector(1 downto 0);
    signal VN1513_in0 : std_logic_vector(1 downto 0);
    signal VN1513_in1 : std_logic_vector(1 downto 0);
    signal VN1513_in2 : std_logic_vector(1 downto 0);
    signal VN1513_in3 : std_logic_vector(1 downto 0);
    signal VN1513_in4 : std_logic_vector(1 downto 0);
    signal VN1513_in5 : std_logic_vector(1 downto 0);
    signal VN1514_in0 : std_logic_vector(1 downto 0);
    signal VN1514_in1 : std_logic_vector(1 downto 0);
    signal VN1514_in2 : std_logic_vector(1 downto 0);
    signal VN1514_in3 : std_logic_vector(1 downto 0);
    signal VN1514_in4 : std_logic_vector(1 downto 0);
    signal VN1514_in5 : std_logic_vector(1 downto 0);
    signal VN1515_in0 : std_logic_vector(1 downto 0);
    signal VN1515_in1 : std_logic_vector(1 downto 0);
    signal VN1515_in2 : std_logic_vector(1 downto 0);
    signal VN1515_in3 : std_logic_vector(1 downto 0);
    signal VN1515_in4 : std_logic_vector(1 downto 0);
    signal VN1515_in5 : std_logic_vector(1 downto 0);
    signal VN1516_in0 : std_logic_vector(1 downto 0);
    signal VN1516_in1 : std_logic_vector(1 downto 0);
    signal VN1516_in2 : std_logic_vector(1 downto 0);
    signal VN1516_in3 : std_logic_vector(1 downto 0);
    signal VN1516_in4 : std_logic_vector(1 downto 0);
    signal VN1516_in5 : std_logic_vector(1 downto 0);
    signal VN1517_in0 : std_logic_vector(1 downto 0);
    signal VN1517_in1 : std_logic_vector(1 downto 0);
    signal VN1517_in2 : std_logic_vector(1 downto 0);
    signal VN1517_in3 : std_logic_vector(1 downto 0);
    signal VN1517_in4 : std_logic_vector(1 downto 0);
    signal VN1517_in5 : std_logic_vector(1 downto 0);
    signal VN1518_in0 : std_logic_vector(1 downto 0);
    signal VN1518_in1 : std_logic_vector(1 downto 0);
    signal VN1518_in2 : std_logic_vector(1 downto 0);
    signal VN1518_in3 : std_logic_vector(1 downto 0);
    signal VN1518_in4 : std_logic_vector(1 downto 0);
    signal VN1518_in5 : std_logic_vector(1 downto 0);
    signal VN1519_in0 : std_logic_vector(1 downto 0);
    signal VN1519_in1 : std_logic_vector(1 downto 0);
    signal VN1519_in2 : std_logic_vector(1 downto 0);
    signal VN1519_in3 : std_logic_vector(1 downto 0);
    signal VN1519_in4 : std_logic_vector(1 downto 0);
    signal VN1519_in5 : std_logic_vector(1 downto 0);
    signal VN1520_in0 : std_logic_vector(1 downto 0);
    signal VN1520_in1 : std_logic_vector(1 downto 0);
    signal VN1520_in2 : std_logic_vector(1 downto 0);
    signal VN1520_in3 : std_logic_vector(1 downto 0);
    signal VN1520_in4 : std_logic_vector(1 downto 0);
    signal VN1520_in5 : std_logic_vector(1 downto 0);
    signal VN1521_in0 : std_logic_vector(1 downto 0);
    signal VN1521_in1 : std_logic_vector(1 downto 0);
    signal VN1521_in2 : std_logic_vector(1 downto 0);
    signal VN1521_in3 : std_logic_vector(1 downto 0);
    signal VN1521_in4 : std_logic_vector(1 downto 0);
    signal VN1521_in5 : std_logic_vector(1 downto 0);
    signal VN1522_in0 : std_logic_vector(1 downto 0);
    signal VN1522_in1 : std_logic_vector(1 downto 0);
    signal VN1522_in2 : std_logic_vector(1 downto 0);
    signal VN1522_in3 : std_logic_vector(1 downto 0);
    signal VN1522_in4 : std_logic_vector(1 downto 0);
    signal VN1522_in5 : std_logic_vector(1 downto 0);
    signal VN1523_in0 : std_logic_vector(1 downto 0);
    signal VN1523_in1 : std_logic_vector(1 downto 0);
    signal VN1523_in2 : std_logic_vector(1 downto 0);
    signal VN1523_in3 : std_logic_vector(1 downto 0);
    signal VN1523_in4 : std_logic_vector(1 downto 0);
    signal VN1523_in5 : std_logic_vector(1 downto 0);
    signal VN1524_in0 : std_logic_vector(1 downto 0);
    signal VN1524_in1 : std_logic_vector(1 downto 0);
    signal VN1524_in2 : std_logic_vector(1 downto 0);
    signal VN1524_in3 : std_logic_vector(1 downto 0);
    signal VN1524_in4 : std_logic_vector(1 downto 0);
    signal VN1524_in5 : std_logic_vector(1 downto 0);
    signal VN1525_in0 : std_logic_vector(1 downto 0);
    signal VN1525_in1 : std_logic_vector(1 downto 0);
    signal VN1525_in2 : std_logic_vector(1 downto 0);
    signal VN1525_in3 : std_logic_vector(1 downto 0);
    signal VN1525_in4 : std_logic_vector(1 downto 0);
    signal VN1525_in5 : std_logic_vector(1 downto 0);
    signal VN1526_in0 : std_logic_vector(1 downto 0);
    signal VN1526_in1 : std_logic_vector(1 downto 0);
    signal VN1526_in2 : std_logic_vector(1 downto 0);
    signal VN1526_in3 : std_logic_vector(1 downto 0);
    signal VN1526_in4 : std_logic_vector(1 downto 0);
    signal VN1526_in5 : std_logic_vector(1 downto 0);
    signal VN1527_in0 : std_logic_vector(1 downto 0);
    signal VN1527_in1 : std_logic_vector(1 downto 0);
    signal VN1527_in2 : std_logic_vector(1 downto 0);
    signal VN1527_in3 : std_logic_vector(1 downto 0);
    signal VN1527_in4 : std_logic_vector(1 downto 0);
    signal VN1527_in5 : std_logic_vector(1 downto 0);
    signal VN1528_in0 : std_logic_vector(1 downto 0);
    signal VN1528_in1 : std_logic_vector(1 downto 0);
    signal VN1528_in2 : std_logic_vector(1 downto 0);
    signal VN1528_in3 : std_logic_vector(1 downto 0);
    signal VN1528_in4 : std_logic_vector(1 downto 0);
    signal VN1528_in5 : std_logic_vector(1 downto 0);
    signal VN1529_in0 : std_logic_vector(1 downto 0);
    signal VN1529_in1 : std_logic_vector(1 downto 0);
    signal VN1529_in2 : std_logic_vector(1 downto 0);
    signal VN1529_in3 : std_logic_vector(1 downto 0);
    signal VN1529_in4 : std_logic_vector(1 downto 0);
    signal VN1529_in5 : std_logic_vector(1 downto 0);
    signal VN1530_in0 : std_logic_vector(1 downto 0);
    signal VN1530_in1 : std_logic_vector(1 downto 0);
    signal VN1530_in2 : std_logic_vector(1 downto 0);
    signal VN1530_in3 : std_logic_vector(1 downto 0);
    signal VN1530_in4 : std_logic_vector(1 downto 0);
    signal VN1530_in5 : std_logic_vector(1 downto 0);
    signal VN1531_in0 : std_logic_vector(1 downto 0);
    signal VN1531_in1 : std_logic_vector(1 downto 0);
    signal VN1531_in2 : std_logic_vector(1 downto 0);
    signal VN1531_in3 : std_logic_vector(1 downto 0);
    signal VN1531_in4 : std_logic_vector(1 downto 0);
    signal VN1531_in5 : std_logic_vector(1 downto 0);
    signal VN1532_in0 : std_logic_vector(1 downto 0);
    signal VN1532_in1 : std_logic_vector(1 downto 0);
    signal VN1532_in2 : std_logic_vector(1 downto 0);
    signal VN1532_in3 : std_logic_vector(1 downto 0);
    signal VN1532_in4 : std_logic_vector(1 downto 0);
    signal VN1532_in5 : std_logic_vector(1 downto 0);
    signal VN1533_in0 : std_logic_vector(1 downto 0);
    signal VN1533_in1 : std_logic_vector(1 downto 0);
    signal VN1533_in2 : std_logic_vector(1 downto 0);
    signal VN1533_in3 : std_logic_vector(1 downto 0);
    signal VN1533_in4 : std_logic_vector(1 downto 0);
    signal VN1533_in5 : std_logic_vector(1 downto 0);
    signal VN1534_in0 : std_logic_vector(1 downto 0);
    signal VN1534_in1 : std_logic_vector(1 downto 0);
    signal VN1534_in2 : std_logic_vector(1 downto 0);
    signal VN1534_in3 : std_logic_vector(1 downto 0);
    signal VN1534_in4 : std_logic_vector(1 downto 0);
    signal VN1534_in5 : std_logic_vector(1 downto 0);
    signal VN1535_in0 : std_logic_vector(1 downto 0);
    signal VN1535_in1 : std_logic_vector(1 downto 0);
    signal VN1535_in2 : std_logic_vector(1 downto 0);
    signal VN1535_in3 : std_logic_vector(1 downto 0);
    signal VN1535_in4 : std_logic_vector(1 downto 0);
    signal VN1535_in5 : std_logic_vector(1 downto 0);
    signal VN1536_in0 : std_logic_vector(1 downto 0);
    signal VN1536_in1 : std_logic_vector(1 downto 0);
    signal VN1536_in2 : std_logic_vector(1 downto 0);
    signal VN1536_in3 : std_logic_vector(1 downto 0);
    signal VN1536_in4 : std_logic_vector(1 downto 0);
    signal VN1536_in5 : std_logic_vector(1 downto 0);
    signal VN1537_in0 : std_logic_vector(1 downto 0);
    signal VN1537_in1 : std_logic_vector(1 downto 0);
    signal VN1537_in2 : std_logic_vector(1 downto 0);
    signal VN1537_in3 : std_logic_vector(1 downto 0);
    signal VN1537_in4 : std_logic_vector(1 downto 0);
    signal VN1537_in5 : std_logic_vector(1 downto 0);
    signal VN1538_in0 : std_logic_vector(1 downto 0);
    signal VN1538_in1 : std_logic_vector(1 downto 0);
    signal VN1538_in2 : std_logic_vector(1 downto 0);
    signal VN1538_in3 : std_logic_vector(1 downto 0);
    signal VN1538_in4 : std_logic_vector(1 downto 0);
    signal VN1538_in5 : std_logic_vector(1 downto 0);
    signal VN1539_in0 : std_logic_vector(1 downto 0);
    signal VN1539_in1 : std_logic_vector(1 downto 0);
    signal VN1539_in2 : std_logic_vector(1 downto 0);
    signal VN1539_in3 : std_logic_vector(1 downto 0);
    signal VN1539_in4 : std_logic_vector(1 downto 0);
    signal VN1539_in5 : std_logic_vector(1 downto 0);
    signal VN1540_in0 : std_logic_vector(1 downto 0);
    signal VN1540_in1 : std_logic_vector(1 downto 0);
    signal VN1540_in2 : std_logic_vector(1 downto 0);
    signal VN1540_in3 : std_logic_vector(1 downto 0);
    signal VN1540_in4 : std_logic_vector(1 downto 0);
    signal VN1540_in5 : std_logic_vector(1 downto 0);
    signal VN1541_in0 : std_logic_vector(1 downto 0);
    signal VN1541_in1 : std_logic_vector(1 downto 0);
    signal VN1541_in2 : std_logic_vector(1 downto 0);
    signal VN1541_in3 : std_logic_vector(1 downto 0);
    signal VN1541_in4 : std_logic_vector(1 downto 0);
    signal VN1541_in5 : std_logic_vector(1 downto 0);
    signal VN1542_in0 : std_logic_vector(1 downto 0);
    signal VN1542_in1 : std_logic_vector(1 downto 0);
    signal VN1542_in2 : std_logic_vector(1 downto 0);
    signal VN1542_in3 : std_logic_vector(1 downto 0);
    signal VN1542_in4 : std_logic_vector(1 downto 0);
    signal VN1542_in5 : std_logic_vector(1 downto 0);
    signal VN1543_in0 : std_logic_vector(1 downto 0);
    signal VN1543_in1 : std_logic_vector(1 downto 0);
    signal VN1543_in2 : std_logic_vector(1 downto 0);
    signal VN1543_in3 : std_logic_vector(1 downto 0);
    signal VN1543_in4 : std_logic_vector(1 downto 0);
    signal VN1543_in5 : std_logic_vector(1 downto 0);
    signal VN1544_in0 : std_logic_vector(1 downto 0);
    signal VN1544_in1 : std_logic_vector(1 downto 0);
    signal VN1544_in2 : std_logic_vector(1 downto 0);
    signal VN1544_in3 : std_logic_vector(1 downto 0);
    signal VN1544_in4 : std_logic_vector(1 downto 0);
    signal VN1544_in5 : std_logic_vector(1 downto 0);
    signal VN1545_in0 : std_logic_vector(1 downto 0);
    signal VN1545_in1 : std_logic_vector(1 downto 0);
    signal VN1545_in2 : std_logic_vector(1 downto 0);
    signal VN1545_in3 : std_logic_vector(1 downto 0);
    signal VN1545_in4 : std_logic_vector(1 downto 0);
    signal VN1545_in5 : std_logic_vector(1 downto 0);
    signal VN1546_in0 : std_logic_vector(1 downto 0);
    signal VN1546_in1 : std_logic_vector(1 downto 0);
    signal VN1546_in2 : std_logic_vector(1 downto 0);
    signal VN1546_in3 : std_logic_vector(1 downto 0);
    signal VN1546_in4 : std_logic_vector(1 downto 0);
    signal VN1546_in5 : std_logic_vector(1 downto 0);
    signal VN1547_in0 : std_logic_vector(1 downto 0);
    signal VN1547_in1 : std_logic_vector(1 downto 0);
    signal VN1547_in2 : std_logic_vector(1 downto 0);
    signal VN1547_in3 : std_logic_vector(1 downto 0);
    signal VN1547_in4 : std_logic_vector(1 downto 0);
    signal VN1547_in5 : std_logic_vector(1 downto 0);
    signal VN1548_in0 : std_logic_vector(1 downto 0);
    signal VN1548_in1 : std_logic_vector(1 downto 0);
    signal VN1548_in2 : std_logic_vector(1 downto 0);
    signal VN1548_in3 : std_logic_vector(1 downto 0);
    signal VN1548_in4 : std_logic_vector(1 downto 0);
    signal VN1548_in5 : std_logic_vector(1 downto 0);
    signal VN1549_in0 : std_logic_vector(1 downto 0);
    signal VN1549_in1 : std_logic_vector(1 downto 0);
    signal VN1549_in2 : std_logic_vector(1 downto 0);
    signal VN1549_in3 : std_logic_vector(1 downto 0);
    signal VN1549_in4 : std_logic_vector(1 downto 0);
    signal VN1549_in5 : std_logic_vector(1 downto 0);
    signal VN1550_in0 : std_logic_vector(1 downto 0);
    signal VN1550_in1 : std_logic_vector(1 downto 0);
    signal VN1550_in2 : std_logic_vector(1 downto 0);
    signal VN1550_in3 : std_logic_vector(1 downto 0);
    signal VN1550_in4 : std_logic_vector(1 downto 0);
    signal VN1550_in5 : std_logic_vector(1 downto 0);
    signal VN1551_in0 : std_logic_vector(1 downto 0);
    signal VN1551_in1 : std_logic_vector(1 downto 0);
    signal VN1551_in2 : std_logic_vector(1 downto 0);
    signal VN1551_in3 : std_logic_vector(1 downto 0);
    signal VN1551_in4 : std_logic_vector(1 downto 0);
    signal VN1551_in5 : std_logic_vector(1 downto 0);
    signal VN1552_in0 : std_logic_vector(1 downto 0);
    signal VN1552_in1 : std_logic_vector(1 downto 0);
    signal VN1552_in2 : std_logic_vector(1 downto 0);
    signal VN1552_in3 : std_logic_vector(1 downto 0);
    signal VN1552_in4 : std_logic_vector(1 downto 0);
    signal VN1552_in5 : std_logic_vector(1 downto 0);
    signal VN1553_in0 : std_logic_vector(1 downto 0);
    signal VN1553_in1 : std_logic_vector(1 downto 0);
    signal VN1553_in2 : std_logic_vector(1 downto 0);
    signal VN1553_in3 : std_logic_vector(1 downto 0);
    signal VN1553_in4 : std_logic_vector(1 downto 0);
    signal VN1553_in5 : std_logic_vector(1 downto 0);
    signal VN1554_in0 : std_logic_vector(1 downto 0);
    signal VN1554_in1 : std_logic_vector(1 downto 0);
    signal VN1554_in2 : std_logic_vector(1 downto 0);
    signal VN1554_in3 : std_logic_vector(1 downto 0);
    signal VN1554_in4 : std_logic_vector(1 downto 0);
    signal VN1554_in5 : std_logic_vector(1 downto 0);
    signal VN1555_in0 : std_logic_vector(1 downto 0);
    signal VN1555_in1 : std_logic_vector(1 downto 0);
    signal VN1555_in2 : std_logic_vector(1 downto 0);
    signal VN1555_in3 : std_logic_vector(1 downto 0);
    signal VN1555_in4 : std_logic_vector(1 downto 0);
    signal VN1555_in5 : std_logic_vector(1 downto 0);
    signal VN1556_in0 : std_logic_vector(1 downto 0);
    signal VN1556_in1 : std_logic_vector(1 downto 0);
    signal VN1556_in2 : std_logic_vector(1 downto 0);
    signal VN1556_in3 : std_logic_vector(1 downto 0);
    signal VN1556_in4 : std_logic_vector(1 downto 0);
    signal VN1556_in5 : std_logic_vector(1 downto 0);
    signal VN1557_in0 : std_logic_vector(1 downto 0);
    signal VN1557_in1 : std_logic_vector(1 downto 0);
    signal VN1557_in2 : std_logic_vector(1 downto 0);
    signal VN1557_in3 : std_logic_vector(1 downto 0);
    signal VN1557_in4 : std_logic_vector(1 downto 0);
    signal VN1557_in5 : std_logic_vector(1 downto 0);
    signal VN1558_in0 : std_logic_vector(1 downto 0);
    signal VN1558_in1 : std_logic_vector(1 downto 0);
    signal VN1558_in2 : std_logic_vector(1 downto 0);
    signal VN1558_in3 : std_logic_vector(1 downto 0);
    signal VN1558_in4 : std_logic_vector(1 downto 0);
    signal VN1558_in5 : std_logic_vector(1 downto 0);
    signal VN1559_in0 : std_logic_vector(1 downto 0);
    signal VN1559_in1 : std_logic_vector(1 downto 0);
    signal VN1559_in2 : std_logic_vector(1 downto 0);
    signal VN1559_in3 : std_logic_vector(1 downto 0);
    signal VN1559_in4 : std_logic_vector(1 downto 0);
    signal VN1559_in5 : std_logic_vector(1 downto 0);
    signal VN1560_in0 : std_logic_vector(1 downto 0);
    signal VN1560_in1 : std_logic_vector(1 downto 0);
    signal VN1560_in2 : std_logic_vector(1 downto 0);
    signal VN1560_in3 : std_logic_vector(1 downto 0);
    signal VN1560_in4 : std_logic_vector(1 downto 0);
    signal VN1560_in5 : std_logic_vector(1 downto 0);
    signal VN1561_in0 : std_logic_vector(1 downto 0);
    signal VN1561_in1 : std_logic_vector(1 downto 0);
    signal VN1561_in2 : std_logic_vector(1 downto 0);
    signal VN1561_in3 : std_logic_vector(1 downto 0);
    signal VN1561_in4 : std_logic_vector(1 downto 0);
    signal VN1561_in5 : std_logic_vector(1 downto 0);
    signal VN1562_in0 : std_logic_vector(1 downto 0);
    signal VN1562_in1 : std_logic_vector(1 downto 0);
    signal VN1562_in2 : std_logic_vector(1 downto 0);
    signal VN1562_in3 : std_logic_vector(1 downto 0);
    signal VN1562_in4 : std_logic_vector(1 downto 0);
    signal VN1562_in5 : std_logic_vector(1 downto 0);
    signal VN1563_in0 : std_logic_vector(1 downto 0);
    signal VN1563_in1 : std_logic_vector(1 downto 0);
    signal VN1563_in2 : std_logic_vector(1 downto 0);
    signal VN1563_in3 : std_logic_vector(1 downto 0);
    signal VN1563_in4 : std_logic_vector(1 downto 0);
    signal VN1563_in5 : std_logic_vector(1 downto 0);
    signal VN1564_in0 : std_logic_vector(1 downto 0);
    signal VN1564_in1 : std_logic_vector(1 downto 0);
    signal VN1564_in2 : std_logic_vector(1 downto 0);
    signal VN1564_in3 : std_logic_vector(1 downto 0);
    signal VN1564_in4 : std_logic_vector(1 downto 0);
    signal VN1564_in5 : std_logic_vector(1 downto 0);
    signal VN1565_in0 : std_logic_vector(1 downto 0);
    signal VN1565_in1 : std_logic_vector(1 downto 0);
    signal VN1565_in2 : std_logic_vector(1 downto 0);
    signal VN1565_in3 : std_logic_vector(1 downto 0);
    signal VN1565_in4 : std_logic_vector(1 downto 0);
    signal VN1565_in5 : std_logic_vector(1 downto 0);
    signal VN1566_in0 : std_logic_vector(1 downto 0);
    signal VN1566_in1 : std_logic_vector(1 downto 0);
    signal VN1566_in2 : std_logic_vector(1 downto 0);
    signal VN1566_in3 : std_logic_vector(1 downto 0);
    signal VN1566_in4 : std_logic_vector(1 downto 0);
    signal VN1566_in5 : std_logic_vector(1 downto 0);
    signal VN1567_in0 : std_logic_vector(1 downto 0);
    signal VN1567_in1 : std_logic_vector(1 downto 0);
    signal VN1567_in2 : std_logic_vector(1 downto 0);
    signal VN1567_in3 : std_logic_vector(1 downto 0);
    signal VN1567_in4 : std_logic_vector(1 downto 0);
    signal VN1567_in5 : std_logic_vector(1 downto 0);
    signal VN1568_in0 : std_logic_vector(1 downto 0);
    signal VN1568_in1 : std_logic_vector(1 downto 0);
    signal VN1568_in2 : std_logic_vector(1 downto 0);
    signal VN1568_in3 : std_logic_vector(1 downto 0);
    signal VN1568_in4 : std_logic_vector(1 downto 0);
    signal VN1568_in5 : std_logic_vector(1 downto 0);
    signal VN1569_in0 : std_logic_vector(1 downto 0);
    signal VN1569_in1 : std_logic_vector(1 downto 0);
    signal VN1569_in2 : std_logic_vector(1 downto 0);
    signal VN1569_in3 : std_logic_vector(1 downto 0);
    signal VN1569_in4 : std_logic_vector(1 downto 0);
    signal VN1569_in5 : std_logic_vector(1 downto 0);
    signal VN1570_in0 : std_logic_vector(1 downto 0);
    signal VN1570_in1 : std_logic_vector(1 downto 0);
    signal VN1570_in2 : std_logic_vector(1 downto 0);
    signal VN1570_in3 : std_logic_vector(1 downto 0);
    signal VN1570_in4 : std_logic_vector(1 downto 0);
    signal VN1570_in5 : std_logic_vector(1 downto 0);
    signal VN1571_in0 : std_logic_vector(1 downto 0);
    signal VN1571_in1 : std_logic_vector(1 downto 0);
    signal VN1571_in2 : std_logic_vector(1 downto 0);
    signal VN1571_in3 : std_logic_vector(1 downto 0);
    signal VN1571_in4 : std_logic_vector(1 downto 0);
    signal VN1571_in5 : std_logic_vector(1 downto 0);
    signal VN1572_in0 : std_logic_vector(1 downto 0);
    signal VN1572_in1 : std_logic_vector(1 downto 0);
    signal VN1572_in2 : std_logic_vector(1 downto 0);
    signal VN1572_in3 : std_logic_vector(1 downto 0);
    signal VN1572_in4 : std_logic_vector(1 downto 0);
    signal VN1572_in5 : std_logic_vector(1 downto 0);
    signal VN1573_in0 : std_logic_vector(1 downto 0);
    signal VN1573_in1 : std_logic_vector(1 downto 0);
    signal VN1573_in2 : std_logic_vector(1 downto 0);
    signal VN1573_in3 : std_logic_vector(1 downto 0);
    signal VN1573_in4 : std_logic_vector(1 downto 0);
    signal VN1573_in5 : std_logic_vector(1 downto 0);
    signal VN1574_in0 : std_logic_vector(1 downto 0);
    signal VN1574_in1 : std_logic_vector(1 downto 0);
    signal VN1574_in2 : std_logic_vector(1 downto 0);
    signal VN1574_in3 : std_logic_vector(1 downto 0);
    signal VN1574_in4 : std_logic_vector(1 downto 0);
    signal VN1574_in5 : std_logic_vector(1 downto 0);
    signal VN1575_in0 : std_logic_vector(1 downto 0);
    signal VN1575_in1 : std_logic_vector(1 downto 0);
    signal VN1575_in2 : std_logic_vector(1 downto 0);
    signal VN1575_in3 : std_logic_vector(1 downto 0);
    signal VN1575_in4 : std_logic_vector(1 downto 0);
    signal VN1575_in5 : std_logic_vector(1 downto 0);
    signal VN1576_in0 : std_logic_vector(1 downto 0);
    signal VN1576_in1 : std_logic_vector(1 downto 0);
    signal VN1576_in2 : std_logic_vector(1 downto 0);
    signal VN1576_in3 : std_logic_vector(1 downto 0);
    signal VN1576_in4 : std_logic_vector(1 downto 0);
    signal VN1576_in5 : std_logic_vector(1 downto 0);
    signal VN1577_in0 : std_logic_vector(1 downto 0);
    signal VN1577_in1 : std_logic_vector(1 downto 0);
    signal VN1577_in2 : std_logic_vector(1 downto 0);
    signal VN1577_in3 : std_logic_vector(1 downto 0);
    signal VN1577_in4 : std_logic_vector(1 downto 0);
    signal VN1577_in5 : std_logic_vector(1 downto 0);
    signal VN1578_in0 : std_logic_vector(1 downto 0);
    signal VN1578_in1 : std_logic_vector(1 downto 0);
    signal VN1578_in2 : std_logic_vector(1 downto 0);
    signal VN1578_in3 : std_logic_vector(1 downto 0);
    signal VN1578_in4 : std_logic_vector(1 downto 0);
    signal VN1578_in5 : std_logic_vector(1 downto 0);
    signal VN1579_in0 : std_logic_vector(1 downto 0);
    signal VN1579_in1 : std_logic_vector(1 downto 0);
    signal VN1579_in2 : std_logic_vector(1 downto 0);
    signal VN1579_in3 : std_logic_vector(1 downto 0);
    signal VN1579_in4 : std_logic_vector(1 downto 0);
    signal VN1579_in5 : std_logic_vector(1 downto 0);
    signal VN1580_in0 : std_logic_vector(1 downto 0);
    signal VN1580_in1 : std_logic_vector(1 downto 0);
    signal VN1580_in2 : std_logic_vector(1 downto 0);
    signal VN1580_in3 : std_logic_vector(1 downto 0);
    signal VN1580_in4 : std_logic_vector(1 downto 0);
    signal VN1580_in5 : std_logic_vector(1 downto 0);
    signal VN1581_in0 : std_logic_vector(1 downto 0);
    signal VN1581_in1 : std_logic_vector(1 downto 0);
    signal VN1581_in2 : std_logic_vector(1 downto 0);
    signal VN1581_in3 : std_logic_vector(1 downto 0);
    signal VN1581_in4 : std_logic_vector(1 downto 0);
    signal VN1581_in5 : std_logic_vector(1 downto 0);
    signal VN1582_in0 : std_logic_vector(1 downto 0);
    signal VN1582_in1 : std_logic_vector(1 downto 0);
    signal VN1582_in2 : std_logic_vector(1 downto 0);
    signal VN1582_in3 : std_logic_vector(1 downto 0);
    signal VN1582_in4 : std_logic_vector(1 downto 0);
    signal VN1582_in5 : std_logic_vector(1 downto 0);
    signal VN1583_in0 : std_logic_vector(1 downto 0);
    signal VN1583_in1 : std_logic_vector(1 downto 0);
    signal VN1583_in2 : std_logic_vector(1 downto 0);
    signal VN1583_in3 : std_logic_vector(1 downto 0);
    signal VN1583_in4 : std_logic_vector(1 downto 0);
    signal VN1583_in5 : std_logic_vector(1 downto 0);
    signal VN1584_in0 : std_logic_vector(1 downto 0);
    signal VN1584_in1 : std_logic_vector(1 downto 0);
    signal VN1584_in2 : std_logic_vector(1 downto 0);
    signal VN1584_in3 : std_logic_vector(1 downto 0);
    signal VN1584_in4 : std_logic_vector(1 downto 0);
    signal VN1584_in5 : std_logic_vector(1 downto 0);
    signal VN1585_in0 : std_logic_vector(1 downto 0);
    signal VN1585_in1 : std_logic_vector(1 downto 0);
    signal VN1585_in2 : std_logic_vector(1 downto 0);
    signal VN1585_in3 : std_logic_vector(1 downto 0);
    signal VN1585_in4 : std_logic_vector(1 downto 0);
    signal VN1585_in5 : std_logic_vector(1 downto 0);
    signal VN1586_in0 : std_logic_vector(1 downto 0);
    signal VN1586_in1 : std_logic_vector(1 downto 0);
    signal VN1586_in2 : std_logic_vector(1 downto 0);
    signal VN1586_in3 : std_logic_vector(1 downto 0);
    signal VN1586_in4 : std_logic_vector(1 downto 0);
    signal VN1586_in5 : std_logic_vector(1 downto 0);
    signal VN1587_in0 : std_logic_vector(1 downto 0);
    signal VN1587_in1 : std_logic_vector(1 downto 0);
    signal VN1587_in2 : std_logic_vector(1 downto 0);
    signal VN1587_in3 : std_logic_vector(1 downto 0);
    signal VN1587_in4 : std_logic_vector(1 downto 0);
    signal VN1587_in5 : std_logic_vector(1 downto 0);
    signal VN1588_in0 : std_logic_vector(1 downto 0);
    signal VN1588_in1 : std_logic_vector(1 downto 0);
    signal VN1588_in2 : std_logic_vector(1 downto 0);
    signal VN1588_in3 : std_logic_vector(1 downto 0);
    signal VN1588_in4 : std_logic_vector(1 downto 0);
    signal VN1588_in5 : std_logic_vector(1 downto 0);
    signal VN1589_in0 : std_logic_vector(1 downto 0);
    signal VN1589_in1 : std_logic_vector(1 downto 0);
    signal VN1589_in2 : std_logic_vector(1 downto 0);
    signal VN1589_in3 : std_logic_vector(1 downto 0);
    signal VN1589_in4 : std_logic_vector(1 downto 0);
    signal VN1589_in5 : std_logic_vector(1 downto 0);
    signal VN1590_in0 : std_logic_vector(1 downto 0);
    signal VN1590_in1 : std_logic_vector(1 downto 0);
    signal VN1590_in2 : std_logic_vector(1 downto 0);
    signal VN1590_in3 : std_logic_vector(1 downto 0);
    signal VN1590_in4 : std_logic_vector(1 downto 0);
    signal VN1590_in5 : std_logic_vector(1 downto 0);
    signal VN1591_in0 : std_logic_vector(1 downto 0);
    signal VN1591_in1 : std_logic_vector(1 downto 0);
    signal VN1591_in2 : std_logic_vector(1 downto 0);
    signal VN1591_in3 : std_logic_vector(1 downto 0);
    signal VN1591_in4 : std_logic_vector(1 downto 0);
    signal VN1591_in5 : std_logic_vector(1 downto 0);
    signal VN1592_in0 : std_logic_vector(1 downto 0);
    signal VN1592_in1 : std_logic_vector(1 downto 0);
    signal VN1592_in2 : std_logic_vector(1 downto 0);
    signal VN1592_in3 : std_logic_vector(1 downto 0);
    signal VN1592_in4 : std_logic_vector(1 downto 0);
    signal VN1592_in5 : std_logic_vector(1 downto 0);
    signal VN1593_in0 : std_logic_vector(1 downto 0);
    signal VN1593_in1 : std_logic_vector(1 downto 0);
    signal VN1593_in2 : std_logic_vector(1 downto 0);
    signal VN1593_in3 : std_logic_vector(1 downto 0);
    signal VN1593_in4 : std_logic_vector(1 downto 0);
    signal VN1593_in5 : std_logic_vector(1 downto 0);
    signal VN1594_in0 : std_logic_vector(1 downto 0);
    signal VN1594_in1 : std_logic_vector(1 downto 0);
    signal VN1594_in2 : std_logic_vector(1 downto 0);
    signal VN1594_in3 : std_logic_vector(1 downto 0);
    signal VN1594_in4 : std_logic_vector(1 downto 0);
    signal VN1594_in5 : std_logic_vector(1 downto 0);
    signal VN1595_in0 : std_logic_vector(1 downto 0);
    signal VN1595_in1 : std_logic_vector(1 downto 0);
    signal VN1595_in2 : std_logic_vector(1 downto 0);
    signal VN1595_in3 : std_logic_vector(1 downto 0);
    signal VN1595_in4 : std_logic_vector(1 downto 0);
    signal VN1595_in5 : std_logic_vector(1 downto 0);
    signal VN1596_in0 : std_logic_vector(1 downto 0);
    signal VN1596_in1 : std_logic_vector(1 downto 0);
    signal VN1596_in2 : std_logic_vector(1 downto 0);
    signal VN1596_in3 : std_logic_vector(1 downto 0);
    signal VN1596_in4 : std_logic_vector(1 downto 0);
    signal VN1596_in5 : std_logic_vector(1 downto 0);
    signal VN1597_in0 : std_logic_vector(1 downto 0);
    signal VN1597_in1 : std_logic_vector(1 downto 0);
    signal VN1597_in2 : std_logic_vector(1 downto 0);
    signal VN1597_in3 : std_logic_vector(1 downto 0);
    signal VN1597_in4 : std_logic_vector(1 downto 0);
    signal VN1597_in5 : std_logic_vector(1 downto 0);
    signal VN1598_in0 : std_logic_vector(1 downto 0);
    signal VN1598_in1 : std_logic_vector(1 downto 0);
    signal VN1598_in2 : std_logic_vector(1 downto 0);
    signal VN1598_in3 : std_logic_vector(1 downto 0);
    signal VN1598_in4 : std_logic_vector(1 downto 0);
    signal VN1598_in5 : std_logic_vector(1 downto 0);
    signal VN1599_in0 : std_logic_vector(1 downto 0);
    signal VN1599_in1 : std_logic_vector(1 downto 0);
    signal VN1599_in2 : std_logic_vector(1 downto 0);
    signal VN1599_in3 : std_logic_vector(1 downto 0);
    signal VN1599_in4 : std_logic_vector(1 downto 0);
    signal VN1599_in5 : std_logic_vector(1 downto 0);
    signal VN1600_in0 : std_logic_vector(1 downto 0);
    signal VN1600_in1 : std_logic_vector(1 downto 0);
    signal VN1600_in2 : std_logic_vector(1 downto 0);
    signal VN1600_in3 : std_logic_vector(1 downto 0);
    signal VN1600_in4 : std_logic_vector(1 downto 0);
    signal VN1600_in5 : std_logic_vector(1 downto 0);
    signal VN1601_in0 : std_logic_vector(1 downto 0);
    signal VN1601_in1 : std_logic_vector(1 downto 0);
    signal VN1601_in2 : std_logic_vector(1 downto 0);
    signal VN1601_in3 : std_logic_vector(1 downto 0);
    signal VN1601_in4 : std_logic_vector(1 downto 0);
    signal VN1601_in5 : std_logic_vector(1 downto 0);
    signal VN1602_in0 : std_logic_vector(1 downto 0);
    signal VN1602_in1 : std_logic_vector(1 downto 0);
    signal VN1602_in2 : std_logic_vector(1 downto 0);
    signal VN1602_in3 : std_logic_vector(1 downto 0);
    signal VN1602_in4 : std_logic_vector(1 downto 0);
    signal VN1602_in5 : std_logic_vector(1 downto 0);
    signal VN1603_in0 : std_logic_vector(1 downto 0);
    signal VN1603_in1 : std_logic_vector(1 downto 0);
    signal VN1603_in2 : std_logic_vector(1 downto 0);
    signal VN1603_in3 : std_logic_vector(1 downto 0);
    signal VN1603_in4 : std_logic_vector(1 downto 0);
    signal VN1603_in5 : std_logic_vector(1 downto 0);
    signal VN1604_in0 : std_logic_vector(1 downto 0);
    signal VN1604_in1 : std_logic_vector(1 downto 0);
    signal VN1604_in2 : std_logic_vector(1 downto 0);
    signal VN1604_in3 : std_logic_vector(1 downto 0);
    signal VN1604_in4 : std_logic_vector(1 downto 0);
    signal VN1604_in5 : std_logic_vector(1 downto 0);
    signal VN1605_in0 : std_logic_vector(1 downto 0);
    signal VN1605_in1 : std_logic_vector(1 downto 0);
    signal VN1605_in2 : std_logic_vector(1 downto 0);
    signal VN1605_in3 : std_logic_vector(1 downto 0);
    signal VN1605_in4 : std_logic_vector(1 downto 0);
    signal VN1605_in5 : std_logic_vector(1 downto 0);
    signal VN1606_in0 : std_logic_vector(1 downto 0);
    signal VN1606_in1 : std_logic_vector(1 downto 0);
    signal VN1606_in2 : std_logic_vector(1 downto 0);
    signal VN1606_in3 : std_logic_vector(1 downto 0);
    signal VN1606_in4 : std_logic_vector(1 downto 0);
    signal VN1606_in5 : std_logic_vector(1 downto 0);
    signal VN1607_in0 : std_logic_vector(1 downto 0);
    signal VN1607_in1 : std_logic_vector(1 downto 0);
    signal VN1607_in2 : std_logic_vector(1 downto 0);
    signal VN1607_in3 : std_logic_vector(1 downto 0);
    signal VN1607_in4 : std_logic_vector(1 downto 0);
    signal VN1607_in5 : std_logic_vector(1 downto 0);
    signal VN1608_in0 : std_logic_vector(1 downto 0);
    signal VN1608_in1 : std_logic_vector(1 downto 0);
    signal VN1608_in2 : std_logic_vector(1 downto 0);
    signal VN1608_in3 : std_logic_vector(1 downto 0);
    signal VN1608_in4 : std_logic_vector(1 downto 0);
    signal VN1608_in5 : std_logic_vector(1 downto 0);
    signal VN1609_in0 : std_logic_vector(1 downto 0);
    signal VN1609_in1 : std_logic_vector(1 downto 0);
    signal VN1609_in2 : std_logic_vector(1 downto 0);
    signal VN1609_in3 : std_logic_vector(1 downto 0);
    signal VN1609_in4 : std_logic_vector(1 downto 0);
    signal VN1609_in5 : std_logic_vector(1 downto 0);
    signal VN1610_in0 : std_logic_vector(1 downto 0);
    signal VN1610_in1 : std_logic_vector(1 downto 0);
    signal VN1610_in2 : std_logic_vector(1 downto 0);
    signal VN1610_in3 : std_logic_vector(1 downto 0);
    signal VN1610_in4 : std_logic_vector(1 downto 0);
    signal VN1610_in5 : std_logic_vector(1 downto 0);
    signal VN1611_in0 : std_logic_vector(1 downto 0);
    signal VN1611_in1 : std_logic_vector(1 downto 0);
    signal VN1611_in2 : std_logic_vector(1 downto 0);
    signal VN1611_in3 : std_logic_vector(1 downto 0);
    signal VN1611_in4 : std_logic_vector(1 downto 0);
    signal VN1611_in5 : std_logic_vector(1 downto 0);
    signal VN1612_in0 : std_logic_vector(1 downto 0);
    signal VN1612_in1 : std_logic_vector(1 downto 0);
    signal VN1612_in2 : std_logic_vector(1 downto 0);
    signal VN1612_in3 : std_logic_vector(1 downto 0);
    signal VN1612_in4 : std_logic_vector(1 downto 0);
    signal VN1612_in5 : std_logic_vector(1 downto 0);
    signal VN1613_in0 : std_logic_vector(1 downto 0);
    signal VN1613_in1 : std_logic_vector(1 downto 0);
    signal VN1613_in2 : std_logic_vector(1 downto 0);
    signal VN1613_in3 : std_logic_vector(1 downto 0);
    signal VN1613_in4 : std_logic_vector(1 downto 0);
    signal VN1613_in5 : std_logic_vector(1 downto 0);
    signal VN1614_in0 : std_logic_vector(1 downto 0);
    signal VN1614_in1 : std_logic_vector(1 downto 0);
    signal VN1614_in2 : std_logic_vector(1 downto 0);
    signal VN1614_in3 : std_logic_vector(1 downto 0);
    signal VN1614_in4 : std_logic_vector(1 downto 0);
    signal VN1614_in5 : std_logic_vector(1 downto 0);
    signal VN1615_in0 : std_logic_vector(1 downto 0);
    signal VN1615_in1 : std_logic_vector(1 downto 0);
    signal VN1615_in2 : std_logic_vector(1 downto 0);
    signal VN1615_in3 : std_logic_vector(1 downto 0);
    signal VN1615_in4 : std_logic_vector(1 downto 0);
    signal VN1615_in5 : std_logic_vector(1 downto 0);
    signal VN1616_in0 : std_logic_vector(1 downto 0);
    signal VN1616_in1 : std_logic_vector(1 downto 0);
    signal VN1616_in2 : std_logic_vector(1 downto 0);
    signal VN1616_in3 : std_logic_vector(1 downto 0);
    signal VN1616_in4 : std_logic_vector(1 downto 0);
    signal VN1616_in5 : std_logic_vector(1 downto 0);
    signal VN1617_in0 : std_logic_vector(1 downto 0);
    signal VN1617_in1 : std_logic_vector(1 downto 0);
    signal VN1617_in2 : std_logic_vector(1 downto 0);
    signal VN1617_in3 : std_logic_vector(1 downto 0);
    signal VN1617_in4 : std_logic_vector(1 downto 0);
    signal VN1617_in5 : std_logic_vector(1 downto 0);
    signal VN1618_in0 : std_logic_vector(1 downto 0);
    signal VN1618_in1 : std_logic_vector(1 downto 0);
    signal VN1618_in2 : std_logic_vector(1 downto 0);
    signal VN1618_in3 : std_logic_vector(1 downto 0);
    signal VN1618_in4 : std_logic_vector(1 downto 0);
    signal VN1618_in5 : std_logic_vector(1 downto 0);
    signal VN1619_in0 : std_logic_vector(1 downto 0);
    signal VN1619_in1 : std_logic_vector(1 downto 0);
    signal VN1619_in2 : std_logic_vector(1 downto 0);
    signal VN1619_in3 : std_logic_vector(1 downto 0);
    signal VN1619_in4 : std_logic_vector(1 downto 0);
    signal VN1619_in5 : std_logic_vector(1 downto 0);
    signal VN1620_in0 : std_logic_vector(1 downto 0);
    signal VN1620_in1 : std_logic_vector(1 downto 0);
    signal VN1620_in2 : std_logic_vector(1 downto 0);
    signal VN1620_in3 : std_logic_vector(1 downto 0);
    signal VN1620_in4 : std_logic_vector(1 downto 0);
    signal VN1620_in5 : std_logic_vector(1 downto 0);
    signal VN1621_in0 : std_logic_vector(1 downto 0);
    signal VN1621_in1 : std_logic_vector(1 downto 0);
    signal VN1621_in2 : std_logic_vector(1 downto 0);
    signal VN1621_in3 : std_logic_vector(1 downto 0);
    signal VN1621_in4 : std_logic_vector(1 downto 0);
    signal VN1621_in5 : std_logic_vector(1 downto 0);
    signal VN1622_in0 : std_logic_vector(1 downto 0);
    signal VN1622_in1 : std_logic_vector(1 downto 0);
    signal VN1622_in2 : std_logic_vector(1 downto 0);
    signal VN1622_in3 : std_logic_vector(1 downto 0);
    signal VN1622_in4 : std_logic_vector(1 downto 0);
    signal VN1622_in5 : std_logic_vector(1 downto 0);
    signal VN1623_in0 : std_logic_vector(1 downto 0);
    signal VN1623_in1 : std_logic_vector(1 downto 0);
    signal VN1623_in2 : std_logic_vector(1 downto 0);
    signal VN1623_in3 : std_logic_vector(1 downto 0);
    signal VN1623_in4 : std_logic_vector(1 downto 0);
    signal VN1623_in5 : std_logic_vector(1 downto 0);
    signal VN1624_in0 : std_logic_vector(1 downto 0);
    signal VN1624_in1 : std_logic_vector(1 downto 0);
    signal VN1624_in2 : std_logic_vector(1 downto 0);
    signal VN1624_in3 : std_logic_vector(1 downto 0);
    signal VN1624_in4 : std_logic_vector(1 downto 0);
    signal VN1624_in5 : std_logic_vector(1 downto 0);
    signal VN1625_in0 : std_logic_vector(1 downto 0);
    signal VN1625_in1 : std_logic_vector(1 downto 0);
    signal VN1625_in2 : std_logic_vector(1 downto 0);
    signal VN1625_in3 : std_logic_vector(1 downto 0);
    signal VN1625_in4 : std_logic_vector(1 downto 0);
    signal VN1625_in5 : std_logic_vector(1 downto 0);
    signal VN1626_in0 : std_logic_vector(1 downto 0);
    signal VN1626_in1 : std_logic_vector(1 downto 0);
    signal VN1626_in2 : std_logic_vector(1 downto 0);
    signal VN1626_in3 : std_logic_vector(1 downto 0);
    signal VN1626_in4 : std_logic_vector(1 downto 0);
    signal VN1626_in5 : std_logic_vector(1 downto 0);
    signal VN1627_in0 : std_logic_vector(1 downto 0);
    signal VN1627_in1 : std_logic_vector(1 downto 0);
    signal VN1627_in2 : std_logic_vector(1 downto 0);
    signal VN1627_in3 : std_logic_vector(1 downto 0);
    signal VN1627_in4 : std_logic_vector(1 downto 0);
    signal VN1627_in5 : std_logic_vector(1 downto 0);
    signal VN1628_in0 : std_logic_vector(1 downto 0);
    signal VN1628_in1 : std_logic_vector(1 downto 0);
    signal VN1628_in2 : std_logic_vector(1 downto 0);
    signal VN1628_in3 : std_logic_vector(1 downto 0);
    signal VN1628_in4 : std_logic_vector(1 downto 0);
    signal VN1628_in5 : std_logic_vector(1 downto 0);
    signal VN1629_in0 : std_logic_vector(1 downto 0);
    signal VN1629_in1 : std_logic_vector(1 downto 0);
    signal VN1629_in2 : std_logic_vector(1 downto 0);
    signal VN1629_in3 : std_logic_vector(1 downto 0);
    signal VN1629_in4 : std_logic_vector(1 downto 0);
    signal VN1629_in5 : std_logic_vector(1 downto 0);
    signal VN1630_in0 : std_logic_vector(1 downto 0);
    signal VN1630_in1 : std_logic_vector(1 downto 0);
    signal VN1630_in2 : std_logic_vector(1 downto 0);
    signal VN1630_in3 : std_logic_vector(1 downto 0);
    signal VN1630_in4 : std_logic_vector(1 downto 0);
    signal VN1630_in5 : std_logic_vector(1 downto 0);
    signal VN1631_in0 : std_logic_vector(1 downto 0);
    signal VN1631_in1 : std_logic_vector(1 downto 0);
    signal VN1631_in2 : std_logic_vector(1 downto 0);
    signal VN1631_in3 : std_logic_vector(1 downto 0);
    signal VN1631_in4 : std_logic_vector(1 downto 0);
    signal VN1631_in5 : std_logic_vector(1 downto 0);
    signal VN1632_in0 : std_logic_vector(1 downto 0);
    signal VN1632_in1 : std_logic_vector(1 downto 0);
    signal VN1632_in2 : std_logic_vector(1 downto 0);
    signal VN1632_in3 : std_logic_vector(1 downto 0);
    signal VN1632_in4 : std_logic_vector(1 downto 0);
    signal VN1632_in5 : std_logic_vector(1 downto 0);
    signal VN1633_in0 : std_logic_vector(1 downto 0);
    signal VN1633_in1 : std_logic_vector(1 downto 0);
    signal VN1633_in2 : std_logic_vector(1 downto 0);
    signal VN1633_in3 : std_logic_vector(1 downto 0);
    signal VN1633_in4 : std_logic_vector(1 downto 0);
    signal VN1633_in5 : std_logic_vector(1 downto 0);
    signal VN1634_in0 : std_logic_vector(1 downto 0);
    signal VN1634_in1 : std_logic_vector(1 downto 0);
    signal VN1634_in2 : std_logic_vector(1 downto 0);
    signal VN1634_in3 : std_logic_vector(1 downto 0);
    signal VN1634_in4 : std_logic_vector(1 downto 0);
    signal VN1634_in5 : std_logic_vector(1 downto 0);
    signal VN1635_in0 : std_logic_vector(1 downto 0);
    signal VN1635_in1 : std_logic_vector(1 downto 0);
    signal VN1635_in2 : std_logic_vector(1 downto 0);
    signal VN1635_in3 : std_logic_vector(1 downto 0);
    signal VN1635_in4 : std_logic_vector(1 downto 0);
    signal VN1635_in5 : std_logic_vector(1 downto 0);
    signal VN1636_in0 : std_logic_vector(1 downto 0);
    signal VN1636_in1 : std_logic_vector(1 downto 0);
    signal VN1636_in2 : std_logic_vector(1 downto 0);
    signal VN1636_in3 : std_logic_vector(1 downto 0);
    signal VN1636_in4 : std_logic_vector(1 downto 0);
    signal VN1636_in5 : std_logic_vector(1 downto 0);
    signal VN1637_in0 : std_logic_vector(1 downto 0);
    signal VN1637_in1 : std_logic_vector(1 downto 0);
    signal VN1637_in2 : std_logic_vector(1 downto 0);
    signal VN1637_in3 : std_logic_vector(1 downto 0);
    signal VN1637_in4 : std_logic_vector(1 downto 0);
    signal VN1637_in5 : std_logic_vector(1 downto 0);
    signal VN1638_in0 : std_logic_vector(1 downto 0);
    signal VN1638_in1 : std_logic_vector(1 downto 0);
    signal VN1638_in2 : std_logic_vector(1 downto 0);
    signal VN1638_in3 : std_logic_vector(1 downto 0);
    signal VN1638_in4 : std_logic_vector(1 downto 0);
    signal VN1638_in5 : std_logic_vector(1 downto 0);
    signal VN1639_in0 : std_logic_vector(1 downto 0);
    signal VN1639_in1 : std_logic_vector(1 downto 0);
    signal VN1639_in2 : std_logic_vector(1 downto 0);
    signal VN1639_in3 : std_logic_vector(1 downto 0);
    signal VN1639_in4 : std_logic_vector(1 downto 0);
    signal VN1639_in5 : std_logic_vector(1 downto 0);
    signal VN1640_in0 : std_logic_vector(1 downto 0);
    signal VN1640_in1 : std_logic_vector(1 downto 0);
    signal VN1640_in2 : std_logic_vector(1 downto 0);
    signal VN1640_in3 : std_logic_vector(1 downto 0);
    signal VN1640_in4 : std_logic_vector(1 downto 0);
    signal VN1640_in5 : std_logic_vector(1 downto 0);
    signal VN1641_in0 : std_logic_vector(1 downto 0);
    signal VN1641_in1 : std_logic_vector(1 downto 0);
    signal VN1641_in2 : std_logic_vector(1 downto 0);
    signal VN1641_in3 : std_logic_vector(1 downto 0);
    signal VN1641_in4 : std_logic_vector(1 downto 0);
    signal VN1641_in5 : std_logic_vector(1 downto 0);
    signal VN1642_in0 : std_logic_vector(1 downto 0);
    signal VN1642_in1 : std_logic_vector(1 downto 0);
    signal VN1642_in2 : std_logic_vector(1 downto 0);
    signal VN1642_in3 : std_logic_vector(1 downto 0);
    signal VN1642_in4 : std_logic_vector(1 downto 0);
    signal VN1642_in5 : std_logic_vector(1 downto 0);
    signal VN1643_in0 : std_logic_vector(1 downto 0);
    signal VN1643_in1 : std_logic_vector(1 downto 0);
    signal VN1643_in2 : std_logic_vector(1 downto 0);
    signal VN1643_in3 : std_logic_vector(1 downto 0);
    signal VN1643_in4 : std_logic_vector(1 downto 0);
    signal VN1643_in5 : std_logic_vector(1 downto 0);
    signal VN1644_in0 : std_logic_vector(1 downto 0);
    signal VN1644_in1 : std_logic_vector(1 downto 0);
    signal VN1644_in2 : std_logic_vector(1 downto 0);
    signal VN1644_in3 : std_logic_vector(1 downto 0);
    signal VN1644_in4 : std_logic_vector(1 downto 0);
    signal VN1644_in5 : std_logic_vector(1 downto 0);
    signal VN1645_in0 : std_logic_vector(1 downto 0);
    signal VN1645_in1 : std_logic_vector(1 downto 0);
    signal VN1645_in2 : std_logic_vector(1 downto 0);
    signal VN1645_in3 : std_logic_vector(1 downto 0);
    signal VN1645_in4 : std_logic_vector(1 downto 0);
    signal VN1645_in5 : std_logic_vector(1 downto 0);
    signal VN1646_in0 : std_logic_vector(1 downto 0);
    signal VN1646_in1 : std_logic_vector(1 downto 0);
    signal VN1646_in2 : std_logic_vector(1 downto 0);
    signal VN1646_in3 : std_logic_vector(1 downto 0);
    signal VN1646_in4 : std_logic_vector(1 downto 0);
    signal VN1646_in5 : std_logic_vector(1 downto 0);
    signal VN1647_in0 : std_logic_vector(1 downto 0);
    signal VN1647_in1 : std_logic_vector(1 downto 0);
    signal VN1647_in2 : std_logic_vector(1 downto 0);
    signal VN1647_in3 : std_logic_vector(1 downto 0);
    signal VN1647_in4 : std_logic_vector(1 downto 0);
    signal VN1647_in5 : std_logic_vector(1 downto 0);
    signal VN1648_in0 : std_logic_vector(1 downto 0);
    signal VN1648_in1 : std_logic_vector(1 downto 0);
    signal VN1648_in2 : std_logic_vector(1 downto 0);
    signal VN1648_in3 : std_logic_vector(1 downto 0);
    signal VN1648_in4 : std_logic_vector(1 downto 0);
    signal VN1648_in5 : std_logic_vector(1 downto 0);
    signal VN1649_in0 : std_logic_vector(1 downto 0);
    signal VN1649_in1 : std_logic_vector(1 downto 0);
    signal VN1649_in2 : std_logic_vector(1 downto 0);
    signal VN1649_in3 : std_logic_vector(1 downto 0);
    signal VN1649_in4 : std_logic_vector(1 downto 0);
    signal VN1649_in5 : std_logic_vector(1 downto 0);
    signal VN1650_in0 : std_logic_vector(1 downto 0);
    signal VN1650_in1 : std_logic_vector(1 downto 0);
    signal VN1650_in2 : std_logic_vector(1 downto 0);
    signal VN1650_in3 : std_logic_vector(1 downto 0);
    signal VN1650_in4 : std_logic_vector(1 downto 0);
    signal VN1650_in5 : std_logic_vector(1 downto 0);
    signal VN1651_in0 : std_logic_vector(1 downto 0);
    signal VN1651_in1 : std_logic_vector(1 downto 0);
    signal VN1651_in2 : std_logic_vector(1 downto 0);
    signal VN1651_in3 : std_logic_vector(1 downto 0);
    signal VN1651_in4 : std_logic_vector(1 downto 0);
    signal VN1651_in5 : std_logic_vector(1 downto 0);
    signal VN1652_in0 : std_logic_vector(1 downto 0);
    signal VN1652_in1 : std_logic_vector(1 downto 0);
    signal VN1652_in2 : std_logic_vector(1 downto 0);
    signal VN1652_in3 : std_logic_vector(1 downto 0);
    signal VN1652_in4 : std_logic_vector(1 downto 0);
    signal VN1652_in5 : std_logic_vector(1 downto 0);
    signal VN1653_in0 : std_logic_vector(1 downto 0);
    signal VN1653_in1 : std_logic_vector(1 downto 0);
    signal VN1653_in2 : std_logic_vector(1 downto 0);
    signal VN1653_in3 : std_logic_vector(1 downto 0);
    signal VN1653_in4 : std_logic_vector(1 downto 0);
    signal VN1653_in5 : std_logic_vector(1 downto 0);
    signal VN1654_in0 : std_logic_vector(1 downto 0);
    signal VN1654_in1 : std_logic_vector(1 downto 0);
    signal VN1654_in2 : std_logic_vector(1 downto 0);
    signal VN1654_in3 : std_logic_vector(1 downto 0);
    signal VN1654_in4 : std_logic_vector(1 downto 0);
    signal VN1654_in5 : std_logic_vector(1 downto 0);
    signal VN1655_in0 : std_logic_vector(1 downto 0);
    signal VN1655_in1 : std_logic_vector(1 downto 0);
    signal VN1655_in2 : std_logic_vector(1 downto 0);
    signal VN1655_in3 : std_logic_vector(1 downto 0);
    signal VN1655_in4 : std_logic_vector(1 downto 0);
    signal VN1655_in5 : std_logic_vector(1 downto 0);
    signal VN1656_in0 : std_logic_vector(1 downto 0);
    signal VN1656_in1 : std_logic_vector(1 downto 0);
    signal VN1656_in2 : std_logic_vector(1 downto 0);
    signal VN1656_in3 : std_logic_vector(1 downto 0);
    signal VN1656_in4 : std_logic_vector(1 downto 0);
    signal VN1656_in5 : std_logic_vector(1 downto 0);
    signal VN1657_in0 : std_logic_vector(1 downto 0);
    signal VN1657_in1 : std_logic_vector(1 downto 0);
    signal VN1657_in2 : std_logic_vector(1 downto 0);
    signal VN1657_in3 : std_logic_vector(1 downto 0);
    signal VN1657_in4 : std_logic_vector(1 downto 0);
    signal VN1657_in5 : std_logic_vector(1 downto 0);
    signal VN1658_in0 : std_logic_vector(1 downto 0);
    signal VN1658_in1 : std_logic_vector(1 downto 0);
    signal VN1658_in2 : std_logic_vector(1 downto 0);
    signal VN1658_in3 : std_logic_vector(1 downto 0);
    signal VN1658_in4 : std_logic_vector(1 downto 0);
    signal VN1658_in5 : std_logic_vector(1 downto 0);
    signal VN1659_in0 : std_logic_vector(1 downto 0);
    signal VN1659_in1 : std_logic_vector(1 downto 0);
    signal VN1659_in2 : std_logic_vector(1 downto 0);
    signal VN1659_in3 : std_logic_vector(1 downto 0);
    signal VN1659_in4 : std_logic_vector(1 downto 0);
    signal VN1659_in5 : std_logic_vector(1 downto 0);
    signal VN1660_in0 : std_logic_vector(1 downto 0);
    signal VN1660_in1 : std_logic_vector(1 downto 0);
    signal VN1660_in2 : std_logic_vector(1 downto 0);
    signal VN1660_in3 : std_logic_vector(1 downto 0);
    signal VN1660_in4 : std_logic_vector(1 downto 0);
    signal VN1660_in5 : std_logic_vector(1 downto 0);
    signal VN1661_in0 : std_logic_vector(1 downto 0);
    signal VN1661_in1 : std_logic_vector(1 downto 0);
    signal VN1661_in2 : std_logic_vector(1 downto 0);
    signal VN1661_in3 : std_logic_vector(1 downto 0);
    signal VN1661_in4 : std_logic_vector(1 downto 0);
    signal VN1661_in5 : std_logic_vector(1 downto 0);
    signal VN1662_in0 : std_logic_vector(1 downto 0);
    signal VN1662_in1 : std_logic_vector(1 downto 0);
    signal VN1662_in2 : std_logic_vector(1 downto 0);
    signal VN1662_in3 : std_logic_vector(1 downto 0);
    signal VN1662_in4 : std_logic_vector(1 downto 0);
    signal VN1662_in5 : std_logic_vector(1 downto 0);
    signal VN1663_in0 : std_logic_vector(1 downto 0);
    signal VN1663_in1 : std_logic_vector(1 downto 0);
    signal VN1663_in2 : std_logic_vector(1 downto 0);
    signal VN1663_in3 : std_logic_vector(1 downto 0);
    signal VN1663_in4 : std_logic_vector(1 downto 0);
    signal VN1663_in5 : std_logic_vector(1 downto 0);
    signal VN1664_in0 : std_logic_vector(1 downto 0);
    signal VN1664_in1 : std_logic_vector(1 downto 0);
    signal VN1664_in2 : std_logic_vector(1 downto 0);
    signal VN1664_in3 : std_logic_vector(1 downto 0);
    signal VN1664_in4 : std_logic_vector(1 downto 0);
    signal VN1664_in5 : std_logic_vector(1 downto 0);
    signal VN1665_in0 : std_logic_vector(1 downto 0);
    signal VN1665_in1 : std_logic_vector(1 downto 0);
    signal VN1665_in2 : std_logic_vector(1 downto 0);
    signal VN1665_in3 : std_logic_vector(1 downto 0);
    signal VN1665_in4 : std_logic_vector(1 downto 0);
    signal VN1665_in5 : std_logic_vector(1 downto 0);
    signal VN1666_in0 : std_logic_vector(1 downto 0);
    signal VN1666_in1 : std_logic_vector(1 downto 0);
    signal VN1666_in2 : std_logic_vector(1 downto 0);
    signal VN1666_in3 : std_logic_vector(1 downto 0);
    signal VN1666_in4 : std_logic_vector(1 downto 0);
    signal VN1666_in5 : std_logic_vector(1 downto 0);
    signal VN1667_in0 : std_logic_vector(1 downto 0);
    signal VN1667_in1 : std_logic_vector(1 downto 0);
    signal VN1667_in2 : std_logic_vector(1 downto 0);
    signal VN1667_in3 : std_logic_vector(1 downto 0);
    signal VN1667_in4 : std_logic_vector(1 downto 0);
    signal VN1667_in5 : std_logic_vector(1 downto 0);
    signal VN1668_in0 : std_logic_vector(1 downto 0);
    signal VN1668_in1 : std_logic_vector(1 downto 0);
    signal VN1668_in2 : std_logic_vector(1 downto 0);
    signal VN1668_in3 : std_logic_vector(1 downto 0);
    signal VN1668_in4 : std_logic_vector(1 downto 0);
    signal VN1668_in5 : std_logic_vector(1 downto 0);
    signal VN1669_in0 : std_logic_vector(1 downto 0);
    signal VN1669_in1 : std_logic_vector(1 downto 0);
    signal VN1669_in2 : std_logic_vector(1 downto 0);
    signal VN1669_in3 : std_logic_vector(1 downto 0);
    signal VN1669_in4 : std_logic_vector(1 downto 0);
    signal VN1669_in5 : std_logic_vector(1 downto 0);
    signal VN1670_in0 : std_logic_vector(1 downto 0);
    signal VN1670_in1 : std_logic_vector(1 downto 0);
    signal VN1670_in2 : std_logic_vector(1 downto 0);
    signal VN1670_in3 : std_logic_vector(1 downto 0);
    signal VN1670_in4 : std_logic_vector(1 downto 0);
    signal VN1670_in5 : std_logic_vector(1 downto 0);
    signal VN1671_in0 : std_logic_vector(1 downto 0);
    signal VN1671_in1 : std_logic_vector(1 downto 0);
    signal VN1671_in2 : std_logic_vector(1 downto 0);
    signal VN1671_in3 : std_logic_vector(1 downto 0);
    signal VN1671_in4 : std_logic_vector(1 downto 0);
    signal VN1671_in5 : std_logic_vector(1 downto 0);
    signal VN1672_in0 : std_logic_vector(1 downto 0);
    signal VN1672_in1 : std_logic_vector(1 downto 0);
    signal VN1672_in2 : std_logic_vector(1 downto 0);
    signal VN1672_in3 : std_logic_vector(1 downto 0);
    signal VN1672_in4 : std_logic_vector(1 downto 0);
    signal VN1672_in5 : std_logic_vector(1 downto 0);
    signal VN1673_in0 : std_logic_vector(1 downto 0);
    signal VN1673_in1 : std_logic_vector(1 downto 0);
    signal VN1673_in2 : std_logic_vector(1 downto 0);
    signal VN1673_in3 : std_logic_vector(1 downto 0);
    signal VN1673_in4 : std_logic_vector(1 downto 0);
    signal VN1673_in5 : std_logic_vector(1 downto 0);
    signal VN1674_in0 : std_logic_vector(1 downto 0);
    signal VN1674_in1 : std_logic_vector(1 downto 0);
    signal VN1674_in2 : std_logic_vector(1 downto 0);
    signal VN1674_in3 : std_logic_vector(1 downto 0);
    signal VN1674_in4 : std_logic_vector(1 downto 0);
    signal VN1674_in5 : std_logic_vector(1 downto 0);
    signal VN1675_in0 : std_logic_vector(1 downto 0);
    signal VN1675_in1 : std_logic_vector(1 downto 0);
    signal VN1675_in2 : std_logic_vector(1 downto 0);
    signal VN1675_in3 : std_logic_vector(1 downto 0);
    signal VN1675_in4 : std_logic_vector(1 downto 0);
    signal VN1675_in5 : std_logic_vector(1 downto 0);
    signal VN1676_in0 : std_logic_vector(1 downto 0);
    signal VN1676_in1 : std_logic_vector(1 downto 0);
    signal VN1676_in2 : std_logic_vector(1 downto 0);
    signal VN1676_in3 : std_logic_vector(1 downto 0);
    signal VN1676_in4 : std_logic_vector(1 downto 0);
    signal VN1676_in5 : std_logic_vector(1 downto 0);
    signal VN1677_in0 : std_logic_vector(1 downto 0);
    signal VN1677_in1 : std_logic_vector(1 downto 0);
    signal VN1677_in2 : std_logic_vector(1 downto 0);
    signal VN1677_in3 : std_logic_vector(1 downto 0);
    signal VN1677_in4 : std_logic_vector(1 downto 0);
    signal VN1677_in5 : std_logic_vector(1 downto 0);
    signal VN1678_in0 : std_logic_vector(1 downto 0);
    signal VN1678_in1 : std_logic_vector(1 downto 0);
    signal VN1678_in2 : std_logic_vector(1 downto 0);
    signal VN1678_in3 : std_logic_vector(1 downto 0);
    signal VN1678_in4 : std_logic_vector(1 downto 0);
    signal VN1678_in5 : std_logic_vector(1 downto 0);
    signal VN1679_in0 : std_logic_vector(1 downto 0);
    signal VN1679_in1 : std_logic_vector(1 downto 0);
    signal VN1679_in2 : std_logic_vector(1 downto 0);
    signal VN1679_in3 : std_logic_vector(1 downto 0);
    signal VN1679_in4 : std_logic_vector(1 downto 0);
    signal VN1679_in5 : std_logic_vector(1 downto 0);
    signal VN1680_in0 : std_logic_vector(1 downto 0);
    signal VN1680_in1 : std_logic_vector(1 downto 0);
    signal VN1680_in2 : std_logic_vector(1 downto 0);
    signal VN1680_in3 : std_logic_vector(1 downto 0);
    signal VN1680_in4 : std_logic_vector(1 downto 0);
    signal VN1680_in5 : std_logic_vector(1 downto 0);
    signal VN1681_in0 : std_logic_vector(1 downto 0);
    signal VN1681_in1 : std_logic_vector(1 downto 0);
    signal VN1681_in2 : std_logic_vector(1 downto 0);
    signal VN1681_in3 : std_logic_vector(1 downto 0);
    signal VN1681_in4 : std_logic_vector(1 downto 0);
    signal VN1681_in5 : std_logic_vector(1 downto 0);
    signal VN1682_in0 : std_logic_vector(1 downto 0);
    signal VN1682_in1 : std_logic_vector(1 downto 0);
    signal VN1682_in2 : std_logic_vector(1 downto 0);
    signal VN1682_in3 : std_logic_vector(1 downto 0);
    signal VN1682_in4 : std_logic_vector(1 downto 0);
    signal VN1682_in5 : std_logic_vector(1 downto 0);
    signal VN1683_in0 : std_logic_vector(1 downto 0);
    signal VN1683_in1 : std_logic_vector(1 downto 0);
    signal VN1683_in2 : std_logic_vector(1 downto 0);
    signal VN1683_in3 : std_logic_vector(1 downto 0);
    signal VN1683_in4 : std_logic_vector(1 downto 0);
    signal VN1683_in5 : std_logic_vector(1 downto 0);
    signal VN1684_in0 : std_logic_vector(1 downto 0);
    signal VN1684_in1 : std_logic_vector(1 downto 0);
    signal VN1684_in2 : std_logic_vector(1 downto 0);
    signal VN1684_in3 : std_logic_vector(1 downto 0);
    signal VN1684_in4 : std_logic_vector(1 downto 0);
    signal VN1684_in5 : std_logic_vector(1 downto 0);
    signal VN1685_in0 : std_logic_vector(1 downto 0);
    signal VN1685_in1 : std_logic_vector(1 downto 0);
    signal VN1685_in2 : std_logic_vector(1 downto 0);
    signal VN1685_in3 : std_logic_vector(1 downto 0);
    signal VN1685_in4 : std_logic_vector(1 downto 0);
    signal VN1685_in5 : std_logic_vector(1 downto 0);
    signal VN1686_in0 : std_logic_vector(1 downto 0);
    signal VN1686_in1 : std_logic_vector(1 downto 0);
    signal VN1686_in2 : std_logic_vector(1 downto 0);
    signal VN1686_in3 : std_logic_vector(1 downto 0);
    signal VN1686_in4 : std_logic_vector(1 downto 0);
    signal VN1686_in5 : std_logic_vector(1 downto 0);
    signal VN1687_in0 : std_logic_vector(1 downto 0);
    signal VN1687_in1 : std_logic_vector(1 downto 0);
    signal VN1687_in2 : std_logic_vector(1 downto 0);
    signal VN1687_in3 : std_logic_vector(1 downto 0);
    signal VN1687_in4 : std_logic_vector(1 downto 0);
    signal VN1687_in5 : std_logic_vector(1 downto 0);
    signal VN1688_in0 : std_logic_vector(1 downto 0);
    signal VN1688_in1 : std_logic_vector(1 downto 0);
    signal VN1688_in2 : std_logic_vector(1 downto 0);
    signal VN1688_in3 : std_logic_vector(1 downto 0);
    signal VN1688_in4 : std_logic_vector(1 downto 0);
    signal VN1688_in5 : std_logic_vector(1 downto 0);
    signal VN1689_in0 : std_logic_vector(1 downto 0);
    signal VN1689_in1 : std_logic_vector(1 downto 0);
    signal VN1689_in2 : std_logic_vector(1 downto 0);
    signal VN1689_in3 : std_logic_vector(1 downto 0);
    signal VN1689_in4 : std_logic_vector(1 downto 0);
    signal VN1689_in5 : std_logic_vector(1 downto 0);
    signal VN1690_in0 : std_logic_vector(1 downto 0);
    signal VN1690_in1 : std_logic_vector(1 downto 0);
    signal VN1690_in2 : std_logic_vector(1 downto 0);
    signal VN1690_in3 : std_logic_vector(1 downto 0);
    signal VN1690_in4 : std_logic_vector(1 downto 0);
    signal VN1690_in5 : std_logic_vector(1 downto 0);
    signal VN1691_in0 : std_logic_vector(1 downto 0);
    signal VN1691_in1 : std_logic_vector(1 downto 0);
    signal VN1691_in2 : std_logic_vector(1 downto 0);
    signal VN1691_in3 : std_logic_vector(1 downto 0);
    signal VN1691_in4 : std_logic_vector(1 downto 0);
    signal VN1691_in5 : std_logic_vector(1 downto 0);
    signal VN1692_in0 : std_logic_vector(1 downto 0);
    signal VN1692_in1 : std_logic_vector(1 downto 0);
    signal VN1692_in2 : std_logic_vector(1 downto 0);
    signal VN1692_in3 : std_logic_vector(1 downto 0);
    signal VN1692_in4 : std_logic_vector(1 downto 0);
    signal VN1692_in5 : std_logic_vector(1 downto 0);
    signal VN1693_in0 : std_logic_vector(1 downto 0);
    signal VN1693_in1 : std_logic_vector(1 downto 0);
    signal VN1693_in2 : std_logic_vector(1 downto 0);
    signal VN1693_in3 : std_logic_vector(1 downto 0);
    signal VN1693_in4 : std_logic_vector(1 downto 0);
    signal VN1693_in5 : std_logic_vector(1 downto 0);
    signal VN1694_in0 : std_logic_vector(1 downto 0);
    signal VN1694_in1 : std_logic_vector(1 downto 0);
    signal VN1694_in2 : std_logic_vector(1 downto 0);
    signal VN1694_in3 : std_logic_vector(1 downto 0);
    signal VN1694_in4 : std_logic_vector(1 downto 0);
    signal VN1694_in5 : std_logic_vector(1 downto 0);
    signal VN1695_in0 : std_logic_vector(1 downto 0);
    signal VN1695_in1 : std_logic_vector(1 downto 0);
    signal VN1695_in2 : std_logic_vector(1 downto 0);
    signal VN1695_in3 : std_logic_vector(1 downto 0);
    signal VN1695_in4 : std_logic_vector(1 downto 0);
    signal VN1695_in5 : std_logic_vector(1 downto 0);
    signal VN1696_in0 : std_logic_vector(1 downto 0);
    signal VN1696_in1 : std_logic_vector(1 downto 0);
    signal VN1696_in2 : std_logic_vector(1 downto 0);
    signal VN1696_in3 : std_logic_vector(1 downto 0);
    signal VN1696_in4 : std_logic_vector(1 downto 0);
    signal VN1696_in5 : std_logic_vector(1 downto 0);
    signal VN1697_in0 : std_logic_vector(1 downto 0);
    signal VN1697_in1 : std_logic_vector(1 downto 0);
    signal VN1697_in2 : std_logic_vector(1 downto 0);
    signal VN1697_in3 : std_logic_vector(1 downto 0);
    signal VN1697_in4 : std_logic_vector(1 downto 0);
    signal VN1697_in5 : std_logic_vector(1 downto 0);
    signal VN1698_in0 : std_logic_vector(1 downto 0);
    signal VN1698_in1 : std_logic_vector(1 downto 0);
    signal VN1698_in2 : std_logic_vector(1 downto 0);
    signal VN1698_in3 : std_logic_vector(1 downto 0);
    signal VN1698_in4 : std_logic_vector(1 downto 0);
    signal VN1698_in5 : std_logic_vector(1 downto 0);
    signal VN1699_in0 : std_logic_vector(1 downto 0);
    signal VN1699_in1 : std_logic_vector(1 downto 0);
    signal VN1699_in2 : std_logic_vector(1 downto 0);
    signal VN1699_in3 : std_logic_vector(1 downto 0);
    signal VN1699_in4 : std_logic_vector(1 downto 0);
    signal VN1699_in5 : std_logic_vector(1 downto 0);
    signal VN1700_in0 : std_logic_vector(1 downto 0);
    signal VN1700_in1 : std_logic_vector(1 downto 0);
    signal VN1700_in2 : std_logic_vector(1 downto 0);
    signal VN1700_in3 : std_logic_vector(1 downto 0);
    signal VN1700_in4 : std_logic_vector(1 downto 0);
    signal VN1700_in5 : std_logic_vector(1 downto 0);
    signal VN1701_in0 : std_logic_vector(1 downto 0);
    signal VN1701_in1 : std_logic_vector(1 downto 0);
    signal VN1701_in2 : std_logic_vector(1 downto 0);
    signal VN1701_in3 : std_logic_vector(1 downto 0);
    signal VN1701_in4 : std_logic_vector(1 downto 0);
    signal VN1701_in5 : std_logic_vector(1 downto 0);
    signal VN1702_in0 : std_logic_vector(1 downto 0);
    signal VN1702_in1 : std_logic_vector(1 downto 0);
    signal VN1702_in2 : std_logic_vector(1 downto 0);
    signal VN1702_in3 : std_logic_vector(1 downto 0);
    signal VN1702_in4 : std_logic_vector(1 downto 0);
    signal VN1702_in5 : std_logic_vector(1 downto 0);
    signal VN1703_in0 : std_logic_vector(1 downto 0);
    signal VN1703_in1 : std_logic_vector(1 downto 0);
    signal VN1703_in2 : std_logic_vector(1 downto 0);
    signal VN1703_in3 : std_logic_vector(1 downto 0);
    signal VN1703_in4 : std_logic_vector(1 downto 0);
    signal VN1703_in5 : std_logic_vector(1 downto 0);
    signal VN1704_in0 : std_logic_vector(1 downto 0);
    signal VN1704_in1 : std_logic_vector(1 downto 0);
    signal VN1704_in2 : std_logic_vector(1 downto 0);
    signal VN1704_in3 : std_logic_vector(1 downto 0);
    signal VN1704_in4 : std_logic_vector(1 downto 0);
    signal VN1704_in5 : std_logic_vector(1 downto 0);
    signal VN1705_in0 : std_logic_vector(1 downto 0);
    signal VN1705_in1 : std_logic_vector(1 downto 0);
    signal VN1705_in2 : std_logic_vector(1 downto 0);
    signal VN1705_in3 : std_logic_vector(1 downto 0);
    signal VN1705_in4 : std_logic_vector(1 downto 0);
    signal VN1705_in5 : std_logic_vector(1 downto 0);
    signal VN1706_in0 : std_logic_vector(1 downto 0);
    signal VN1706_in1 : std_logic_vector(1 downto 0);
    signal VN1706_in2 : std_logic_vector(1 downto 0);
    signal VN1706_in3 : std_logic_vector(1 downto 0);
    signal VN1706_in4 : std_logic_vector(1 downto 0);
    signal VN1706_in5 : std_logic_vector(1 downto 0);
    signal VN1707_in0 : std_logic_vector(1 downto 0);
    signal VN1707_in1 : std_logic_vector(1 downto 0);
    signal VN1707_in2 : std_logic_vector(1 downto 0);
    signal VN1707_in3 : std_logic_vector(1 downto 0);
    signal VN1707_in4 : std_logic_vector(1 downto 0);
    signal VN1707_in5 : std_logic_vector(1 downto 0);
    signal VN1708_in0 : std_logic_vector(1 downto 0);
    signal VN1708_in1 : std_logic_vector(1 downto 0);
    signal VN1708_in2 : std_logic_vector(1 downto 0);
    signal VN1708_in3 : std_logic_vector(1 downto 0);
    signal VN1708_in4 : std_logic_vector(1 downto 0);
    signal VN1708_in5 : std_logic_vector(1 downto 0);
    signal VN1709_in0 : std_logic_vector(1 downto 0);
    signal VN1709_in1 : std_logic_vector(1 downto 0);
    signal VN1709_in2 : std_logic_vector(1 downto 0);
    signal VN1709_in3 : std_logic_vector(1 downto 0);
    signal VN1709_in4 : std_logic_vector(1 downto 0);
    signal VN1709_in5 : std_logic_vector(1 downto 0);
    signal VN1710_in0 : std_logic_vector(1 downto 0);
    signal VN1710_in1 : std_logic_vector(1 downto 0);
    signal VN1710_in2 : std_logic_vector(1 downto 0);
    signal VN1710_in3 : std_logic_vector(1 downto 0);
    signal VN1710_in4 : std_logic_vector(1 downto 0);
    signal VN1710_in5 : std_logic_vector(1 downto 0);
    signal VN1711_in0 : std_logic_vector(1 downto 0);
    signal VN1711_in1 : std_logic_vector(1 downto 0);
    signal VN1711_in2 : std_logic_vector(1 downto 0);
    signal VN1711_in3 : std_logic_vector(1 downto 0);
    signal VN1711_in4 : std_logic_vector(1 downto 0);
    signal VN1711_in5 : std_logic_vector(1 downto 0);
    signal VN1712_in0 : std_logic_vector(1 downto 0);
    signal VN1712_in1 : std_logic_vector(1 downto 0);
    signal VN1712_in2 : std_logic_vector(1 downto 0);
    signal VN1712_in3 : std_logic_vector(1 downto 0);
    signal VN1712_in4 : std_logic_vector(1 downto 0);
    signal VN1712_in5 : std_logic_vector(1 downto 0);
    signal VN1713_in0 : std_logic_vector(1 downto 0);
    signal VN1713_in1 : std_logic_vector(1 downto 0);
    signal VN1713_in2 : std_logic_vector(1 downto 0);
    signal VN1713_in3 : std_logic_vector(1 downto 0);
    signal VN1713_in4 : std_logic_vector(1 downto 0);
    signal VN1713_in5 : std_logic_vector(1 downto 0);
    signal VN1714_in0 : std_logic_vector(1 downto 0);
    signal VN1714_in1 : std_logic_vector(1 downto 0);
    signal VN1714_in2 : std_logic_vector(1 downto 0);
    signal VN1714_in3 : std_logic_vector(1 downto 0);
    signal VN1714_in4 : std_logic_vector(1 downto 0);
    signal VN1714_in5 : std_logic_vector(1 downto 0);
    signal VN1715_in0 : std_logic_vector(1 downto 0);
    signal VN1715_in1 : std_logic_vector(1 downto 0);
    signal VN1715_in2 : std_logic_vector(1 downto 0);
    signal VN1715_in3 : std_logic_vector(1 downto 0);
    signal VN1715_in4 : std_logic_vector(1 downto 0);
    signal VN1715_in5 : std_logic_vector(1 downto 0);
    signal VN1716_in0 : std_logic_vector(1 downto 0);
    signal VN1716_in1 : std_logic_vector(1 downto 0);
    signal VN1716_in2 : std_logic_vector(1 downto 0);
    signal VN1716_in3 : std_logic_vector(1 downto 0);
    signal VN1716_in4 : std_logic_vector(1 downto 0);
    signal VN1716_in5 : std_logic_vector(1 downto 0);
    signal VN1717_in0 : std_logic_vector(1 downto 0);
    signal VN1717_in1 : std_logic_vector(1 downto 0);
    signal VN1717_in2 : std_logic_vector(1 downto 0);
    signal VN1717_in3 : std_logic_vector(1 downto 0);
    signal VN1717_in4 : std_logic_vector(1 downto 0);
    signal VN1717_in5 : std_logic_vector(1 downto 0);
    signal VN1718_in0 : std_logic_vector(1 downto 0);
    signal VN1718_in1 : std_logic_vector(1 downto 0);
    signal VN1718_in2 : std_logic_vector(1 downto 0);
    signal VN1718_in3 : std_logic_vector(1 downto 0);
    signal VN1718_in4 : std_logic_vector(1 downto 0);
    signal VN1718_in5 : std_logic_vector(1 downto 0);
    signal VN1719_in0 : std_logic_vector(1 downto 0);
    signal VN1719_in1 : std_logic_vector(1 downto 0);
    signal VN1719_in2 : std_logic_vector(1 downto 0);
    signal VN1719_in3 : std_logic_vector(1 downto 0);
    signal VN1719_in4 : std_logic_vector(1 downto 0);
    signal VN1719_in5 : std_logic_vector(1 downto 0);
    signal VN1720_in0 : std_logic_vector(1 downto 0);
    signal VN1720_in1 : std_logic_vector(1 downto 0);
    signal VN1720_in2 : std_logic_vector(1 downto 0);
    signal VN1720_in3 : std_logic_vector(1 downto 0);
    signal VN1720_in4 : std_logic_vector(1 downto 0);
    signal VN1720_in5 : std_logic_vector(1 downto 0);
    signal VN1721_in0 : std_logic_vector(1 downto 0);
    signal VN1721_in1 : std_logic_vector(1 downto 0);
    signal VN1721_in2 : std_logic_vector(1 downto 0);
    signal VN1721_in3 : std_logic_vector(1 downto 0);
    signal VN1721_in4 : std_logic_vector(1 downto 0);
    signal VN1721_in5 : std_logic_vector(1 downto 0);
    signal VN1722_in0 : std_logic_vector(1 downto 0);
    signal VN1722_in1 : std_logic_vector(1 downto 0);
    signal VN1722_in2 : std_logic_vector(1 downto 0);
    signal VN1722_in3 : std_logic_vector(1 downto 0);
    signal VN1722_in4 : std_logic_vector(1 downto 0);
    signal VN1722_in5 : std_logic_vector(1 downto 0);
    signal VN1723_in0 : std_logic_vector(1 downto 0);
    signal VN1723_in1 : std_logic_vector(1 downto 0);
    signal VN1723_in2 : std_logic_vector(1 downto 0);
    signal VN1723_in3 : std_logic_vector(1 downto 0);
    signal VN1723_in4 : std_logic_vector(1 downto 0);
    signal VN1723_in5 : std_logic_vector(1 downto 0);
    signal VN1724_in0 : std_logic_vector(1 downto 0);
    signal VN1724_in1 : std_logic_vector(1 downto 0);
    signal VN1724_in2 : std_logic_vector(1 downto 0);
    signal VN1724_in3 : std_logic_vector(1 downto 0);
    signal VN1724_in4 : std_logic_vector(1 downto 0);
    signal VN1724_in5 : std_logic_vector(1 downto 0);
    signal VN1725_in0 : std_logic_vector(1 downto 0);
    signal VN1725_in1 : std_logic_vector(1 downto 0);
    signal VN1725_in2 : std_logic_vector(1 downto 0);
    signal VN1725_in3 : std_logic_vector(1 downto 0);
    signal VN1725_in4 : std_logic_vector(1 downto 0);
    signal VN1725_in5 : std_logic_vector(1 downto 0);
    signal VN1726_in0 : std_logic_vector(1 downto 0);
    signal VN1726_in1 : std_logic_vector(1 downto 0);
    signal VN1726_in2 : std_logic_vector(1 downto 0);
    signal VN1726_in3 : std_logic_vector(1 downto 0);
    signal VN1726_in4 : std_logic_vector(1 downto 0);
    signal VN1726_in5 : std_logic_vector(1 downto 0);
    signal VN1727_in0 : std_logic_vector(1 downto 0);
    signal VN1727_in1 : std_logic_vector(1 downto 0);
    signal VN1727_in2 : std_logic_vector(1 downto 0);
    signal VN1727_in3 : std_logic_vector(1 downto 0);
    signal VN1727_in4 : std_logic_vector(1 downto 0);
    signal VN1727_in5 : std_logic_vector(1 downto 0);
    signal VN1728_in0 : std_logic_vector(1 downto 0);
    signal VN1728_in1 : std_logic_vector(1 downto 0);
    signal VN1728_in2 : std_logic_vector(1 downto 0);
    signal VN1728_in3 : std_logic_vector(1 downto 0);
    signal VN1728_in4 : std_logic_vector(1 downto 0);
    signal VN1728_in5 : std_logic_vector(1 downto 0);
    signal VN1729_in0 : std_logic_vector(1 downto 0);
    signal VN1729_in1 : std_logic_vector(1 downto 0);
    signal VN1729_in2 : std_logic_vector(1 downto 0);
    signal VN1729_in3 : std_logic_vector(1 downto 0);
    signal VN1729_in4 : std_logic_vector(1 downto 0);
    signal VN1729_in5 : std_logic_vector(1 downto 0);
    signal VN1730_in0 : std_logic_vector(1 downto 0);
    signal VN1730_in1 : std_logic_vector(1 downto 0);
    signal VN1730_in2 : std_logic_vector(1 downto 0);
    signal VN1730_in3 : std_logic_vector(1 downto 0);
    signal VN1730_in4 : std_logic_vector(1 downto 0);
    signal VN1730_in5 : std_logic_vector(1 downto 0);
    signal VN1731_in0 : std_logic_vector(1 downto 0);
    signal VN1731_in1 : std_logic_vector(1 downto 0);
    signal VN1731_in2 : std_logic_vector(1 downto 0);
    signal VN1731_in3 : std_logic_vector(1 downto 0);
    signal VN1731_in4 : std_logic_vector(1 downto 0);
    signal VN1731_in5 : std_logic_vector(1 downto 0);
    signal VN1732_in0 : std_logic_vector(1 downto 0);
    signal VN1732_in1 : std_logic_vector(1 downto 0);
    signal VN1732_in2 : std_logic_vector(1 downto 0);
    signal VN1732_in3 : std_logic_vector(1 downto 0);
    signal VN1732_in4 : std_logic_vector(1 downto 0);
    signal VN1732_in5 : std_logic_vector(1 downto 0);
    signal VN1733_in0 : std_logic_vector(1 downto 0);
    signal VN1733_in1 : std_logic_vector(1 downto 0);
    signal VN1733_in2 : std_logic_vector(1 downto 0);
    signal VN1733_in3 : std_logic_vector(1 downto 0);
    signal VN1733_in4 : std_logic_vector(1 downto 0);
    signal VN1733_in5 : std_logic_vector(1 downto 0);
    signal VN1734_in0 : std_logic_vector(1 downto 0);
    signal VN1734_in1 : std_logic_vector(1 downto 0);
    signal VN1734_in2 : std_logic_vector(1 downto 0);
    signal VN1734_in3 : std_logic_vector(1 downto 0);
    signal VN1734_in4 : std_logic_vector(1 downto 0);
    signal VN1734_in5 : std_logic_vector(1 downto 0);
    signal VN1735_in0 : std_logic_vector(1 downto 0);
    signal VN1735_in1 : std_logic_vector(1 downto 0);
    signal VN1735_in2 : std_logic_vector(1 downto 0);
    signal VN1735_in3 : std_logic_vector(1 downto 0);
    signal VN1735_in4 : std_logic_vector(1 downto 0);
    signal VN1735_in5 : std_logic_vector(1 downto 0);
    signal VN1736_in0 : std_logic_vector(1 downto 0);
    signal VN1736_in1 : std_logic_vector(1 downto 0);
    signal VN1736_in2 : std_logic_vector(1 downto 0);
    signal VN1736_in3 : std_logic_vector(1 downto 0);
    signal VN1736_in4 : std_logic_vector(1 downto 0);
    signal VN1736_in5 : std_logic_vector(1 downto 0);
    signal VN1737_in0 : std_logic_vector(1 downto 0);
    signal VN1737_in1 : std_logic_vector(1 downto 0);
    signal VN1737_in2 : std_logic_vector(1 downto 0);
    signal VN1737_in3 : std_logic_vector(1 downto 0);
    signal VN1737_in4 : std_logic_vector(1 downto 0);
    signal VN1737_in5 : std_logic_vector(1 downto 0);
    signal VN1738_in0 : std_logic_vector(1 downto 0);
    signal VN1738_in1 : std_logic_vector(1 downto 0);
    signal VN1738_in2 : std_logic_vector(1 downto 0);
    signal VN1738_in3 : std_logic_vector(1 downto 0);
    signal VN1738_in4 : std_logic_vector(1 downto 0);
    signal VN1738_in5 : std_logic_vector(1 downto 0);
    signal VN1739_in0 : std_logic_vector(1 downto 0);
    signal VN1739_in1 : std_logic_vector(1 downto 0);
    signal VN1739_in2 : std_logic_vector(1 downto 0);
    signal VN1739_in3 : std_logic_vector(1 downto 0);
    signal VN1739_in4 : std_logic_vector(1 downto 0);
    signal VN1739_in5 : std_logic_vector(1 downto 0);
    signal VN1740_in0 : std_logic_vector(1 downto 0);
    signal VN1740_in1 : std_logic_vector(1 downto 0);
    signal VN1740_in2 : std_logic_vector(1 downto 0);
    signal VN1740_in3 : std_logic_vector(1 downto 0);
    signal VN1740_in4 : std_logic_vector(1 downto 0);
    signal VN1740_in5 : std_logic_vector(1 downto 0);
    signal VN1741_in0 : std_logic_vector(1 downto 0);
    signal VN1741_in1 : std_logic_vector(1 downto 0);
    signal VN1741_in2 : std_logic_vector(1 downto 0);
    signal VN1741_in3 : std_logic_vector(1 downto 0);
    signal VN1741_in4 : std_logic_vector(1 downto 0);
    signal VN1741_in5 : std_logic_vector(1 downto 0);
    signal VN1742_in0 : std_logic_vector(1 downto 0);
    signal VN1742_in1 : std_logic_vector(1 downto 0);
    signal VN1742_in2 : std_logic_vector(1 downto 0);
    signal VN1742_in3 : std_logic_vector(1 downto 0);
    signal VN1742_in4 : std_logic_vector(1 downto 0);
    signal VN1742_in5 : std_logic_vector(1 downto 0);
    signal VN1743_in0 : std_logic_vector(1 downto 0);
    signal VN1743_in1 : std_logic_vector(1 downto 0);
    signal VN1743_in2 : std_logic_vector(1 downto 0);
    signal VN1743_in3 : std_logic_vector(1 downto 0);
    signal VN1743_in4 : std_logic_vector(1 downto 0);
    signal VN1743_in5 : std_logic_vector(1 downto 0);
    signal VN1744_in0 : std_logic_vector(1 downto 0);
    signal VN1744_in1 : std_logic_vector(1 downto 0);
    signal VN1744_in2 : std_logic_vector(1 downto 0);
    signal VN1744_in3 : std_logic_vector(1 downto 0);
    signal VN1744_in4 : std_logic_vector(1 downto 0);
    signal VN1744_in5 : std_logic_vector(1 downto 0);
    signal VN1745_in0 : std_logic_vector(1 downto 0);
    signal VN1745_in1 : std_logic_vector(1 downto 0);
    signal VN1745_in2 : std_logic_vector(1 downto 0);
    signal VN1745_in3 : std_logic_vector(1 downto 0);
    signal VN1745_in4 : std_logic_vector(1 downto 0);
    signal VN1745_in5 : std_logic_vector(1 downto 0);
    signal VN1746_in0 : std_logic_vector(1 downto 0);
    signal VN1746_in1 : std_logic_vector(1 downto 0);
    signal VN1746_in2 : std_logic_vector(1 downto 0);
    signal VN1746_in3 : std_logic_vector(1 downto 0);
    signal VN1746_in4 : std_logic_vector(1 downto 0);
    signal VN1746_in5 : std_logic_vector(1 downto 0);
    signal VN1747_in0 : std_logic_vector(1 downto 0);
    signal VN1747_in1 : std_logic_vector(1 downto 0);
    signal VN1747_in2 : std_logic_vector(1 downto 0);
    signal VN1747_in3 : std_logic_vector(1 downto 0);
    signal VN1747_in4 : std_logic_vector(1 downto 0);
    signal VN1747_in5 : std_logic_vector(1 downto 0);
    signal VN1748_in0 : std_logic_vector(1 downto 0);
    signal VN1748_in1 : std_logic_vector(1 downto 0);
    signal VN1748_in2 : std_logic_vector(1 downto 0);
    signal VN1748_in3 : std_logic_vector(1 downto 0);
    signal VN1748_in4 : std_logic_vector(1 downto 0);
    signal VN1748_in5 : std_logic_vector(1 downto 0);
    signal VN1749_in0 : std_logic_vector(1 downto 0);
    signal VN1749_in1 : std_logic_vector(1 downto 0);
    signal VN1749_in2 : std_logic_vector(1 downto 0);
    signal VN1749_in3 : std_logic_vector(1 downto 0);
    signal VN1749_in4 : std_logic_vector(1 downto 0);
    signal VN1749_in5 : std_logic_vector(1 downto 0);
    signal VN1750_in0 : std_logic_vector(1 downto 0);
    signal VN1750_in1 : std_logic_vector(1 downto 0);
    signal VN1750_in2 : std_logic_vector(1 downto 0);
    signal VN1750_in3 : std_logic_vector(1 downto 0);
    signal VN1750_in4 : std_logic_vector(1 downto 0);
    signal VN1750_in5 : std_logic_vector(1 downto 0);
    signal VN1751_in0 : std_logic_vector(1 downto 0);
    signal VN1751_in1 : std_logic_vector(1 downto 0);
    signal VN1751_in2 : std_logic_vector(1 downto 0);
    signal VN1751_in3 : std_logic_vector(1 downto 0);
    signal VN1751_in4 : std_logic_vector(1 downto 0);
    signal VN1751_in5 : std_logic_vector(1 downto 0);
    signal VN1752_in0 : std_logic_vector(1 downto 0);
    signal VN1752_in1 : std_logic_vector(1 downto 0);
    signal VN1752_in2 : std_logic_vector(1 downto 0);
    signal VN1752_in3 : std_logic_vector(1 downto 0);
    signal VN1752_in4 : std_logic_vector(1 downto 0);
    signal VN1752_in5 : std_logic_vector(1 downto 0);
    signal VN1753_in0 : std_logic_vector(1 downto 0);
    signal VN1753_in1 : std_logic_vector(1 downto 0);
    signal VN1753_in2 : std_logic_vector(1 downto 0);
    signal VN1753_in3 : std_logic_vector(1 downto 0);
    signal VN1753_in4 : std_logic_vector(1 downto 0);
    signal VN1753_in5 : std_logic_vector(1 downto 0);
    signal VN1754_in0 : std_logic_vector(1 downto 0);
    signal VN1754_in1 : std_logic_vector(1 downto 0);
    signal VN1754_in2 : std_logic_vector(1 downto 0);
    signal VN1754_in3 : std_logic_vector(1 downto 0);
    signal VN1754_in4 : std_logic_vector(1 downto 0);
    signal VN1754_in5 : std_logic_vector(1 downto 0);
    signal VN1755_in0 : std_logic_vector(1 downto 0);
    signal VN1755_in1 : std_logic_vector(1 downto 0);
    signal VN1755_in2 : std_logic_vector(1 downto 0);
    signal VN1755_in3 : std_logic_vector(1 downto 0);
    signal VN1755_in4 : std_logic_vector(1 downto 0);
    signal VN1755_in5 : std_logic_vector(1 downto 0);
    signal VN1756_in0 : std_logic_vector(1 downto 0);
    signal VN1756_in1 : std_logic_vector(1 downto 0);
    signal VN1756_in2 : std_logic_vector(1 downto 0);
    signal VN1756_in3 : std_logic_vector(1 downto 0);
    signal VN1756_in4 : std_logic_vector(1 downto 0);
    signal VN1756_in5 : std_logic_vector(1 downto 0);
    signal VN1757_in0 : std_logic_vector(1 downto 0);
    signal VN1757_in1 : std_logic_vector(1 downto 0);
    signal VN1757_in2 : std_logic_vector(1 downto 0);
    signal VN1757_in3 : std_logic_vector(1 downto 0);
    signal VN1757_in4 : std_logic_vector(1 downto 0);
    signal VN1757_in5 : std_logic_vector(1 downto 0);
    signal VN1758_in0 : std_logic_vector(1 downto 0);
    signal VN1758_in1 : std_logic_vector(1 downto 0);
    signal VN1758_in2 : std_logic_vector(1 downto 0);
    signal VN1758_in3 : std_logic_vector(1 downto 0);
    signal VN1758_in4 : std_logic_vector(1 downto 0);
    signal VN1758_in5 : std_logic_vector(1 downto 0);
    signal VN1759_in0 : std_logic_vector(1 downto 0);
    signal VN1759_in1 : std_logic_vector(1 downto 0);
    signal VN1759_in2 : std_logic_vector(1 downto 0);
    signal VN1759_in3 : std_logic_vector(1 downto 0);
    signal VN1759_in4 : std_logic_vector(1 downto 0);
    signal VN1759_in5 : std_logic_vector(1 downto 0);
    signal VN1760_in0 : std_logic_vector(1 downto 0);
    signal VN1760_in1 : std_logic_vector(1 downto 0);
    signal VN1760_in2 : std_logic_vector(1 downto 0);
    signal VN1760_in3 : std_logic_vector(1 downto 0);
    signal VN1760_in4 : std_logic_vector(1 downto 0);
    signal VN1760_in5 : std_logic_vector(1 downto 0);
    signal VN1761_in0 : std_logic_vector(1 downto 0);
    signal VN1761_in1 : std_logic_vector(1 downto 0);
    signal VN1761_in2 : std_logic_vector(1 downto 0);
    signal VN1761_in3 : std_logic_vector(1 downto 0);
    signal VN1761_in4 : std_logic_vector(1 downto 0);
    signal VN1761_in5 : std_logic_vector(1 downto 0);
    signal VN1762_in0 : std_logic_vector(1 downto 0);
    signal VN1762_in1 : std_logic_vector(1 downto 0);
    signal VN1762_in2 : std_logic_vector(1 downto 0);
    signal VN1762_in3 : std_logic_vector(1 downto 0);
    signal VN1762_in4 : std_logic_vector(1 downto 0);
    signal VN1762_in5 : std_logic_vector(1 downto 0);
    signal VN1763_in0 : std_logic_vector(1 downto 0);
    signal VN1763_in1 : std_logic_vector(1 downto 0);
    signal VN1763_in2 : std_logic_vector(1 downto 0);
    signal VN1763_in3 : std_logic_vector(1 downto 0);
    signal VN1763_in4 : std_logic_vector(1 downto 0);
    signal VN1763_in5 : std_logic_vector(1 downto 0);
    signal VN1764_in0 : std_logic_vector(1 downto 0);
    signal VN1764_in1 : std_logic_vector(1 downto 0);
    signal VN1764_in2 : std_logic_vector(1 downto 0);
    signal VN1764_in3 : std_logic_vector(1 downto 0);
    signal VN1764_in4 : std_logic_vector(1 downto 0);
    signal VN1764_in5 : std_logic_vector(1 downto 0);
    signal VN1765_in0 : std_logic_vector(1 downto 0);
    signal VN1765_in1 : std_logic_vector(1 downto 0);
    signal VN1765_in2 : std_logic_vector(1 downto 0);
    signal VN1765_in3 : std_logic_vector(1 downto 0);
    signal VN1765_in4 : std_logic_vector(1 downto 0);
    signal VN1765_in5 : std_logic_vector(1 downto 0);
    signal VN1766_in0 : std_logic_vector(1 downto 0);
    signal VN1766_in1 : std_logic_vector(1 downto 0);
    signal VN1766_in2 : std_logic_vector(1 downto 0);
    signal VN1766_in3 : std_logic_vector(1 downto 0);
    signal VN1766_in4 : std_logic_vector(1 downto 0);
    signal VN1766_in5 : std_logic_vector(1 downto 0);
    signal VN1767_in0 : std_logic_vector(1 downto 0);
    signal VN1767_in1 : std_logic_vector(1 downto 0);
    signal VN1767_in2 : std_logic_vector(1 downto 0);
    signal VN1767_in3 : std_logic_vector(1 downto 0);
    signal VN1767_in4 : std_logic_vector(1 downto 0);
    signal VN1767_in5 : std_logic_vector(1 downto 0);
    signal VN1768_in0 : std_logic_vector(1 downto 0);
    signal VN1768_in1 : std_logic_vector(1 downto 0);
    signal VN1768_in2 : std_logic_vector(1 downto 0);
    signal VN1768_in3 : std_logic_vector(1 downto 0);
    signal VN1768_in4 : std_logic_vector(1 downto 0);
    signal VN1768_in5 : std_logic_vector(1 downto 0);
    signal VN1769_in0 : std_logic_vector(1 downto 0);
    signal VN1769_in1 : std_logic_vector(1 downto 0);
    signal VN1769_in2 : std_logic_vector(1 downto 0);
    signal VN1769_in3 : std_logic_vector(1 downto 0);
    signal VN1769_in4 : std_logic_vector(1 downto 0);
    signal VN1769_in5 : std_logic_vector(1 downto 0);
    signal VN1770_in0 : std_logic_vector(1 downto 0);
    signal VN1770_in1 : std_logic_vector(1 downto 0);
    signal VN1770_in2 : std_logic_vector(1 downto 0);
    signal VN1770_in3 : std_logic_vector(1 downto 0);
    signal VN1770_in4 : std_logic_vector(1 downto 0);
    signal VN1770_in5 : std_logic_vector(1 downto 0);
    signal VN1771_in0 : std_logic_vector(1 downto 0);
    signal VN1771_in1 : std_logic_vector(1 downto 0);
    signal VN1771_in2 : std_logic_vector(1 downto 0);
    signal VN1771_in3 : std_logic_vector(1 downto 0);
    signal VN1771_in4 : std_logic_vector(1 downto 0);
    signal VN1771_in5 : std_logic_vector(1 downto 0);
    signal VN1772_in0 : std_logic_vector(1 downto 0);
    signal VN1772_in1 : std_logic_vector(1 downto 0);
    signal VN1772_in2 : std_logic_vector(1 downto 0);
    signal VN1772_in3 : std_logic_vector(1 downto 0);
    signal VN1772_in4 : std_logic_vector(1 downto 0);
    signal VN1772_in5 : std_logic_vector(1 downto 0);
    signal VN1773_in0 : std_logic_vector(1 downto 0);
    signal VN1773_in1 : std_logic_vector(1 downto 0);
    signal VN1773_in2 : std_logic_vector(1 downto 0);
    signal VN1773_in3 : std_logic_vector(1 downto 0);
    signal VN1773_in4 : std_logic_vector(1 downto 0);
    signal VN1773_in5 : std_logic_vector(1 downto 0);
    signal VN1774_in0 : std_logic_vector(1 downto 0);
    signal VN1774_in1 : std_logic_vector(1 downto 0);
    signal VN1774_in2 : std_logic_vector(1 downto 0);
    signal VN1774_in3 : std_logic_vector(1 downto 0);
    signal VN1774_in4 : std_logic_vector(1 downto 0);
    signal VN1774_in5 : std_logic_vector(1 downto 0);
    signal VN1775_in0 : std_logic_vector(1 downto 0);
    signal VN1775_in1 : std_logic_vector(1 downto 0);
    signal VN1775_in2 : std_logic_vector(1 downto 0);
    signal VN1775_in3 : std_logic_vector(1 downto 0);
    signal VN1775_in4 : std_logic_vector(1 downto 0);
    signal VN1775_in5 : std_logic_vector(1 downto 0);
    signal VN1776_in0 : std_logic_vector(1 downto 0);
    signal VN1776_in1 : std_logic_vector(1 downto 0);
    signal VN1776_in2 : std_logic_vector(1 downto 0);
    signal VN1776_in3 : std_logic_vector(1 downto 0);
    signal VN1776_in4 : std_logic_vector(1 downto 0);
    signal VN1776_in5 : std_logic_vector(1 downto 0);
    signal VN1777_in0 : std_logic_vector(1 downto 0);
    signal VN1777_in1 : std_logic_vector(1 downto 0);
    signal VN1777_in2 : std_logic_vector(1 downto 0);
    signal VN1777_in3 : std_logic_vector(1 downto 0);
    signal VN1777_in4 : std_logic_vector(1 downto 0);
    signal VN1777_in5 : std_logic_vector(1 downto 0);
    signal VN1778_in0 : std_logic_vector(1 downto 0);
    signal VN1778_in1 : std_logic_vector(1 downto 0);
    signal VN1778_in2 : std_logic_vector(1 downto 0);
    signal VN1778_in3 : std_logic_vector(1 downto 0);
    signal VN1778_in4 : std_logic_vector(1 downto 0);
    signal VN1778_in5 : std_logic_vector(1 downto 0);
    signal VN1779_in0 : std_logic_vector(1 downto 0);
    signal VN1779_in1 : std_logic_vector(1 downto 0);
    signal VN1779_in2 : std_logic_vector(1 downto 0);
    signal VN1779_in3 : std_logic_vector(1 downto 0);
    signal VN1779_in4 : std_logic_vector(1 downto 0);
    signal VN1779_in5 : std_logic_vector(1 downto 0);
    signal VN1780_in0 : std_logic_vector(1 downto 0);
    signal VN1780_in1 : std_logic_vector(1 downto 0);
    signal VN1780_in2 : std_logic_vector(1 downto 0);
    signal VN1780_in3 : std_logic_vector(1 downto 0);
    signal VN1780_in4 : std_logic_vector(1 downto 0);
    signal VN1780_in5 : std_logic_vector(1 downto 0);
    signal VN1781_in0 : std_logic_vector(1 downto 0);
    signal VN1781_in1 : std_logic_vector(1 downto 0);
    signal VN1781_in2 : std_logic_vector(1 downto 0);
    signal VN1781_in3 : std_logic_vector(1 downto 0);
    signal VN1781_in4 : std_logic_vector(1 downto 0);
    signal VN1781_in5 : std_logic_vector(1 downto 0);
    signal VN1782_in0 : std_logic_vector(1 downto 0);
    signal VN1782_in1 : std_logic_vector(1 downto 0);
    signal VN1782_in2 : std_logic_vector(1 downto 0);
    signal VN1782_in3 : std_logic_vector(1 downto 0);
    signal VN1782_in4 : std_logic_vector(1 downto 0);
    signal VN1782_in5 : std_logic_vector(1 downto 0);
    signal VN1783_in0 : std_logic_vector(1 downto 0);
    signal VN1783_in1 : std_logic_vector(1 downto 0);
    signal VN1783_in2 : std_logic_vector(1 downto 0);
    signal VN1783_in3 : std_logic_vector(1 downto 0);
    signal VN1783_in4 : std_logic_vector(1 downto 0);
    signal VN1783_in5 : std_logic_vector(1 downto 0);
    signal VN1784_in0 : std_logic_vector(1 downto 0);
    signal VN1784_in1 : std_logic_vector(1 downto 0);
    signal VN1784_in2 : std_logic_vector(1 downto 0);
    signal VN1784_in3 : std_logic_vector(1 downto 0);
    signal VN1784_in4 : std_logic_vector(1 downto 0);
    signal VN1784_in5 : std_logic_vector(1 downto 0);
    signal VN1785_in0 : std_logic_vector(1 downto 0);
    signal VN1785_in1 : std_logic_vector(1 downto 0);
    signal VN1785_in2 : std_logic_vector(1 downto 0);
    signal VN1785_in3 : std_logic_vector(1 downto 0);
    signal VN1785_in4 : std_logic_vector(1 downto 0);
    signal VN1785_in5 : std_logic_vector(1 downto 0);
    signal VN1786_in0 : std_logic_vector(1 downto 0);
    signal VN1786_in1 : std_logic_vector(1 downto 0);
    signal VN1786_in2 : std_logic_vector(1 downto 0);
    signal VN1786_in3 : std_logic_vector(1 downto 0);
    signal VN1786_in4 : std_logic_vector(1 downto 0);
    signal VN1786_in5 : std_logic_vector(1 downto 0);
    signal VN1787_in0 : std_logic_vector(1 downto 0);
    signal VN1787_in1 : std_logic_vector(1 downto 0);
    signal VN1787_in2 : std_logic_vector(1 downto 0);
    signal VN1787_in3 : std_logic_vector(1 downto 0);
    signal VN1787_in4 : std_logic_vector(1 downto 0);
    signal VN1787_in5 : std_logic_vector(1 downto 0);
    signal VN1788_in0 : std_logic_vector(1 downto 0);
    signal VN1788_in1 : std_logic_vector(1 downto 0);
    signal VN1788_in2 : std_logic_vector(1 downto 0);
    signal VN1788_in3 : std_logic_vector(1 downto 0);
    signal VN1788_in4 : std_logic_vector(1 downto 0);
    signal VN1788_in5 : std_logic_vector(1 downto 0);
    signal VN1789_in0 : std_logic_vector(1 downto 0);
    signal VN1789_in1 : std_logic_vector(1 downto 0);
    signal VN1789_in2 : std_logic_vector(1 downto 0);
    signal VN1789_in3 : std_logic_vector(1 downto 0);
    signal VN1789_in4 : std_logic_vector(1 downto 0);
    signal VN1789_in5 : std_logic_vector(1 downto 0);
    signal VN1790_in0 : std_logic_vector(1 downto 0);
    signal VN1790_in1 : std_logic_vector(1 downto 0);
    signal VN1790_in2 : std_logic_vector(1 downto 0);
    signal VN1790_in3 : std_logic_vector(1 downto 0);
    signal VN1790_in4 : std_logic_vector(1 downto 0);
    signal VN1790_in5 : std_logic_vector(1 downto 0);
    signal VN1791_in0 : std_logic_vector(1 downto 0);
    signal VN1791_in1 : std_logic_vector(1 downto 0);
    signal VN1791_in2 : std_logic_vector(1 downto 0);
    signal VN1791_in3 : std_logic_vector(1 downto 0);
    signal VN1791_in4 : std_logic_vector(1 downto 0);
    signal VN1791_in5 : std_logic_vector(1 downto 0);
    signal VN1792_in0 : std_logic_vector(1 downto 0);
    signal VN1792_in1 : std_logic_vector(1 downto 0);
    signal VN1792_in2 : std_logic_vector(1 downto 0);
    signal VN1792_in3 : std_logic_vector(1 downto 0);
    signal VN1792_in4 : std_logic_vector(1 downto 0);
    signal VN1792_in5 : std_logic_vector(1 downto 0);
    signal VN1793_in0 : std_logic_vector(1 downto 0);
    signal VN1793_in1 : std_logic_vector(1 downto 0);
    signal VN1793_in2 : std_logic_vector(1 downto 0);
    signal VN1793_in3 : std_logic_vector(1 downto 0);
    signal VN1793_in4 : std_logic_vector(1 downto 0);
    signal VN1793_in5 : std_logic_vector(1 downto 0);
    signal VN1794_in0 : std_logic_vector(1 downto 0);
    signal VN1794_in1 : std_logic_vector(1 downto 0);
    signal VN1794_in2 : std_logic_vector(1 downto 0);
    signal VN1794_in3 : std_logic_vector(1 downto 0);
    signal VN1794_in4 : std_logic_vector(1 downto 0);
    signal VN1794_in5 : std_logic_vector(1 downto 0);
    signal VN1795_in0 : std_logic_vector(1 downto 0);
    signal VN1795_in1 : std_logic_vector(1 downto 0);
    signal VN1795_in2 : std_logic_vector(1 downto 0);
    signal VN1795_in3 : std_logic_vector(1 downto 0);
    signal VN1795_in4 : std_logic_vector(1 downto 0);
    signal VN1795_in5 : std_logic_vector(1 downto 0);
    signal VN1796_in0 : std_logic_vector(1 downto 0);
    signal VN1796_in1 : std_logic_vector(1 downto 0);
    signal VN1796_in2 : std_logic_vector(1 downto 0);
    signal VN1796_in3 : std_logic_vector(1 downto 0);
    signal VN1796_in4 : std_logic_vector(1 downto 0);
    signal VN1796_in5 : std_logic_vector(1 downto 0);
    signal VN1797_in0 : std_logic_vector(1 downto 0);
    signal VN1797_in1 : std_logic_vector(1 downto 0);
    signal VN1797_in2 : std_logic_vector(1 downto 0);
    signal VN1797_in3 : std_logic_vector(1 downto 0);
    signal VN1797_in4 : std_logic_vector(1 downto 0);
    signal VN1797_in5 : std_logic_vector(1 downto 0);
    signal VN1798_in0 : std_logic_vector(1 downto 0);
    signal VN1798_in1 : std_logic_vector(1 downto 0);
    signal VN1798_in2 : std_logic_vector(1 downto 0);
    signal VN1798_in3 : std_logic_vector(1 downto 0);
    signal VN1798_in4 : std_logic_vector(1 downto 0);
    signal VN1798_in5 : std_logic_vector(1 downto 0);
    signal VN1799_in0 : std_logic_vector(1 downto 0);
    signal VN1799_in1 : std_logic_vector(1 downto 0);
    signal VN1799_in2 : std_logic_vector(1 downto 0);
    signal VN1799_in3 : std_logic_vector(1 downto 0);
    signal VN1799_in4 : std_logic_vector(1 downto 0);
    signal VN1799_in5 : std_logic_vector(1 downto 0);
    signal VN1800_in0 : std_logic_vector(1 downto 0);
    signal VN1800_in1 : std_logic_vector(1 downto 0);
    signal VN1800_in2 : std_logic_vector(1 downto 0);
    signal VN1800_in3 : std_logic_vector(1 downto 0);
    signal VN1800_in4 : std_logic_vector(1 downto 0);
    signal VN1800_in5 : std_logic_vector(1 downto 0);
    signal VN1801_in0 : std_logic_vector(1 downto 0);
    signal VN1801_in1 : std_logic_vector(1 downto 0);
    signal VN1801_in2 : std_logic_vector(1 downto 0);
    signal VN1801_in3 : std_logic_vector(1 downto 0);
    signal VN1801_in4 : std_logic_vector(1 downto 0);
    signal VN1801_in5 : std_logic_vector(1 downto 0);
    signal VN1802_in0 : std_logic_vector(1 downto 0);
    signal VN1802_in1 : std_logic_vector(1 downto 0);
    signal VN1802_in2 : std_logic_vector(1 downto 0);
    signal VN1802_in3 : std_logic_vector(1 downto 0);
    signal VN1802_in4 : std_logic_vector(1 downto 0);
    signal VN1802_in5 : std_logic_vector(1 downto 0);
    signal VN1803_in0 : std_logic_vector(1 downto 0);
    signal VN1803_in1 : std_logic_vector(1 downto 0);
    signal VN1803_in2 : std_logic_vector(1 downto 0);
    signal VN1803_in3 : std_logic_vector(1 downto 0);
    signal VN1803_in4 : std_logic_vector(1 downto 0);
    signal VN1803_in5 : std_logic_vector(1 downto 0);
    signal VN1804_in0 : std_logic_vector(1 downto 0);
    signal VN1804_in1 : std_logic_vector(1 downto 0);
    signal VN1804_in2 : std_logic_vector(1 downto 0);
    signal VN1804_in3 : std_logic_vector(1 downto 0);
    signal VN1804_in4 : std_logic_vector(1 downto 0);
    signal VN1804_in5 : std_logic_vector(1 downto 0);
    signal VN1805_in0 : std_logic_vector(1 downto 0);
    signal VN1805_in1 : std_logic_vector(1 downto 0);
    signal VN1805_in2 : std_logic_vector(1 downto 0);
    signal VN1805_in3 : std_logic_vector(1 downto 0);
    signal VN1805_in4 : std_logic_vector(1 downto 0);
    signal VN1805_in5 : std_logic_vector(1 downto 0);
    signal VN1806_in0 : std_logic_vector(1 downto 0);
    signal VN1806_in1 : std_logic_vector(1 downto 0);
    signal VN1806_in2 : std_logic_vector(1 downto 0);
    signal VN1806_in3 : std_logic_vector(1 downto 0);
    signal VN1806_in4 : std_logic_vector(1 downto 0);
    signal VN1806_in5 : std_logic_vector(1 downto 0);
    signal VN1807_in0 : std_logic_vector(1 downto 0);
    signal VN1807_in1 : std_logic_vector(1 downto 0);
    signal VN1807_in2 : std_logic_vector(1 downto 0);
    signal VN1807_in3 : std_logic_vector(1 downto 0);
    signal VN1807_in4 : std_logic_vector(1 downto 0);
    signal VN1807_in5 : std_logic_vector(1 downto 0);
    signal VN1808_in0 : std_logic_vector(1 downto 0);
    signal VN1808_in1 : std_logic_vector(1 downto 0);
    signal VN1808_in2 : std_logic_vector(1 downto 0);
    signal VN1808_in3 : std_logic_vector(1 downto 0);
    signal VN1808_in4 : std_logic_vector(1 downto 0);
    signal VN1808_in5 : std_logic_vector(1 downto 0);
    signal VN1809_in0 : std_logic_vector(1 downto 0);
    signal VN1809_in1 : std_logic_vector(1 downto 0);
    signal VN1809_in2 : std_logic_vector(1 downto 0);
    signal VN1809_in3 : std_logic_vector(1 downto 0);
    signal VN1809_in4 : std_logic_vector(1 downto 0);
    signal VN1809_in5 : std_logic_vector(1 downto 0);
    signal VN1810_in0 : std_logic_vector(1 downto 0);
    signal VN1810_in1 : std_logic_vector(1 downto 0);
    signal VN1810_in2 : std_logic_vector(1 downto 0);
    signal VN1810_in3 : std_logic_vector(1 downto 0);
    signal VN1810_in4 : std_logic_vector(1 downto 0);
    signal VN1810_in5 : std_logic_vector(1 downto 0);
    signal VN1811_in0 : std_logic_vector(1 downto 0);
    signal VN1811_in1 : std_logic_vector(1 downto 0);
    signal VN1811_in2 : std_logic_vector(1 downto 0);
    signal VN1811_in3 : std_logic_vector(1 downto 0);
    signal VN1811_in4 : std_logic_vector(1 downto 0);
    signal VN1811_in5 : std_logic_vector(1 downto 0);
    signal VN1812_in0 : std_logic_vector(1 downto 0);
    signal VN1812_in1 : std_logic_vector(1 downto 0);
    signal VN1812_in2 : std_logic_vector(1 downto 0);
    signal VN1812_in3 : std_logic_vector(1 downto 0);
    signal VN1812_in4 : std_logic_vector(1 downto 0);
    signal VN1812_in5 : std_logic_vector(1 downto 0);
    signal VN1813_in0 : std_logic_vector(1 downto 0);
    signal VN1813_in1 : std_logic_vector(1 downto 0);
    signal VN1813_in2 : std_logic_vector(1 downto 0);
    signal VN1813_in3 : std_logic_vector(1 downto 0);
    signal VN1813_in4 : std_logic_vector(1 downto 0);
    signal VN1813_in5 : std_logic_vector(1 downto 0);
    signal VN1814_in0 : std_logic_vector(1 downto 0);
    signal VN1814_in1 : std_logic_vector(1 downto 0);
    signal VN1814_in2 : std_logic_vector(1 downto 0);
    signal VN1814_in3 : std_logic_vector(1 downto 0);
    signal VN1814_in4 : std_logic_vector(1 downto 0);
    signal VN1814_in5 : std_logic_vector(1 downto 0);
    signal VN1815_in0 : std_logic_vector(1 downto 0);
    signal VN1815_in1 : std_logic_vector(1 downto 0);
    signal VN1815_in2 : std_logic_vector(1 downto 0);
    signal VN1815_in3 : std_logic_vector(1 downto 0);
    signal VN1815_in4 : std_logic_vector(1 downto 0);
    signal VN1815_in5 : std_logic_vector(1 downto 0);
    signal VN1816_in0 : std_logic_vector(1 downto 0);
    signal VN1816_in1 : std_logic_vector(1 downto 0);
    signal VN1816_in2 : std_logic_vector(1 downto 0);
    signal VN1816_in3 : std_logic_vector(1 downto 0);
    signal VN1816_in4 : std_logic_vector(1 downto 0);
    signal VN1816_in5 : std_logic_vector(1 downto 0);
    signal VN1817_in0 : std_logic_vector(1 downto 0);
    signal VN1817_in1 : std_logic_vector(1 downto 0);
    signal VN1817_in2 : std_logic_vector(1 downto 0);
    signal VN1817_in3 : std_logic_vector(1 downto 0);
    signal VN1817_in4 : std_logic_vector(1 downto 0);
    signal VN1817_in5 : std_logic_vector(1 downto 0);
    signal VN1818_in0 : std_logic_vector(1 downto 0);
    signal VN1818_in1 : std_logic_vector(1 downto 0);
    signal VN1818_in2 : std_logic_vector(1 downto 0);
    signal VN1818_in3 : std_logic_vector(1 downto 0);
    signal VN1818_in4 : std_logic_vector(1 downto 0);
    signal VN1818_in5 : std_logic_vector(1 downto 0);
    signal VN1819_in0 : std_logic_vector(1 downto 0);
    signal VN1819_in1 : std_logic_vector(1 downto 0);
    signal VN1819_in2 : std_logic_vector(1 downto 0);
    signal VN1819_in3 : std_logic_vector(1 downto 0);
    signal VN1819_in4 : std_logic_vector(1 downto 0);
    signal VN1819_in5 : std_logic_vector(1 downto 0);
    signal VN1820_in0 : std_logic_vector(1 downto 0);
    signal VN1820_in1 : std_logic_vector(1 downto 0);
    signal VN1820_in2 : std_logic_vector(1 downto 0);
    signal VN1820_in3 : std_logic_vector(1 downto 0);
    signal VN1820_in4 : std_logic_vector(1 downto 0);
    signal VN1820_in5 : std_logic_vector(1 downto 0);
    signal VN1821_in0 : std_logic_vector(1 downto 0);
    signal VN1821_in1 : std_logic_vector(1 downto 0);
    signal VN1821_in2 : std_logic_vector(1 downto 0);
    signal VN1821_in3 : std_logic_vector(1 downto 0);
    signal VN1821_in4 : std_logic_vector(1 downto 0);
    signal VN1821_in5 : std_logic_vector(1 downto 0);
    signal VN1822_in0 : std_logic_vector(1 downto 0);
    signal VN1822_in1 : std_logic_vector(1 downto 0);
    signal VN1822_in2 : std_logic_vector(1 downto 0);
    signal VN1822_in3 : std_logic_vector(1 downto 0);
    signal VN1822_in4 : std_logic_vector(1 downto 0);
    signal VN1822_in5 : std_logic_vector(1 downto 0);
    signal VN1823_in0 : std_logic_vector(1 downto 0);
    signal VN1823_in1 : std_logic_vector(1 downto 0);
    signal VN1823_in2 : std_logic_vector(1 downto 0);
    signal VN1823_in3 : std_logic_vector(1 downto 0);
    signal VN1823_in4 : std_logic_vector(1 downto 0);
    signal VN1823_in5 : std_logic_vector(1 downto 0);
    signal VN1824_in0 : std_logic_vector(1 downto 0);
    signal VN1824_in1 : std_logic_vector(1 downto 0);
    signal VN1824_in2 : std_logic_vector(1 downto 0);
    signal VN1824_in3 : std_logic_vector(1 downto 0);
    signal VN1824_in4 : std_logic_vector(1 downto 0);
    signal VN1824_in5 : std_logic_vector(1 downto 0);
    signal VN1825_in0 : std_logic_vector(1 downto 0);
    signal VN1825_in1 : std_logic_vector(1 downto 0);
    signal VN1825_in2 : std_logic_vector(1 downto 0);
    signal VN1825_in3 : std_logic_vector(1 downto 0);
    signal VN1825_in4 : std_logic_vector(1 downto 0);
    signal VN1825_in5 : std_logic_vector(1 downto 0);
    signal VN1826_in0 : std_logic_vector(1 downto 0);
    signal VN1826_in1 : std_logic_vector(1 downto 0);
    signal VN1826_in2 : std_logic_vector(1 downto 0);
    signal VN1826_in3 : std_logic_vector(1 downto 0);
    signal VN1826_in4 : std_logic_vector(1 downto 0);
    signal VN1826_in5 : std_logic_vector(1 downto 0);
    signal VN1827_in0 : std_logic_vector(1 downto 0);
    signal VN1827_in1 : std_logic_vector(1 downto 0);
    signal VN1827_in2 : std_logic_vector(1 downto 0);
    signal VN1827_in3 : std_logic_vector(1 downto 0);
    signal VN1827_in4 : std_logic_vector(1 downto 0);
    signal VN1827_in5 : std_logic_vector(1 downto 0);
    signal VN1828_in0 : std_logic_vector(1 downto 0);
    signal VN1828_in1 : std_logic_vector(1 downto 0);
    signal VN1828_in2 : std_logic_vector(1 downto 0);
    signal VN1828_in3 : std_logic_vector(1 downto 0);
    signal VN1828_in4 : std_logic_vector(1 downto 0);
    signal VN1828_in5 : std_logic_vector(1 downto 0);
    signal VN1829_in0 : std_logic_vector(1 downto 0);
    signal VN1829_in1 : std_logic_vector(1 downto 0);
    signal VN1829_in2 : std_logic_vector(1 downto 0);
    signal VN1829_in3 : std_logic_vector(1 downto 0);
    signal VN1829_in4 : std_logic_vector(1 downto 0);
    signal VN1829_in5 : std_logic_vector(1 downto 0);
    signal VN1830_in0 : std_logic_vector(1 downto 0);
    signal VN1830_in1 : std_logic_vector(1 downto 0);
    signal VN1830_in2 : std_logic_vector(1 downto 0);
    signal VN1830_in3 : std_logic_vector(1 downto 0);
    signal VN1830_in4 : std_logic_vector(1 downto 0);
    signal VN1830_in5 : std_logic_vector(1 downto 0);
    signal VN1831_in0 : std_logic_vector(1 downto 0);
    signal VN1831_in1 : std_logic_vector(1 downto 0);
    signal VN1831_in2 : std_logic_vector(1 downto 0);
    signal VN1831_in3 : std_logic_vector(1 downto 0);
    signal VN1831_in4 : std_logic_vector(1 downto 0);
    signal VN1831_in5 : std_logic_vector(1 downto 0);
    signal VN1832_in0 : std_logic_vector(1 downto 0);
    signal VN1832_in1 : std_logic_vector(1 downto 0);
    signal VN1832_in2 : std_logic_vector(1 downto 0);
    signal VN1832_in3 : std_logic_vector(1 downto 0);
    signal VN1832_in4 : std_logic_vector(1 downto 0);
    signal VN1832_in5 : std_logic_vector(1 downto 0);
    signal VN1833_in0 : std_logic_vector(1 downto 0);
    signal VN1833_in1 : std_logic_vector(1 downto 0);
    signal VN1833_in2 : std_logic_vector(1 downto 0);
    signal VN1833_in3 : std_logic_vector(1 downto 0);
    signal VN1833_in4 : std_logic_vector(1 downto 0);
    signal VN1833_in5 : std_logic_vector(1 downto 0);
    signal VN1834_in0 : std_logic_vector(1 downto 0);
    signal VN1834_in1 : std_logic_vector(1 downto 0);
    signal VN1834_in2 : std_logic_vector(1 downto 0);
    signal VN1834_in3 : std_logic_vector(1 downto 0);
    signal VN1834_in4 : std_logic_vector(1 downto 0);
    signal VN1834_in5 : std_logic_vector(1 downto 0);
    signal VN1835_in0 : std_logic_vector(1 downto 0);
    signal VN1835_in1 : std_logic_vector(1 downto 0);
    signal VN1835_in2 : std_logic_vector(1 downto 0);
    signal VN1835_in3 : std_logic_vector(1 downto 0);
    signal VN1835_in4 : std_logic_vector(1 downto 0);
    signal VN1835_in5 : std_logic_vector(1 downto 0);
    signal VN1836_in0 : std_logic_vector(1 downto 0);
    signal VN1836_in1 : std_logic_vector(1 downto 0);
    signal VN1836_in2 : std_logic_vector(1 downto 0);
    signal VN1836_in3 : std_logic_vector(1 downto 0);
    signal VN1836_in4 : std_logic_vector(1 downto 0);
    signal VN1836_in5 : std_logic_vector(1 downto 0);
    signal VN1837_in0 : std_logic_vector(1 downto 0);
    signal VN1837_in1 : std_logic_vector(1 downto 0);
    signal VN1837_in2 : std_logic_vector(1 downto 0);
    signal VN1837_in3 : std_logic_vector(1 downto 0);
    signal VN1837_in4 : std_logic_vector(1 downto 0);
    signal VN1837_in5 : std_logic_vector(1 downto 0);
    signal VN1838_in0 : std_logic_vector(1 downto 0);
    signal VN1838_in1 : std_logic_vector(1 downto 0);
    signal VN1838_in2 : std_logic_vector(1 downto 0);
    signal VN1838_in3 : std_logic_vector(1 downto 0);
    signal VN1838_in4 : std_logic_vector(1 downto 0);
    signal VN1838_in5 : std_logic_vector(1 downto 0);
    signal VN1839_in0 : std_logic_vector(1 downto 0);
    signal VN1839_in1 : std_logic_vector(1 downto 0);
    signal VN1839_in2 : std_logic_vector(1 downto 0);
    signal VN1839_in3 : std_logic_vector(1 downto 0);
    signal VN1839_in4 : std_logic_vector(1 downto 0);
    signal VN1839_in5 : std_logic_vector(1 downto 0);
    signal VN1840_in0 : std_logic_vector(1 downto 0);
    signal VN1840_in1 : std_logic_vector(1 downto 0);
    signal VN1840_in2 : std_logic_vector(1 downto 0);
    signal VN1840_in3 : std_logic_vector(1 downto 0);
    signal VN1840_in4 : std_logic_vector(1 downto 0);
    signal VN1840_in5 : std_logic_vector(1 downto 0);
    signal VN1841_in0 : std_logic_vector(1 downto 0);
    signal VN1841_in1 : std_logic_vector(1 downto 0);
    signal VN1841_in2 : std_logic_vector(1 downto 0);
    signal VN1841_in3 : std_logic_vector(1 downto 0);
    signal VN1841_in4 : std_logic_vector(1 downto 0);
    signal VN1841_in5 : std_logic_vector(1 downto 0);
    signal VN1842_in0 : std_logic_vector(1 downto 0);
    signal VN1842_in1 : std_logic_vector(1 downto 0);
    signal VN1842_in2 : std_logic_vector(1 downto 0);
    signal VN1842_in3 : std_logic_vector(1 downto 0);
    signal VN1842_in4 : std_logic_vector(1 downto 0);
    signal VN1842_in5 : std_logic_vector(1 downto 0);
    signal VN1843_in0 : std_logic_vector(1 downto 0);
    signal VN1843_in1 : std_logic_vector(1 downto 0);
    signal VN1843_in2 : std_logic_vector(1 downto 0);
    signal VN1843_in3 : std_logic_vector(1 downto 0);
    signal VN1843_in4 : std_logic_vector(1 downto 0);
    signal VN1843_in5 : std_logic_vector(1 downto 0);
    signal VN1844_in0 : std_logic_vector(1 downto 0);
    signal VN1844_in1 : std_logic_vector(1 downto 0);
    signal VN1844_in2 : std_logic_vector(1 downto 0);
    signal VN1844_in3 : std_logic_vector(1 downto 0);
    signal VN1844_in4 : std_logic_vector(1 downto 0);
    signal VN1844_in5 : std_logic_vector(1 downto 0);
    signal VN1845_in0 : std_logic_vector(1 downto 0);
    signal VN1845_in1 : std_logic_vector(1 downto 0);
    signal VN1845_in2 : std_logic_vector(1 downto 0);
    signal VN1845_in3 : std_logic_vector(1 downto 0);
    signal VN1845_in4 : std_logic_vector(1 downto 0);
    signal VN1845_in5 : std_logic_vector(1 downto 0);
    signal VN1846_in0 : std_logic_vector(1 downto 0);
    signal VN1846_in1 : std_logic_vector(1 downto 0);
    signal VN1846_in2 : std_logic_vector(1 downto 0);
    signal VN1846_in3 : std_logic_vector(1 downto 0);
    signal VN1846_in4 : std_logic_vector(1 downto 0);
    signal VN1846_in5 : std_logic_vector(1 downto 0);
    signal VN1847_in0 : std_logic_vector(1 downto 0);
    signal VN1847_in1 : std_logic_vector(1 downto 0);
    signal VN1847_in2 : std_logic_vector(1 downto 0);
    signal VN1847_in3 : std_logic_vector(1 downto 0);
    signal VN1847_in4 : std_logic_vector(1 downto 0);
    signal VN1847_in5 : std_logic_vector(1 downto 0);
    signal VN1848_in0 : std_logic_vector(1 downto 0);
    signal VN1848_in1 : std_logic_vector(1 downto 0);
    signal VN1848_in2 : std_logic_vector(1 downto 0);
    signal VN1848_in3 : std_logic_vector(1 downto 0);
    signal VN1848_in4 : std_logic_vector(1 downto 0);
    signal VN1848_in5 : std_logic_vector(1 downto 0);
    signal VN1849_in0 : std_logic_vector(1 downto 0);
    signal VN1849_in1 : std_logic_vector(1 downto 0);
    signal VN1849_in2 : std_logic_vector(1 downto 0);
    signal VN1849_in3 : std_logic_vector(1 downto 0);
    signal VN1849_in4 : std_logic_vector(1 downto 0);
    signal VN1849_in5 : std_logic_vector(1 downto 0);
    signal VN1850_in0 : std_logic_vector(1 downto 0);
    signal VN1850_in1 : std_logic_vector(1 downto 0);
    signal VN1850_in2 : std_logic_vector(1 downto 0);
    signal VN1850_in3 : std_logic_vector(1 downto 0);
    signal VN1850_in4 : std_logic_vector(1 downto 0);
    signal VN1850_in5 : std_logic_vector(1 downto 0);
    signal VN1851_in0 : std_logic_vector(1 downto 0);
    signal VN1851_in1 : std_logic_vector(1 downto 0);
    signal VN1851_in2 : std_logic_vector(1 downto 0);
    signal VN1851_in3 : std_logic_vector(1 downto 0);
    signal VN1851_in4 : std_logic_vector(1 downto 0);
    signal VN1851_in5 : std_logic_vector(1 downto 0);
    signal VN1852_in0 : std_logic_vector(1 downto 0);
    signal VN1852_in1 : std_logic_vector(1 downto 0);
    signal VN1852_in2 : std_logic_vector(1 downto 0);
    signal VN1852_in3 : std_logic_vector(1 downto 0);
    signal VN1852_in4 : std_logic_vector(1 downto 0);
    signal VN1852_in5 : std_logic_vector(1 downto 0);
    signal VN1853_in0 : std_logic_vector(1 downto 0);
    signal VN1853_in1 : std_logic_vector(1 downto 0);
    signal VN1853_in2 : std_logic_vector(1 downto 0);
    signal VN1853_in3 : std_logic_vector(1 downto 0);
    signal VN1853_in4 : std_logic_vector(1 downto 0);
    signal VN1853_in5 : std_logic_vector(1 downto 0);
    signal VN1854_in0 : std_logic_vector(1 downto 0);
    signal VN1854_in1 : std_logic_vector(1 downto 0);
    signal VN1854_in2 : std_logic_vector(1 downto 0);
    signal VN1854_in3 : std_logic_vector(1 downto 0);
    signal VN1854_in4 : std_logic_vector(1 downto 0);
    signal VN1854_in5 : std_logic_vector(1 downto 0);
    signal VN1855_in0 : std_logic_vector(1 downto 0);
    signal VN1855_in1 : std_logic_vector(1 downto 0);
    signal VN1855_in2 : std_logic_vector(1 downto 0);
    signal VN1855_in3 : std_logic_vector(1 downto 0);
    signal VN1855_in4 : std_logic_vector(1 downto 0);
    signal VN1855_in5 : std_logic_vector(1 downto 0);
    signal VN1856_in0 : std_logic_vector(1 downto 0);
    signal VN1856_in1 : std_logic_vector(1 downto 0);
    signal VN1856_in2 : std_logic_vector(1 downto 0);
    signal VN1856_in3 : std_logic_vector(1 downto 0);
    signal VN1856_in4 : std_logic_vector(1 downto 0);
    signal VN1856_in5 : std_logic_vector(1 downto 0);
    signal VN1857_in0 : std_logic_vector(1 downto 0);
    signal VN1857_in1 : std_logic_vector(1 downto 0);
    signal VN1857_in2 : std_logic_vector(1 downto 0);
    signal VN1857_in3 : std_logic_vector(1 downto 0);
    signal VN1857_in4 : std_logic_vector(1 downto 0);
    signal VN1857_in5 : std_logic_vector(1 downto 0);
    signal VN1858_in0 : std_logic_vector(1 downto 0);
    signal VN1858_in1 : std_logic_vector(1 downto 0);
    signal VN1858_in2 : std_logic_vector(1 downto 0);
    signal VN1858_in3 : std_logic_vector(1 downto 0);
    signal VN1858_in4 : std_logic_vector(1 downto 0);
    signal VN1858_in5 : std_logic_vector(1 downto 0);
    signal VN1859_in0 : std_logic_vector(1 downto 0);
    signal VN1859_in1 : std_logic_vector(1 downto 0);
    signal VN1859_in2 : std_logic_vector(1 downto 0);
    signal VN1859_in3 : std_logic_vector(1 downto 0);
    signal VN1859_in4 : std_logic_vector(1 downto 0);
    signal VN1859_in5 : std_logic_vector(1 downto 0);
    signal VN1860_in0 : std_logic_vector(1 downto 0);
    signal VN1860_in1 : std_logic_vector(1 downto 0);
    signal VN1860_in2 : std_logic_vector(1 downto 0);
    signal VN1860_in3 : std_logic_vector(1 downto 0);
    signal VN1860_in4 : std_logic_vector(1 downto 0);
    signal VN1860_in5 : std_logic_vector(1 downto 0);
    signal VN1861_in0 : std_logic_vector(1 downto 0);
    signal VN1861_in1 : std_logic_vector(1 downto 0);
    signal VN1861_in2 : std_logic_vector(1 downto 0);
    signal VN1861_in3 : std_logic_vector(1 downto 0);
    signal VN1861_in4 : std_logic_vector(1 downto 0);
    signal VN1861_in5 : std_logic_vector(1 downto 0);
    signal VN1862_in0 : std_logic_vector(1 downto 0);
    signal VN1862_in1 : std_logic_vector(1 downto 0);
    signal VN1862_in2 : std_logic_vector(1 downto 0);
    signal VN1862_in3 : std_logic_vector(1 downto 0);
    signal VN1862_in4 : std_logic_vector(1 downto 0);
    signal VN1862_in5 : std_logic_vector(1 downto 0);
    signal VN1863_in0 : std_logic_vector(1 downto 0);
    signal VN1863_in1 : std_logic_vector(1 downto 0);
    signal VN1863_in2 : std_logic_vector(1 downto 0);
    signal VN1863_in3 : std_logic_vector(1 downto 0);
    signal VN1863_in4 : std_logic_vector(1 downto 0);
    signal VN1863_in5 : std_logic_vector(1 downto 0);
    signal VN1864_in0 : std_logic_vector(1 downto 0);
    signal VN1864_in1 : std_logic_vector(1 downto 0);
    signal VN1864_in2 : std_logic_vector(1 downto 0);
    signal VN1864_in3 : std_logic_vector(1 downto 0);
    signal VN1864_in4 : std_logic_vector(1 downto 0);
    signal VN1864_in5 : std_logic_vector(1 downto 0);
    signal VN1865_in0 : std_logic_vector(1 downto 0);
    signal VN1865_in1 : std_logic_vector(1 downto 0);
    signal VN1865_in2 : std_logic_vector(1 downto 0);
    signal VN1865_in3 : std_logic_vector(1 downto 0);
    signal VN1865_in4 : std_logic_vector(1 downto 0);
    signal VN1865_in5 : std_logic_vector(1 downto 0);
    signal VN1866_in0 : std_logic_vector(1 downto 0);
    signal VN1866_in1 : std_logic_vector(1 downto 0);
    signal VN1866_in2 : std_logic_vector(1 downto 0);
    signal VN1866_in3 : std_logic_vector(1 downto 0);
    signal VN1866_in4 : std_logic_vector(1 downto 0);
    signal VN1866_in5 : std_logic_vector(1 downto 0);
    signal VN1867_in0 : std_logic_vector(1 downto 0);
    signal VN1867_in1 : std_logic_vector(1 downto 0);
    signal VN1867_in2 : std_logic_vector(1 downto 0);
    signal VN1867_in3 : std_logic_vector(1 downto 0);
    signal VN1867_in4 : std_logic_vector(1 downto 0);
    signal VN1867_in5 : std_logic_vector(1 downto 0);
    signal VN1868_in0 : std_logic_vector(1 downto 0);
    signal VN1868_in1 : std_logic_vector(1 downto 0);
    signal VN1868_in2 : std_logic_vector(1 downto 0);
    signal VN1868_in3 : std_logic_vector(1 downto 0);
    signal VN1868_in4 : std_logic_vector(1 downto 0);
    signal VN1868_in5 : std_logic_vector(1 downto 0);
    signal VN1869_in0 : std_logic_vector(1 downto 0);
    signal VN1869_in1 : std_logic_vector(1 downto 0);
    signal VN1869_in2 : std_logic_vector(1 downto 0);
    signal VN1869_in3 : std_logic_vector(1 downto 0);
    signal VN1869_in4 : std_logic_vector(1 downto 0);
    signal VN1869_in5 : std_logic_vector(1 downto 0);
    signal VN1870_in0 : std_logic_vector(1 downto 0);
    signal VN1870_in1 : std_logic_vector(1 downto 0);
    signal VN1870_in2 : std_logic_vector(1 downto 0);
    signal VN1870_in3 : std_logic_vector(1 downto 0);
    signal VN1870_in4 : std_logic_vector(1 downto 0);
    signal VN1870_in5 : std_logic_vector(1 downto 0);
    signal VN1871_in0 : std_logic_vector(1 downto 0);
    signal VN1871_in1 : std_logic_vector(1 downto 0);
    signal VN1871_in2 : std_logic_vector(1 downto 0);
    signal VN1871_in3 : std_logic_vector(1 downto 0);
    signal VN1871_in4 : std_logic_vector(1 downto 0);
    signal VN1871_in5 : std_logic_vector(1 downto 0);
    signal VN1872_in0 : std_logic_vector(1 downto 0);
    signal VN1872_in1 : std_logic_vector(1 downto 0);
    signal VN1872_in2 : std_logic_vector(1 downto 0);
    signal VN1872_in3 : std_logic_vector(1 downto 0);
    signal VN1872_in4 : std_logic_vector(1 downto 0);
    signal VN1872_in5 : std_logic_vector(1 downto 0);
    signal VN1873_in0 : std_logic_vector(1 downto 0);
    signal VN1873_in1 : std_logic_vector(1 downto 0);
    signal VN1873_in2 : std_logic_vector(1 downto 0);
    signal VN1873_in3 : std_logic_vector(1 downto 0);
    signal VN1873_in4 : std_logic_vector(1 downto 0);
    signal VN1873_in5 : std_logic_vector(1 downto 0);
    signal VN1874_in0 : std_logic_vector(1 downto 0);
    signal VN1874_in1 : std_logic_vector(1 downto 0);
    signal VN1874_in2 : std_logic_vector(1 downto 0);
    signal VN1874_in3 : std_logic_vector(1 downto 0);
    signal VN1874_in4 : std_logic_vector(1 downto 0);
    signal VN1874_in5 : std_logic_vector(1 downto 0);
    signal VN1875_in0 : std_logic_vector(1 downto 0);
    signal VN1875_in1 : std_logic_vector(1 downto 0);
    signal VN1875_in2 : std_logic_vector(1 downto 0);
    signal VN1875_in3 : std_logic_vector(1 downto 0);
    signal VN1875_in4 : std_logic_vector(1 downto 0);
    signal VN1875_in5 : std_logic_vector(1 downto 0);
    signal VN1876_in0 : std_logic_vector(1 downto 0);
    signal VN1876_in1 : std_logic_vector(1 downto 0);
    signal VN1876_in2 : std_logic_vector(1 downto 0);
    signal VN1876_in3 : std_logic_vector(1 downto 0);
    signal VN1876_in4 : std_logic_vector(1 downto 0);
    signal VN1876_in5 : std_logic_vector(1 downto 0);
    signal VN1877_in0 : std_logic_vector(1 downto 0);
    signal VN1877_in1 : std_logic_vector(1 downto 0);
    signal VN1877_in2 : std_logic_vector(1 downto 0);
    signal VN1877_in3 : std_logic_vector(1 downto 0);
    signal VN1877_in4 : std_logic_vector(1 downto 0);
    signal VN1877_in5 : std_logic_vector(1 downto 0);
    signal VN1878_in0 : std_logic_vector(1 downto 0);
    signal VN1878_in1 : std_logic_vector(1 downto 0);
    signal VN1878_in2 : std_logic_vector(1 downto 0);
    signal VN1878_in3 : std_logic_vector(1 downto 0);
    signal VN1878_in4 : std_logic_vector(1 downto 0);
    signal VN1878_in5 : std_logic_vector(1 downto 0);
    signal VN1879_in0 : std_logic_vector(1 downto 0);
    signal VN1879_in1 : std_logic_vector(1 downto 0);
    signal VN1879_in2 : std_logic_vector(1 downto 0);
    signal VN1879_in3 : std_logic_vector(1 downto 0);
    signal VN1879_in4 : std_logic_vector(1 downto 0);
    signal VN1879_in5 : std_logic_vector(1 downto 0);
    signal VN1880_in0 : std_logic_vector(1 downto 0);
    signal VN1880_in1 : std_logic_vector(1 downto 0);
    signal VN1880_in2 : std_logic_vector(1 downto 0);
    signal VN1880_in3 : std_logic_vector(1 downto 0);
    signal VN1880_in4 : std_logic_vector(1 downto 0);
    signal VN1880_in5 : std_logic_vector(1 downto 0);
    signal VN1881_in0 : std_logic_vector(1 downto 0);
    signal VN1881_in1 : std_logic_vector(1 downto 0);
    signal VN1881_in2 : std_logic_vector(1 downto 0);
    signal VN1881_in3 : std_logic_vector(1 downto 0);
    signal VN1881_in4 : std_logic_vector(1 downto 0);
    signal VN1881_in5 : std_logic_vector(1 downto 0);
    signal VN1882_in0 : std_logic_vector(1 downto 0);
    signal VN1882_in1 : std_logic_vector(1 downto 0);
    signal VN1882_in2 : std_logic_vector(1 downto 0);
    signal VN1882_in3 : std_logic_vector(1 downto 0);
    signal VN1882_in4 : std_logic_vector(1 downto 0);
    signal VN1882_in5 : std_logic_vector(1 downto 0);
    signal VN1883_in0 : std_logic_vector(1 downto 0);
    signal VN1883_in1 : std_logic_vector(1 downto 0);
    signal VN1883_in2 : std_logic_vector(1 downto 0);
    signal VN1883_in3 : std_logic_vector(1 downto 0);
    signal VN1883_in4 : std_logic_vector(1 downto 0);
    signal VN1883_in5 : std_logic_vector(1 downto 0);
    signal VN1884_in0 : std_logic_vector(1 downto 0);
    signal VN1884_in1 : std_logic_vector(1 downto 0);
    signal VN1884_in2 : std_logic_vector(1 downto 0);
    signal VN1884_in3 : std_logic_vector(1 downto 0);
    signal VN1884_in4 : std_logic_vector(1 downto 0);
    signal VN1884_in5 : std_logic_vector(1 downto 0);
    signal VN1885_in0 : std_logic_vector(1 downto 0);
    signal VN1885_in1 : std_logic_vector(1 downto 0);
    signal VN1885_in2 : std_logic_vector(1 downto 0);
    signal VN1885_in3 : std_logic_vector(1 downto 0);
    signal VN1885_in4 : std_logic_vector(1 downto 0);
    signal VN1885_in5 : std_logic_vector(1 downto 0);
    signal VN1886_in0 : std_logic_vector(1 downto 0);
    signal VN1886_in1 : std_logic_vector(1 downto 0);
    signal VN1886_in2 : std_logic_vector(1 downto 0);
    signal VN1886_in3 : std_logic_vector(1 downto 0);
    signal VN1886_in4 : std_logic_vector(1 downto 0);
    signal VN1886_in5 : std_logic_vector(1 downto 0);
    signal VN1887_in0 : std_logic_vector(1 downto 0);
    signal VN1887_in1 : std_logic_vector(1 downto 0);
    signal VN1887_in2 : std_logic_vector(1 downto 0);
    signal VN1887_in3 : std_logic_vector(1 downto 0);
    signal VN1887_in4 : std_logic_vector(1 downto 0);
    signal VN1887_in5 : std_logic_vector(1 downto 0);
    signal VN1888_in0 : std_logic_vector(1 downto 0);
    signal VN1888_in1 : std_logic_vector(1 downto 0);
    signal VN1888_in2 : std_logic_vector(1 downto 0);
    signal VN1888_in3 : std_logic_vector(1 downto 0);
    signal VN1888_in4 : std_logic_vector(1 downto 0);
    signal VN1888_in5 : std_logic_vector(1 downto 0);
    signal VN1889_in0 : std_logic_vector(1 downto 0);
    signal VN1889_in1 : std_logic_vector(1 downto 0);
    signal VN1889_in2 : std_logic_vector(1 downto 0);
    signal VN1889_in3 : std_logic_vector(1 downto 0);
    signal VN1889_in4 : std_logic_vector(1 downto 0);
    signal VN1889_in5 : std_logic_vector(1 downto 0);
    signal VN1890_in0 : std_logic_vector(1 downto 0);
    signal VN1890_in1 : std_logic_vector(1 downto 0);
    signal VN1890_in2 : std_logic_vector(1 downto 0);
    signal VN1890_in3 : std_logic_vector(1 downto 0);
    signal VN1890_in4 : std_logic_vector(1 downto 0);
    signal VN1890_in5 : std_logic_vector(1 downto 0);
    signal VN1891_in0 : std_logic_vector(1 downto 0);
    signal VN1891_in1 : std_logic_vector(1 downto 0);
    signal VN1891_in2 : std_logic_vector(1 downto 0);
    signal VN1891_in3 : std_logic_vector(1 downto 0);
    signal VN1891_in4 : std_logic_vector(1 downto 0);
    signal VN1891_in5 : std_logic_vector(1 downto 0);
    signal VN1892_in0 : std_logic_vector(1 downto 0);
    signal VN1892_in1 : std_logic_vector(1 downto 0);
    signal VN1892_in2 : std_logic_vector(1 downto 0);
    signal VN1892_in3 : std_logic_vector(1 downto 0);
    signal VN1892_in4 : std_logic_vector(1 downto 0);
    signal VN1892_in5 : std_logic_vector(1 downto 0);
    signal VN1893_in0 : std_logic_vector(1 downto 0);
    signal VN1893_in1 : std_logic_vector(1 downto 0);
    signal VN1893_in2 : std_logic_vector(1 downto 0);
    signal VN1893_in3 : std_logic_vector(1 downto 0);
    signal VN1893_in4 : std_logic_vector(1 downto 0);
    signal VN1893_in5 : std_logic_vector(1 downto 0);
    signal VN1894_in0 : std_logic_vector(1 downto 0);
    signal VN1894_in1 : std_logic_vector(1 downto 0);
    signal VN1894_in2 : std_logic_vector(1 downto 0);
    signal VN1894_in3 : std_logic_vector(1 downto 0);
    signal VN1894_in4 : std_logic_vector(1 downto 0);
    signal VN1894_in5 : std_logic_vector(1 downto 0);
    signal VN1895_in0 : std_logic_vector(1 downto 0);
    signal VN1895_in1 : std_logic_vector(1 downto 0);
    signal VN1895_in2 : std_logic_vector(1 downto 0);
    signal VN1895_in3 : std_logic_vector(1 downto 0);
    signal VN1895_in4 : std_logic_vector(1 downto 0);
    signal VN1895_in5 : std_logic_vector(1 downto 0);
    signal VN1896_in0 : std_logic_vector(1 downto 0);
    signal VN1896_in1 : std_logic_vector(1 downto 0);
    signal VN1896_in2 : std_logic_vector(1 downto 0);
    signal VN1896_in3 : std_logic_vector(1 downto 0);
    signal VN1896_in4 : std_logic_vector(1 downto 0);
    signal VN1896_in5 : std_logic_vector(1 downto 0);
    signal VN1897_in0 : std_logic_vector(1 downto 0);
    signal VN1897_in1 : std_logic_vector(1 downto 0);
    signal VN1897_in2 : std_logic_vector(1 downto 0);
    signal VN1897_in3 : std_logic_vector(1 downto 0);
    signal VN1897_in4 : std_logic_vector(1 downto 0);
    signal VN1897_in5 : std_logic_vector(1 downto 0);
    signal VN1898_in0 : std_logic_vector(1 downto 0);
    signal VN1898_in1 : std_logic_vector(1 downto 0);
    signal VN1898_in2 : std_logic_vector(1 downto 0);
    signal VN1898_in3 : std_logic_vector(1 downto 0);
    signal VN1898_in4 : std_logic_vector(1 downto 0);
    signal VN1898_in5 : std_logic_vector(1 downto 0);
    signal VN1899_in0 : std_logic_vector(1 downto 0);
    signal VN1899_in1 : std_logic_vector(1 downto 0);
    signal VN1899_in2 : std_logic_vector(1 downto 0);
    signal VN1899_in3 : std_logic_vector(1 downto 0);
    signal VN1899_in4 : std_logic_vector(1 downto 0);
    signal VN1899_in5 : std_logic_vector(1 downto 0);
    signal VN1900_in0 : std_logic_vector(1 downto 0);
    signal VN1900_in1 : std_logic_vector(1 downto 0);
    signal VN1900_in2 : std_logic_vector(1 downto 0);
    signal VN1900_in3 : std_logic_vector(1 downto 0);
    signal VN1900_in4 : std_logic_vector(1 downto 0);
    signal VN1900_in5 : std_logic_vector(1 downto 0);
    signal VN1901_in0 : std_logic_vector(1 downto 0);
    signal VN1901_in1 : std_logic_vector(1 downto 0);
    signal VN1901_in2 : std_logic_vector(1 downto 0);
    signal VN1901_in3 : std_logic_vector(1 downto 0);
    signal VN1901_in4 : std_logic_vector(1 downto 0);
    signal VN1901_in5 : std_logic_vector(1 downto 0);
    signal VN1902_in0 : std_logic_vector(1 downto 0);
    signal VN1902_in1 : std_logic_vector(1 downto 0);
    signal VN1902_in2 : std_logic_vector(1 downto 0);
    signal VN1902_in3 : std_logic_vector(1 downto 0);
    signal VN1902_in4 : std_logic_vector(1 downto 0);
    signal VN1902_in5 : std_logic_vector(1 downto 0);
    signal VN1903_in0 : std_logic_vector(1 downto 0);
    signal VN1903_in1 : std_logic_vector(1 downto 0);
    signal VN1903_in2 : std_logic_vector(1 downto 0);
    signal VN1903_in3 : std_logic_vector(1 downto 0);
    signal VN1903_in4 : std_logic_vector(1 downto 0);
    signal VN1903_in5 : std_logic_vector(1 downto 0);
    signal VN1904_in0 : std_logic_vector(1 downto 0);
    signal VN1904_in1 : std_logic_vector(1 downto 0);
    signal VN1904_in2 : std_logic_vector(1 downto 0);
    signal VN1904_in3 : std_logic_vector(1 downto 0);
    signal VN1904_in4 : std_logic_vector(1 downto 0);
    signal VN1904_in5 : std_logic_vector(1 downto 0);
    signal VN1905_in0 : std_logic_vector(1 downto 0);
    signal VN1905_in1 : std_logic_vector(1 downto 0);
    signal VN1905_in2 : std_logic_vector(1 downto 0);
    signal VN1905_in3 : std_logic_vector(1 downto 0);
    signal VN1905_in4 : std_logic_vector(1 downto 0);
    signal VN1905_in5 : std_logic_vector(1 downto 0);
    signal VN1906_in0 : std_logic_vector(1 downto 0);
    signal VN1906_in1 : std_logic_vector(1 downto 0);
    signal VN1906_in2 : std_logic_vector(1 downto 0);
    signal VN1906_in3 : std_logic_vector(1 downto 0);
    signal VN1906_in4 : std_logic_vector(1 downto 0);
    signal VN1906_in5 : std_logic_vector(1 downto 0);
    signal VN1907_in0 : std_logic_vector(1 downto 0);
    signal VN1907_in1 : std_logic_vector(1 downto 0);
    signal VN1907_in2 : std_logic_vector(1 downto 0);
    signal VN1907_in3 : std_logic_vector(1 downto 0);
    signal VN1907_in4 : std_logic_vector(1 downto 0);
    signal VN1907_in5 : std_logic_vector(1 downto 0);
    signal VN1908_in0 : std_logic_vector(1 downto 0);
    signal VN1908_in1 : std_logic_vector(1 downto 0);
    signal VN1908_in2 : std_logic_vector(1 downto 0);
    signal VN1908_in3 : std_logic_vector(1 downto 0);
    signal VN1908_in4 : std_logic_vector(1 downto 0);
    signal VN1908_in5 : std_logic_vector(1 downto 0);
    signal VN1909_in0 : std_logic_vector(1 downto 0);
    signal VN1909_in1 : std_logic_vector(1 downto 0);
    signal VN1909_in2 : std_logic_vector(1 downto 0);
    signal VN1909_in3 : std_logic_vector(1 downto 0);
    signal VN1909_in4 : std_logic_vector(1 downto 0);
    signal VN1909_in5 : std_logic_vector(1 downto 0);
    signal VN1910_in0 : std_logic_vector(1 downto 0);
    signal VN1910_in1 : std_logic_vector(1 downto 0);
    signal VN1910_in2 : std_logic_vector(1 downto 0);
    signal VN1910_in3 : std_logic_vector(1 downto 0);
    signal VN1910_in4 : std_logic_vector(1 downto 0);
    signal VN1910_in5 : std_logic_vector(1 downto 0);
    signal VN1911_in0 : std_logic_vector(1 downto 0);
    signal VN1911_in1 : std_logic_vector(1 downto 0);
    signal VN1911_in2 : std_logic_vector(1 downto 0);
    signal VN1911_in3 : std_logic_vector(1 downto 0);
    signal VN1911_in4 : std_logic_vector(1 downto 0);
    signal VN1911_in5 : std_logic_vector(1 downto 0);
    signal VN1912_in0 : std_logic_vector(1 downto 0);
    signal VN1912_in1 : std_logic_vector(1 downto 0);
    signal VN1912_in2 : std_logic_vector(1 downto 0);
    signal VN1912_in3 : std_logic_vector(1 downto 0);
    signal VN1912_in4 : std_logic_vector(1 downto 0);
    signal VN1912_in5 : std_logic_vector(1 downto 0);
    signal VN1913_in0 : std_logic_vector(1 downto 0);
    signal VN1913_in1 : std_logic_vector(1 downto 0);
    signal VN1913_in2 : std_logic_vector(1 downto 0);
    signal VN1913_in3 : std_logic_vector(1 downto 0);
    signal VN1913_in4 : std_logic_vector(1 downto 0);
    signal VN1913_in5 : std_logic_vector(1 downto 0);
    signal VN1914_in0 : std_logic_vector(1 downto 0);
    signal VN1914_in1 : std_logic_vector(1 downto 0);
    signal VN1914_in2 : std_logic_vector(1 downto 0);
    signal VN1914_in3 : std_logic_vector(1 downto 0);
    signal VN1914_in4 : std_logic_vector(1 downto 0);
    signal VN1914_in5 : std_logic_vector(1 downto 0);
    signal VN1915_in0 : std_logic_vector(1 downto 0);
    signal VN1915_in1 : std_logic_vector(1 downto 0);
    signal VN1915_in2 : std_logic_vector(1 downto 0);
    signal VN1915_in3 : std_logic_vector(1 downto 0);
    signal VN1915_in4 : std_logic_vector(1 downto 0);
    signal VN1915_in5 : std_logic_vector(1 downto 0);
    signal VN1916_in0 : std_logic_vector(1 downto 0);
    signal VN1916_in1 : std_logic_vector(1 downto 0);
    signal VN1916_in2 : std_logic_vector(1 downto 0);
    signal VN1916_in3 : std_logic_vector(1 downto 0);
    signal VN1916_in4 : std_logic_vector(1 downto 0);
    signal VN1916_in5 : std_logic_vector(1 downto 0);
    signal VN1917_in0 : std_logic_vector(1 downto 0);
    signal VN1917_in1 : std_logic_vector(1 downto 0);
    signal VN1917_in2 : std_logic_vector(1 downto 0);
    signal VN1917_in3 : std_logic_vector(1 downto 0);
    signal VN1917_in4 : std_logic_vector(1 downto 0);
    signal VN1917_in5 : std_logic_vector(1 downto 0);
    signal VN1918_in0 : std_logic_vector(1 downto 0);
    signal VN1918_in1 : std_logic_vector(1 downto 0);
    signal VN1918_in2 : std_logic_vector(1 downto 0);
    signal VN1918_in3 : std_logic_vector(1 downto 0);
    signal VN1918_in4 : std_logic_vector(1 downto 0);
    signal VN1918_in5 : std_logic_vector(1 downto 0);
    signal VN1919_in0 : std_logic_vector(1 downto 0);
    signal VN1919_in1 : std_logic_vector(1 downto 0);
    signal VN1919_in2 : std_logic_vector(1 downto 0);
    signal VN1919_in3 : std_logic_vector(1 downto 0);
    signal VN1919_in4 : std_logic_vector(1 downto 0);
    signal VN1919_in5 : std_logic_vector(1 downto 0);
    signal VN1920_in0 : std_logic_vector(1 downto 0);
    signal VN1920_in1 : std_logic_vector(1 downto 0);
    signal VN1920_in2 : std_logic_vector(1 downto 0);
    signal VN1920_in3 : std_logic_vector(1 downto 0);
    signal VN1920_in4 : std_logic_vector(1 downto 0);
    signal VN1920_in5 : std_logic_vector(1 downto 0);
    signal VN1921_in0 : std_logic_vector(1 downto 0);
    signal VN1921_in1 : std_logic_vector(1 downto 0);
    signal VN1921_in2 : std_logic_vector(1 downto 0);
    signal VN1921_in3 : std_logic_vector(1 downto 0);
    signal VN1921_in4 : std_logic_vector(1 downto 0);
    signal VN1921_in5 : std_logic_vector(1 downto 0);
    signal VN1922_in0 : std_logic_vector(1 downto 0);
    signal VN1922_in1 : std_logic_vector(1 downto 0);
    signal VN1922_in2 : std_logic_vector(1 downto 0);
    signal VN1922_in3 : std_logic_vector(1 downto 0);
    signal VN1922_in4 : std_logic_vector(1 downto 0);
    signal VN1922_in5 : std_logic_vector(1 downto 0);
    signal VN1923_in0 : std_logic_vector(1 downto 0);
    signal VN1923_in1 : std_logic_vector(1 downto 0);
    signal VN1923_in2 : std_logic_vector(1 downto 0);
    signal VN1923_in3 : std_logic_vector(1 downto 0);
    signal VN1923_in4 : std_logic_vector(1 downto 0);
    signal VN1923_in5 : std_logic_vector(1 downto 0);
    signal VN1924_in0 : std_logic_vector(1 downto 0);
    signal VN1924_in1 : std_logic_vector(1 downto 0);
    signal VN1924_in2 : std_logic_vector(1 downto 0);
    signal VN1924_in3 : std_logic_vector(1 downto 0);
    signal VN1924_in4 : std_logic_vector(1 downto 0);
    signal VN1924_in5 : std_logic_vector(1 downto 0);
    signal VN1925_in0 : std_logic_vector(1 downto 0);
    signal VN1925_in1 : std_logic_vector(1 downto 0);
    signal VN1925_in2 : std_logic_vector(1 downto 0);
    signal VN1925_in3 : std_logic_vector(1 downto 0);
    signal VN1925_in4 : std_logic_vector(1 downto 0);
    signal VN1925_in5 : std_logic_vector(1 downto 0);
    signal VN1926_in0 : std_logic_vector(1 downto 0);
    signal VN1926_in1 : std_logic_vector(1 downto 0);
    signal VN1926_in2 : std_logic_vector(1 downto 0);
    signal VN1926_in3 : std_logic_vector(1 downto 0);
    signal VN1926_in4 : std_logic_vector(1 downto 0);
    signal VN1926_in5 : std_logic_vector(1 downto 0);
    signal VN1927_in0 : std_logic_vector(1 downto 0);
    signal VN1927_in1 : std_logic_vector(1 downto 0);
    signal VN1927_in2 : std_logic_vector(1 downto 0);
    signal VN1927_in3 : std_logic_vector(1 downto 0);
    signal VN1927_in4 : std_logic_vector(1 downto 0);
    signal VN1927_in5 : std_logic_vector(1 downto 0);
    signal VN1928_in0 : std_logic_vector(1 downto 0);
    signal VN1928_in1 : std_logic_vector(1 downto 0);
    signal VN1928_in2 : std_logic_vector(1 downto 0);
    signal VN1928_in3 : std_logic_vector(1 downto 0);
    signal VN1928_in4 : std_logic_vector(1 downto 0);
    signal VN1928_in5 : std_logic_vector(1 downto 0);
    signal VN1929_in0 : std_logic_vector(1 downto 0);
    signal VN1929_in1 : std_logic_vector(1 downto 0);
    signal VN1929_in2 : std_logic_vector(1 downto 0);
    signal VN1929_in3 : std_logic_vector(1 downto 0);
    signal VN1929_in4 : std_logic_vector(1 downto 0);
    signal VN1929_in5 : std_logic_vector(1 downto 0);
    signal VN1930_in0 : std_logic_vector(1 downto 0);
    signal VN1930_in1 : std_logic_vector(1 downto 0);
    signal VN1930_in2 : std_logic_vector(1 downto 0);
    signal VN1930_in3 : std_logic_vector(1 downto 0);
    signal VN1930_in4 : std_logic_vector(1 downto 0);
    signal VN1930_in5 : std_logic_vector(1 downto 0);
    signal VN1931_in0 : std_logic_vector(1 downto 0);
    signal VN1931_in1 : std_logic_vector(1 downto 0);
    signal VN1931_in2 : std_logic_vector(1 downto 0);
    signal VN1931_in3 : std_logic_vector(1 downto 0);
    signal VN1931_in4 : std_logic_vector(1 downto 0);
    signal VN1931_in5 : std_logic_vector(1 downto 0);
    signal VN1932_in0 : std_logic_vector(1 downto 0);
    signal VN1932_in1 : std_logic_vector(1 downto 0);
    signal VN1932_in2 : std_logic_vector(1 downto 0);
    signal VN1932_in3 : std_logic_vector(1 downto 0);
    signal VN1932_in4 : std_logic_vector(1 downto 0);
    signal VN1932_in5 : std_logic_vector(1 downto 0);
    signal VN1933_in0 : std_logic_vector(1 downto 0);
    signal VN1933_in1 : std_logic_vector(1 downto 0);
    signal VN1933_in2 : std_logic_vector(1 downto 0);
    signal VN1933_in3 : std_logic_vector(1 downto 0);
    signal VN1933_in4 : std_logic_vector(1 downto 0);
    signal VN1933_in5 : std_logic_vector(1 downto 0);
    signal VN1934_in0 : std_logic_vector(1 downto 0);
    signal VN1934_in1 : std_logic_vector(1 downto 0);
    signal VN1934_in2 : std_logic_vector(1 downto 0);
    signal VN1934_in3 : std_logic_vector(1 downto 0);
    signal VN1934_in4 : std_logic_vector(1 downto 0);
    signal VN1934_in5 : std_logic_vector(1 downto 0);
    signal VN1935_in0 : std_logic_vector(1 downto 0);
    signal VN1935_in1 : std_logic_vector(1 downto 0);
    signal VN1935_in2 : std_logic_vector(1 downto 0);
    signal VN1935_in3 : std_logic_vector(1 downto 0);
    signal VN1935_in4 : std_logic_vector(1 downto 0);
    signal VN1935_in5 : std_logic_vector(1 downto 0);
    signal VN1936_in0 : std_logic_vector(1 downto 0);
    signal VN1936_in1 : std_logic_vector(1 downto 0);
    signal VN1936_in2 : std_logic_vector(1 downto 0);
    signal VN1936_in3 : std_logic_vector(1 downto 0);
    signal VN1936_in4 : std_logic_vector(1 downto 0);
    signal VN1936_in5 : std_logic_vector(1 downto 0);
    signal VN1937_in0 : std_logic_vector(1 downto 0);
    signal VN1937_in1 : std_logic_vector(1 downto 0);
    signal VN1937_in2 : std_logic_vector(1 downto 0);
    signal VN1937_in3 : std_logic_vector(1 downto 0);
    signal VN1937_in4 : std_logic_vector(1 downto 0);
    signal VN1937_in5 : std_logic_vector(1 downto 0);
    signal VN1938_in0 : std_logic_vector(1 downto 0);
    signal VN1938_in1 : std_logic_vector(1 downto 0);
    signal VN1938_in2 : std_logic_vector(1 downto 0);
    signal VN1938_in3 : std_logic_vector(1 downto 0);
    signal VN1938_in4 : std_logic_vector(1 downto 0);
    signal VN1938_in5 : std_logic_vector(1 downto 0);
    signal VN1939_in0 : std_logic_vector(1 downto 0);
    signal VN1939_in1 : std_logic_vector(1 downto 0);
    signal VN1939_in2 : std_logic_vector(1 downto 0);
    signal VN1939_in3 : std_logic_vector(1 downto 0);
    signal VN1939_in4 : std_logic_vector(1 downto 0);
    signal VN1939_in5 : std_logic_vector(1 downto 0);
    signal VN1940_in0 : std_logic_vector(1 downto 0);
    signal VN1940_in1 : std_logic_vector(1 downto 0);
    signal VN1940_in2 : std_logic_vector(1 downto 0);
    signal VN1940_in3 : std_logic_vector(1 downto 0);
    signal VN1940_in4 : std_logic_vector(1 downto 0);
    signal VN1940_in5 : std_logic_vector(1 downto 0);
    signal VN1941_in0 : std_logic_vector(1 downto 0);
    signal VN1941_in1 : std_logic_vector(1 downto 0);
    signal VN1941_in2 : std_logic_vector(1 downto 0);
    signal VN1941_in3 : std_logic_vector(1 downto 0);
    signal VN1941_in4 : std_logic_vector(1 downto 0);
    signal VN1941_in5 : std_logic_vector(1 downto 0);
    signal VN1942_in0 : std_logic_vector(1 downto 0);
    signal VN1942_in1 : std_logic_vector(1 downto 0);
    signal VN1942_in2 : std_logic_vector(1 downto 0);
    signal VN1942_in3 : std_logic_vector(1 downto 0);
    signal VN1942_in4 : std_logic_vector(1 downto 0);
    signal VN1942_in5 : std_logic_vector(1 downto 0);
    signal VN1943_in0 : std_logic_vector(1 downto 0);
    signal VN1943_in1 : std_logic_vector(1 downto 0);
    signal VN1943_in2 : std_logic_vector(1 downto 0);
    signal VN1943_in3 : std_logic_vector(1 downto 0);
    signal VN1943_in4 : std_logic_vector(1 downto 0);
    signal VN1943_in5 : std_logic_vector(1 downto 0);
    signal VN1944_in0 : std_logic_vector(1 downto 0);
    signal VN1944_in1 : std_logic_vector(1 downto 0);
    signal VN1944_in2 : std_logic_vector(1 downto 0);
    signal VN1944_in3 : std_logic_vector(1 downto 0);
    signal VN1944_in4 : std_logic_vector(1 downto 0);
    signal VN1944_in5 : std_logic_vector(1 downto 0);
    signal VN1945_in0 : std_logic_vector(1 downto 0);
    signal VN1945_in1 : std_logic_vector(1 downto 0);
    signal VN1945_in2 : std_logic_vector(1 downto 0);
    signal VN1945_in3 : std_logic_vector(1 downto 0);
    signal VN1945_in4 : std_logic_vector(1 downto 0);
    signal VN1945_in5 : std_logic_vector(1 downto 0);
    signal VN1946_in0 : std_logic_vector(1 downto 0);
    signal VN1946_in1 : std_logic_vector(1 downto 0);
    signal VN1946_in2 : std_logic_vector(1 downto 0);
    signal VN1946_in3 : std_logic_vector(1 downto 0);
    signal VN1946_in4 : std_logic_vector(1 downto 0);
    signal VN1946_in5 : std_logic_vector(1 downto 0);
    signal VN1947_in0 : std_logic_vector(1 downto 0);
    signal VN1947_in1 : std_logic_vector(1 downto 0);
    signal VN1947_in2 : std_logic_vector(1 downto 0);
    signal VN1947_in3 : std_logic_vector(1 downto 0);
    signal VN1947_in4 : std_logic_vector(1 downto 0);
    signal VN1947_in5 : std_logic_vector(1 downto 0);
    signal VN1948_in0 : std_logic_vector(1 downto 0);
    signal VN1948_in1 : std_logic_vector(1 downto 0);
    signal VN1948_in2 : std_logic_vector(1 downto 0);
    signal VN1948_in3 : std_logic_vector(1 downto 0);
    signal VN1948_in4 : std_logic_vector(1 downto 0);
    signal VN1948_in5 : std_logic_vector(1 downto 0);
    signal VN1949_in0 : std_logic_vector(1 downto 0);
    signal VN1949_in1 : std_logic_vector(1 downto 0);
    signal VN1949_in2 : std_logic_vector(1 downto 0);
    signal VN1949_in3 : std_logic_vector(1 downto 0);
    signal VN1949_in4 : std_logic_vector(1 downto 0);
    signal VN1949_in5 : std_logic_vector(1 downto 0);
    signal VN1950_in0 : std_logic_vector(1 downto 0);
    signal VN1950_in1 : std_logic_vector(1 downto 0);
    signal VN1950_in2 : std_logic_vector(1 downto 0);
    signal VN1950_in3 : std_logic_vector(1 downto 0);
    signal VN1950_in4 : std_logic_vector(1 downto 0);
    signal VN1950_in5 : std_logic_vector(1 downto 0);
    signal VN1951_in0 : std_logic_vector(1 downto 0);
    signal VN1951_in1 : std_logic_vector(1 downto 0);
    signal VN1951_in2 : std_logic_vector(1 downto 0);
    signal VN1951_in3 : std_logic_vector(1 downto 0);
    signal VN1951_in4 : std_logic_vector(1 downto 0);
    signal VN1951_in5 : std_logic_vector(1 downto 0);
    signal VN1952_in0 : std_logic_vector(1 downto 0);
    signal VN1952_in1 : std_logic_vector(1 downto 0);
    signal VN1952_in2 : std_logic_vector(1 downto 0);
    signal VN1952_in3 : std_logic_vector(1 downto 0);
    signal VN1952_in4 : std_logic_vector(1 downto 0);
    signal VN1952_in5 : std_logic_vector(1 downto 0);
    signal VN1953_in0 : std_logic_vector(1 downto 0);
    signal VN1953_in1 : std_logic_vector(1 downto 0);
    signal VN1953_in2 : std_logic_vector(1 downto 0);
    signal VN1953_in3 : std_logic_vector(1 downto 0);
    signal VN1953_in4 : std_logic_vector(1 downto 0);
    signal VN1953_in5 : std_logic_vector(1 downto 0);
    signal VN1954_in0 : std_logic_vector(1 downto 0);
    signal VN1954_in1 : std_logic_vector(1 downto 0);
    signal VN1954_in2 : std_logic_vector(1 downto 0);
    signal VN1954_in3 : std_logic_vector(1 downto 0);
    signal VN1954_in4 : std_logic_vector(1 downto 0);
    signal VN1954_in5 : std_logic_vector(1 downto 0);
    signal VN1955_in0 : std_logic_vector(1 downto 0);
    signal VN1955_in1 : std_logic_vector(1 downto 0);
    signal VN1955_in2 : std_logic_vector(1 downto 0);
    signal VN1955_in3 : std_logic_vector(1 downto 0);
    signal VN1955_in4 : std_logic_vector(1 downto 0);
    signal VN1955_in5 : std_logic_vector(1 downto 0);
    signal VN1956_in0 : std_logic_vector(1 downto 0);
    signal VN1956_in1 : std_logic_vector(1 downto 0);
    signal VN1956_in2 : std_logic_vector(1 downto 0);
    signal VN1956_in3 : std_logic_vector(1 downto 0);
    signal VN1956_in4 : std_logic_vector(1 downto 0);
    signal VN1956_in5 : std_logic_vector(1 downto 0);
    signal VN1957_in0 : std_logic_vector(1 downto 0);
    signal VN1957_in1 : std_logic_vector(1 downto 0);
    signal VN1957_in2 : std_logic_vector(1 downto 0);
    signal VN1957_in3 : std_logic_vector(1 downto 0);
    signal VN1957_in4 : std_logic_vector(1 downto 0);
    signal VN1957_in5 : std_logic_vector(1 downto 0);
    signal VN1958_in0 : std_logic_vector(1 downto 0);
    signal VN1958_in1 : std_logic_vector(1 downto 0);
    signal VN1958_in2 : std_logic_vector(1 downto 0);
    signal VN1958_in3 : std_logic_vector(1 downto 0);
    signal VN1958_in4 : std_logic_vector(1 downto 0);
    signal VN1958_in5 : std_logic_vector(1 downto 0);
    signal VN1959_in0 : std_logic_vector(1 downto 0);
    signal VN1959_in1 : std_logic_vector(1 downto 0);
    signal VN1959_in2 : std_logic_vector(1 downto 0);
    signal VN1959_in3 : std_logic_vector(1 downto 0);
    signal VN1959_in4 : std_logic_vector(1 downto 0);
    signal VN1959_in5 : std_logic_vector(1 downto 0);
    signal VN1960_in0 : std_logic_vector(1 downto 0);
    signal VN1960_in1 : std_logic_vector(1 downto 0);
    signal VN1960_in2 : std_logic_vector(1 downto 0);
    signal VN1960_in3 : std_logic_vector(1 downto 0);
    signal VN1960_in4 : std_logic_vector(1 downto 0);
    signal VN1960_in5 : std_logic_vector(1 downto 0);
    signal VN1961_in0 : std_logic_vector(1 downto 0);
    signal VN1961_in1 : std_logic_vector(1 downto 0);
    signal VN1961_in2 : std_logic_vector(1 downto 0);
    signal VN1961_in3 : std_logic_vector(1 downto 0);
    signal VN1961_in4 : std_logic_vector(1 downto 0);
    signal VN1961_in5 : std_logic_vector(1 downto 0);
    signal VN1962_in0 : std_logic_vector(1 downto 0);
    signal VN1962_in1 : std_logic_vector(1 downto 0);
    signal VN1962_in2 : std_logic_vector(1 downto 0);
    signal VN1962_in3 : std_logic_vector(1 downto 0);
    signal VN1962_in4 : std_logic_vector(1 downto 0);
    signal VN1962_in5 : std_logic_vector(1 downto 0);
    signal VN1963_in0 : std_logic_vector(1 downto 0);
    signal VN1963_in1 : std_logic_vector(1 downto 0);
    signal VN1963_in2 : std_logic_vector(1 downto 0);
    signal VN1963_in3 : std_logic_vector(1 downto 0);
    signal VN1963_in4 : std_logic_vector(1 downto 0);
    signal VN1963_in5 : std_logic_vector(1 downto 0);
    signal VN1964_in0 : std_logic_vector(1 downto 0);
    signal VN1964_in1 : std_logic_vector(1 downto 0);
    signal VN1964_in2 : std_logic_vector(1 downto 0);
    signal VN1964_in3 : std_logic_vector(1 downto 0);
    signal VN1964_in4 : std_logic_vector(1 downto 0);
    signal VN1964_in5 : std_logic_vector(1 downto 0);
    signal VN1965_in0 : std_logic_vector(1 downto 0);
    signal VN1965_in1 : std_logic_vector(1 downto 0);
    signal VN1965_in2 : std_logic_vector(1 downto 0);
    signal VN1965_in3 : std_logic_vector(1 downto 0);
    signal VN1965_in4 : std_logic_vector(1 downto 0);
    signal VN1965_in5 : std_logic_vector(1 downto 0);
    signal VN1966_in0 : std_logic_vector(1 downto 0);
    signal VN1966_in1 : std_logic_vector(1 downto 0);
    signal VN1966_in2 : std_logic_vector(1 downto 0);
    signal VN1966_in3 : std_logic_vector(1 downto 0);
    signal VN1966_in4 : std_logic_vector(1 downto 0);
    signal VN1966_in5 : std_logic_vector(1 downto 0);
    signal VN1967_in0 : std_logic_vector(1 downto 0);
    signal VN1967_in1 : std_logic_vector(1 downto 0);
    signal VN1967_in2 : std_logic_vector(1 downto 0);
    signal VN1967_in3 : std_logic_vector(1 downto 0);
    signal VN1967_in4 : std_logic_vector(1 downto 0);
    signal VN1967_in5 : std_logic_vector(1 downto 0);
    signal VN1968_in0 : std_logic_vector(1 downto 0);
    signal VN1968_in1 : std_logic_vector(1 downto 0);
    signal VN1968_in2 : std_logic_vector(1 downto 0);
    signal VN1968_in3 : std_logic_vector(1 downto 0);
    signal VN1968_in4 : std_logic_vector(1 downto 0);
    signal VN1968_in5 : std_logic_vector(1 downto 0);
    signal VN1969_in0 : std_logic_vector(1 downto 0);
    signal VN1969_in1 : std_logic_vector(1 downto 0);
    signal VN1969_in2 : std_logic_vector(1 downto 0);
    signal VN1969_in3 : std_logic_vector(1 downto 0);
    signal VN1969_in4 : std_logic_vector(1 downto 0);
    signal VN1969_in5 : std_logic_vector(1 downto 0);
    signal VN1970_in0 : std_logic_vector(1 downto 0);
    signal VN1970_in1 : std_logic_vector(1 downto 0);
    signal VN1970_in2 : std_logic_vector(1 downto 0);
    signal VN1970_in3 : std_logic_vector(1 downto 0);
    signal VN1970_in4 : std_logic_vector(1 downto 0);
    signal VN1970_in5 : std_logic_vector(1 downto 0);
    signal VN1971_in0 : std_logic_vector(1 downto 0);
    signal VN1971_in1 : std_logic_vector(1 downto 0);
    signal VN1971_in2 : std_logic_vector(1 downto 0);
    signal VN1971_in3 : std_logic_vector(1 downto 0);
    signal VN1971_in4 : std_logic_vector(1 downto 0);
    signal VN1971_in5 : std_logic_vector(1 downto 0);
    signal VN1972_in0 : std_logic_vector(1 downto 0);
    signal VN1972_in1 : std_logic_vector(1 downto 0);
    signal VN1972_in2 : std_logic_vector(1 downto 0);
    signal VN1972_in3 : std_logic_vector(1 downto 0);
    signal VN1972_in4 : std_logic_vector(1 downto 0);
    signal VN1972_in5 : std_logic_vector(1 downto 0);
    signal VN1973_in0 : std_logic_vector(1 downto 0);
    signal VN1973_in1 : std_logic_vector(1 downto 0);
    signal VN1973_in2 : std_logic_vector(1 downto 0);
    signal VN1973_in3 : std_logic_vector(1 downto 0);
    signal VN1973_in4 : std_logic_vector(1 downto 0);
    signal VN1973_in5 : std_logic_vector(1 downto 0);
    signal VN1974_in0 : std_logic_vector(1 downto 0);
    signal VN1974_in1 : std_logic_vector(1 downto 0);
    signal VN1974_in2 : std_logic_vector(1 downto 0);
    signal VN1974_in3 : std_logic_vector(1 downto 0);
    signal VN1974_in4 : std_logic_vector(1 downto 0);
    signal VN1974_in5 : std_logic_vector(1 downto 0);
    signal VN1975_in0 : std_logic_vector(1 downto 0);
    signal VN1975_in1 : std_logic_vector(1 downto 0);
    signal VN1975_in2 : std_logic_vector(1 downto 0);
    signal VN1975_in3 : std_logic_vector(1 downto 0);
    signal VN1975_in4 : std_logic_vector(1 downto 0);
    signal VN1975_in5 : std_logic_vector(1 downto 0);
    signal VN1976_in0 : std_logic_vector(1 downto 0);
    signal VN1976_in1 : std_logic_vector(1 downto 0);
    signal VN1976_in2 : std_logic_vector(1 downto 0);
    signal VN1976_in3 : std_logic_vector(1 downto 0);
    signal VN1976_in4 : std_logic_vector(1 downto 0);
    signal VN1976_in5 : std_logic_vector(1 downto 0);
    signal VN1977_in0 : std_logic_vector(1 downto 0);
    signal VN1977_in1 : std_logic_vector(1 downto 0);
    signal VN1977_in2 : std_logic_vector(1 downto 0);
    signal VN1977_in3 : std_logic_vector(1 downto 0);
    signal VN1977_in4 : std_logic_vector(1 downto 0);
    signal VN1977_in5 : std_logic_vector(1 downto 0);
    signal VN1978_in0 : std_logic_vector(1 downto 0);
    signal VN1978_in1 : std_logic_vector(1 downto 0);
    signal VN1978_in2 : std_logic_vector(1 downto 0);
    signal VN1978_in3 : std_logic_vector(1 downto 0);
    signal VN1978_in4 : std_logic_vector(1 downto 0);
    signal VN1978_in5 : std_logic_vector(1 downto 0);
    signal VN1979_in0 : std_logic_vector(1 downto 0);
    signal VN1979_in1 : std_logic_vector(1 downto 0);
    signal VN1979_in2 : std_logic_vector(1 downto 0);
    signal VN1979_in3 : std_logic_vector(1 downto 0);
    signal VN1979_in4 : std_logic_vector(1 downto 0);
    signal VN1979_in5 : std_logic_vector(1 downto 0);
    signal VN1980_in0 : std_logic_vector(1 downto 0);
    signal VN1980_in1 : std_logic_vector(1 downto 0);
    signal VN1980_in2 : std_logic_vector(1 downto 0);
    signal VN1980_in3 : std_logic_vector(1 downto 0);
    signal VN1980_in4 : std_logic_vector(1 downto 0);
    signal VN1980_in5 : std_logic_vector(1 downto 0);
    signal VN1981_in0 : std_logic_vector(1 downto 0);
    signal VN1981_in1 : std_logic_vector(1 downto 0);
    signal VN1981_in2 : std_logic_vector(1 downto 0);
    signal VN1981_in3 : std_logic_vector(1 downto 0);
    signal VN1981_in4 : std_logic_vector(1 downto 0);
    signal VN1981_in5 : std_logic_vector(1 downto 0);
    signal VN1982_in0 : std_logic_vector(1 downto 0);
    signal VN1982_in1 : std_logic_vector(1 downto 0);
    signal VN1982_in2 : std_logic_vector(1 downto 0);
    signal VN1982_in3 : std_logic_vector(1 downto 0);
    signal VN1982_in4 : std_logic_vector(1 downto 0);
    signal VN1982_in5 : std_logic_vector(1 downto 0);
    signal VN1983_in0 : std_logic_vector(1 downto 0);
    signal VN1983_in1 : std_logic_vector(1 downto 0);
    signal VN1983_in2 : std_logic_vector(1 downto 0);
    signal VN1983_in3 : std_logic_vector(1 downto 0);
    signal VN1983_in4 : std_logic_vector(1 downto 0);
    signal VN1983_in5 : std_logic_vector(1 downto 0);
    signal VN1984_in0 : std_logic_vector(1 downto 0);
    signal VN1984_in1 : std_logic_vector(1 downto 0);
    signal VN1984_in2 : std_logic_vector(1 downto 0);
    signal VN1984_in3 : std_logic_vector(1 downto 0);
    signal VN1984_in4 : std_logic_vector(1 downto 0);
    signal VN1984_in5 : std_logic_vector(1 downto 0);
    signal VN1985_in0 : std_logic_vector(1 downto 0);
    signal VN1985_in1 : std_logic_vector(1 downto 0);
    signal VN1985_in2 : std_logic_vector(1 downto 0);
    signal VN1985_in3 : std_logic_vector(1 downto 0);
    signal VN1985_in4 : std_logic_vector(1 downto 0);
    signal VN1985_in5 : std_logic_vector(1 downto 0);
    signal VN1986_in0 : std_logic_vector(1 downto 0);
    signal VN1986_in1 : std_logic_vector(1 downto 0);
    signal VN1986_in2 : std_logic_vector(1 downto 0);
    signal VN1986_in3 : std_logic_vector(1 downto 0);
    signal VN1986_in4 : std_logic_vector(1 downto 0);
    signal VN1986_in5 : std_logic_vector(1 downto 0);
    signal VN1987_in0 : std_logic_vector(1 downto 0);
    signal VN1987_in1 : std_logic_vector(1 downto 0);
    signal VN1987_in2 : std_logic_vector(1 downto 0);
    signal VN1987_in3 : std_logic_vector(1 downto 0);
    signal VN1987_in4 : std_logic_vector(1 downto 0);
    signal VN1987_in5 : std_logic_vector(1 downto 0);
    signal VN1988_in0 : std_logic_vector(1 downto 0);
    signal VN1988_in1 : std_logic_vector(1 downto 0);
    signal VN1988_in2 : std_logic_vector(1 downto 0);
    signal VN1988_in3 : std_logic_vector(1 downto 0);
    signal VN1988_in4 : std_logic_vector(1 downto 0);
    signal VN1988_in5 : std_logic_vector(1 downto 0);
    signal VN1989_in0 : std_logic_vector(1 downto 0);
    signal VN1989_in1 : std_logic_vector(1 downto 0);
    signal VN1989_in2 : std_logic_vector(1 downto 0);
    signal VN1989_in3 : std_logic_vector(1 downto 0);
    signal VN1989_in4 : std_logic_vector(1 downto 0);
    signal VN1989_in5 : std_logic_vector(1 downto 0);
    signal VN1990_in0 : std_logic_vector(1 downto 0);
    signal VN1990_in1 : std_logic_vector(1 downto 0);
    signal VN1990_in2 : std_logic_vector(1 downto 0);
    signal VN1990_in3 : std_logic_vector(1 downto 0);
    signal VN1990_in4 : std_logic_vector(1 downto 0);
    signal VN1990_in5 : std_logic_vector(1 downto 0);
    signal VN1991_in0 : std_logic_vector(1 downto 0);
    signal VN1991_in1 : std_logic_vector(1 downto 0);
    signal VN1991_in2 : std_logic_vector(1 downto 0);
    signal VN1991_in3 : std_logic_vector(1 downto 0);
    signal VN1991_in4 : std_logic_vector(1 downto 0);
    signal VN1991_in5 : std_logic_vector(1 downto 0);
    signal VN1992_in0 : std_logic_vector(1 downto 0);
    signal VN1992_in1 : std_logic_vector(1 downto 0);
    signal VN1992_in2 : std_logic_vector(1 downto 0);
    signal VN1992_in3 : std_logic_vector(1 downto 0);
    signal VN1992_in4 : std_logic_vector(1 downto 0);
    signal VN1992_in5 : std_logic_vector(1 downto 0);
    signal VN1993_in0 : std_logic_vector(1 downto 0);
    signal VN1993_in1 : std_logic_vector(1 downto 0);
    signal VN1993_in2 : std_logic_vector(1 downto 0);
    signal VN1993_in3 : std_logic_vector(1 downto 0);
    signal VN1993_in4 : std_logic_vector(1 downto 0);
    signal VN1993_in5 : std_logic_vector(1 downto 0);
    signal VN1994_in0 : std_logic_vector(1 downto 0);
    signal VN1994_in1 : std_logic_vector(1 downto 0);
    signal VN1994_in2 : std_logic_vector(1 downto 0);
    signal VN1994_in3 : std_logic_vector(1 downto 0);
    signal VN1994_in4 : std_logic_vector(1 downto 0);
    signal VN1994_in5 : std_logic_vector(1 downto 0);
    signal VN1995_in0 : std_logic_vector(1 downto 0);
    signal VN1995_in1 : std_logic_vector(1 downto 0);
    signal VN1995_in2 : std_logic_vector(1 downto 0);
    signal VN1995_in3 : std_logic_vector(1 downto 0);
    signal VN1995_in4 : std_logic_vector(1 downto 0);
    signal VN1995_in5 : std_logic_vector(1 downto 0);
    signal VN1996_in0 : std_logic_vector(1 downto 0);
    signal VN1996_in1 : std_logic_vector(1 downto 0);
    signal VN1996_in2 : std_logic_vector(1 downto 0);
    signal VN1996_in3 : std_logic_vector(1 downto 0);
    signal VN1996_in4 : std_logic_vector(1 downto 0);
    signal VN1996_in5 : std_logic_vector(1 downto 0);
    signal VN1997_in0 : std_logic_vector(1 downto 0);
    signal VN1997_in1 : std_logic_vector(1 downto 0);
    signal VN1997_in2 : std_logic_vector(1 downto 0);
    signal VN1997_in3 : std_logic_vector(1 downto 0);
    signal VN1997_in4 : std_logic_vector(1 downto 0);
    signal VN1997_in5 : std_logic_vector(1 downto 0);
    signal VN1998_in0 : std_logic_vector(1 downto 0);
    signal VN1998_in1 : std_logic_vector(1 downto 0);
    signal VN1998_in2 : std_logic_vector(1 downto 0);
    signal VN1998_in3 : std_logic_vector(1 downto 0);
    signal VN1998_in4 : std_logic_vector(1 downto 0);
    signal VN1998_in5 : std_logic_vector(1 downto 0);
    signal VN1999_in0 : std_logic_vector(1 downto 0);
    signal VN1999_in1 : std_logic_vector(1 downto 0);
    signal VN1999_in2 : std_logic_vector(1 downto 0);
    signal VN1999_in3 : std_logic_vector(1 downto 0);
    signal VN1999_in4 : std_logic_vector(1 downto 0);
    signal VN1999_in5 : std_logic_vector(1 downto 0);
    signal VN2000_in0 : std_logic_vector(1 downto 0);
    signal VN2000_in1 : std_logic_vector(1 downto 0);
    signal VN2000_in2 : std_logic_vector(1 downto 0);
    signal VN2000_in3 : std_logic_vector(1 downto 0);
    signal VN2000_in4 : std_logic_vector(1 downto 0);
    signal VN2000_in5 : std_logic_vector(1 downto 0);
    signal VN2001_in0 : std_logic_vector(1 downto 0);
    signal VN2001_in1 : std_logic_vector(1 downto 0);
    signal VN2001_in2 : std_logic_vector(1 downto 0);
    signal VN2001_in3 : std_logic_vector(1 downto 0);
    signal VN2001_in4 : std_logic_vector(1 downto 0);
    signal VN2001_in5 : std_logic_vector(1 downto 0);
    signal VN2002_in0 : std_logic_vector(1 downto 0);
    signal VN2002_in1 : std_logic_vector(1 downto 0);
    signal VN2002_in2 : std_logic_vector(1 downto 0);
    signal VN2002_in3 : std_logic_vector(1 downto 0);
    signal VN2002_in4 : std_logic_vector(1 downto 0);
    signal VN2002_in5 : std_logic_vector(1 downto 0);
    signal VN2003_in0 : std_logic_vector(1 downto 0);
    signal VN2003_in1 : std_logic_vector(1 downto 0);
    signal VN2003_in2 : std_logic_vector(1 downto 0);
    signal VN2003_in3 : std_logic_vector(1 downto 0);
    signal VN2003_in4 : std_logic_vector(1 downto 0);
    signal VN2003_in5 : std_logic_vector(1 downto 0);
    signal VN2004_in0 : std_logic_vector(1 downto 0);
    signal VN2004_in1 : std_logic_vector(1 downto 0);
    signal VN2004_in2 : std_logic_vector(1 downto 0);
    signal VN2004_in3 : std_logic_vector(1 downto 0);
    signal VN2004_in4 : std_logic_vector(1 downto 0);
    signal VN2004_in5 : std_logic_vector(1 downto 0);
    signal VN2005_in0 : std_logic_vector(1 downto 0);
    signal VN2005_in1 : std_logic_vector(1 downto 0);
    signal VN2005_in2 : std_logic_vector(1 downto 0);
    signal VN2005_in3 : std_logic_vector(1 downto 0);
    signal VN2005_in4 : std_logic_vector(1 downto 0);
    signal VN2005_in5 : std_logic_vector(1 downto 0);
    signal VN2006_in0 : std_logic_vector(1 downto 0);
    signal VN2006_in1 : std_logic_vector(1 downto 0);
    signal VN2006_in2 : std_logic_vector(1 downto 0);
    signal VN2006_in3 : std_logic_vector(1 downto 0);
    signal VN2006_in4 : std_logic_vector(1 downto 0);
    signal VN2006_in5 : std_logic_vector(1 downto 0);
    signal VN2007_in0 : std_logic_vector(1 downto 0);
    signal VN2007_in1 : std_logic_vector(1 downto 0);
    signal VN2007_in2 : std_logic_vector(1 downto 0);
    signal VN2007_in3 : std_logic_vector(1 downto 0);
    signal VN2007_in4 : std_logic_vector(1 downto 0);
    signal VN2007_in5 : std_logic_vector(1 downto 0);
    signal VN2008_in0 : std_logic_vector(1 downto 0);
    signal VN2008_in1 : std_logic_vector(1 downto 0);
    signal VN2008_in2 : std_logic_vector(1 downto 0);
    signal VN2008_in3 : std_logic_vector(1 downto 0);
    signal VN2008_in4 : std_logic_vector(1 downto 0);
    signal VN2008_in5 : std_logic_vector(1 downto 0);
    signal VN2009_in0 : std_logic_vector(1 downto 0);
    signal VN2009_in1 : std_logic_vector(1 downto 0);
    signal VN2009_in2 : std_logic_vector(1 downto 0);
    signal VN2009_in3 : std_logic_vector(1 downto 0);
    signal VN2009_in4 : std_logic_vector(1 downto 0);
    signal VN2009_in5 : std_logic_vector(1 downto 0);
    signal VN2010_in0 : std_logic_vector(1 downto 0);
    signal VN2010_in1 : std_logic_vector(1 downto 0);
    signal VN2010_in2 : std_logic_vector(1 downto 0);
    signal VN2010_in3 : std_logic_vector(1 downto 0);
    signal VN2010_in4 : std_logic_vector(1 downto 0);
    signal VN2010_in5 : std_logic_vector(1 downto 0);
    signal VN2011_in0 : std_logic_vector(1 downto 0);
    signal VN2011_in1 : std_logic_vector(1 downto 0);
    signal VN2011_in2 : std_logic_vector(1 downto 0);
    signal VN2011_in3 : std_logic_vector(1 downto 0);
    signal VN2011_in4 : std_logic_vector(1 downto 0);
    signal VN2011_in5 : std_logic_vector(1 downto 0);
    signal VN2012_in0 : std_logic_vector(1 downto 0);
    signal VN2012_in1 : std_logic_vector(1 downto 0);
    signal VN2012_in2 : std_logic_vector(1 downto 0);
    signal VN2012_in3 : std_logic_vector(1 downto 0);
    signal VN2012_in4 : std_logic_vector(1 downto 0);
    signal VN2012_in5 : std_logic_vector(1 downto 0);
    signal VN2013_in0 : std_logic_vector(1 downto 0);
    signal VN2013_in1 : std_logic_vector(1 downto 0);
    signal VN2013_in2 : std_logic_vector(1 downto 0);
    signal VN2013_in3 : std_logic_vector(1 downto 0);
    signal VN2013_in4 : std_logic_vector(1 downto 0);
    signal VN2013_in5 : std_logic_vector(1 downto 0);
    signal VN2014_in0 : std_logic_vector(1 downto 0);
    signal VN2014_in1 : std_logic_vector(1 downto 0);
    signal VN2014_in2 : std_logic_vector(1 downto 0);
    signal VN2014_in3 : std_logic_vector(1 downto 0);
    signal VN2014_in4 : std_logic_vector(1 downto 0);
    signal VN2014_in5 : std_logic_vector(1 downto 0);
    signal VN2015_in0 : std_logic_vector(1 downto 0);
    signal VN2015_in1 : std_logic_vector(1 downto 0);
    signal VN2015_in2 : std_logic_vector(1 downto 0);
    signal VN2015_in3 : std_logic_vector(1 downto 0);
    signal VN2015_in4 : std_logic_vector(1 downto 0);
    signal VN2015_in5 : std_logic_vector(1 downto 0);
    signal VN2016_in0 : std_logic_vector(1 downto 0);
    signal VN2016_in1 : std_logic_vector(1 downto 0);
    signal VN2016_in2 : std_logic_vector(1 downto 0);
    signal VN2016_in3 : std_logic_vector(1 downto 0);
    signal VN2016_in4 : std_logic_vector(1 downto 0);
    signal VN2016_in5 : std_logic_vector(1 downto 0);
    signal VN2017_in0 : std_logic_vector(1 downto 0);
    signal VN2017_in1 : std_logic_vector(1 downto 0);
    signal VN2017_in2 : std_logic_vector(1 downto 0);
    signal VN2017_in3 : std_logic_vector(1 downto 0);
    signal VN2017_in4 : std_logic_vector(1 downto 0);
    signal VN2017_in5 : std_logic_vector(1 downto 0);
    signal VN2018_in0 : std_logic_vector(1 downto 0);
    signal VN2018_in1 : std_logic_vector(1 downto 0);
    signal VN2018_in2 : std_logic_vector(1 downto 0);
    signal VN2018_in3 : std_logic_vector(1 downto 0);
    signal VN2018_in4 : std_logic_vector(1 downto 0);
    signal VN2018_in5 : std_logic_vector(1 downto 0);
    signal VN2019_in0 : std_logic_vector(1 downto 0);
    signal VN2019_in1 : std_logic_vector(1 downto 0);
    signal VN2019_in2 : std_logic_vector(1 downto 0);
    signal VN2019_in3 : std_logic_vector(1 downto 0);
    signal VN2019_in4 : std_logic_vector(1 downto 0);
    signal VN2019_in5 : std_logic_vector(1 downto 0);
    signal VN2020_in0 : std_logic_vector(1 downto 0);
    signal VN2020_in1 : std_logic_vector(1 downto 0);
    signal VN2020_in2 : std_logic_vector(1 downto 0);
    signal VN2020_in3 : std_logic_vector(1 downto 0);
    signal VN2020_in4 : std_logic_vector(1 downto 0);
    signal VN2020_in5 : std_logic_vector(1 downto 0);
    signal VN2021_in0 : std_logic_vector(1 downto 0);
    signal VN2021_in1 : std_logic_vector(1 downto 0);
    signal VN2021_in2 : std_logic_vector(1 downto 0);
    signal VN2021_in3 : std_logic_vector(1 downto 0);
    signal VN2021_in4 : std_logic_vector(1 downto 0);
    signal VN2021_in5 : std_logic_vector(1 downto 0);
    signal VN2022_in0 : std_logic_vector(1 downto 0);
    signal VN2022_in1 : std_logic_vector(1 downto 0);
    signal VN2022_in2 : std_logic_vector(1 downto 0);
    signal VN2022_in3 : std_logic_vector(1 downto 0);
    signal VN2022_in4 : std_logic_vector(1 downto 0);
    signal VN2022_in5 : std_logic_vector(1 downto 0);
    signal VN2023_in0 : std_logic_vector(1 downto 0);
    signal VN2023_in1 : std_logic_vector(1 downto 0);
    signal VN2023_in2 : std_logic_vector(1 downto 0);
    signal VN2023_in3 : std_logic_vector(1 downto 0);
    signal VN2023_in4 : std_logic_vector(1 downto 0);
    signal VN2023_in5 : std_logic_vector(1 downto 0);
    signal VN2024_in0 : std_logic_vector(1 downto 0);
    signal VN2024_in1 : std_logic_vector(1 downto 0);
    signal VN2024_in2 : std_logic_vector(1 downto 0);
    signal VN2024_in3 : std_logic_vector(1 downto 0);
    signal VN2024_in4 : std_logic_vector(1 downto 0);
    signal VN2024_in5 : std_logic_vector(1 downto 0);
    signal VN2025_in0 : std_logic_vector(1 downto 0);
    signal VN2025_in1 : std_logic_vector(1 downto 0);
    signal VN2025_in2 : std_logic_vector(1 downto 0);
    signal VN2025_in3 : std_logic_vector(1 downto 0);
    signal VN2025_in4 : std_logic_vector(1 downto 0);
    signal VN2025_in5 : std_logic_vector(1 downto 0);
    signal VN2026_in0 : std_logic_vector(1 downto 0);
    signal VN2026_in1 : std_logic_vector(1 downto 0);
    signal VN2026_in2 : std_logic_vector(1 downto 0);
    signal VN2026_in3 : std_logic_vector(1 downto 0);
    signal VN2026_in4 : std_logic_vector(1 downto 0);
    signal VN2026_in5 : std_logic_vector(1 downto 0);
    signal VN2027_in0 : std_logic_vector(1 downto 0);
    signal VN2027_in1 : std_logic_vector(1 downto 0);
    signal VN2027_in2 : std_logic_vector(1 downto 0);
    signal VN2027_in3 : std_logic_vector(1 downto 0);
    signal VN2027_in4 : std_logic_vector(1 downto 0);
    signal VN2027_in5 : std_logic_vector(1 downto 0);
    signal VN2028_in0 : std_logic_vector(1 downto 0);
    signal VN2028_in1 : std_logic_vector(1 downto 0);
    signal VN2028_in2 : std_logic_vector(1 downto 0);
    signal VN2028_in3 : std_logic_vector(1 downto 0);
    signal VN2028_in4 : std_logic_vector(1 downto 0);
    signal VN2028_in5 : std_logic_vector(1 downto 0);
    signal VN2029_in0 : std_logic_vector(1 downto 0);
    signal VN2029_in1 : std_logic_vector(1 downto 0);
    signal VN2029_in2 : std_logic_vector(1 downto 0);
    signal VN2029_in3 : std_logic_vector(1 downto 0);
    signal VN2029_in4 : std_logic_vector(1 downto 0);
    signal VN2029_in5 : std_logic_vector(1 downto 0);
    signal VN2030_in0 : std_logic_vector(1 downto 0);
    signal VN2030_in1 : std_logic_vector(1 downto 0);
    signal VN2030_in2 : std_logic_vector(1 downto 0);
    signal VN2030_in3 : std_logic_vector(1 downto 0);
    signal VN2030_in4 : std_logic_vector(1 downto 0);
    signal VN2030_in5 : std_logic_vector(1 downto 0);
    signal VN2031_in0 : std_logic_vector(1 downto 0);
    signal VN2031_in1 : std_logic_vector(1 downto 0);
    signal VN2031_in2 : std_logic_vector(1 downto 0);
    signal VN2031_in3 : std_logic_vector(1 downto 0);
    signal VN2031_in4 : std_logic_vector(1 downto 0);
    signal VN2031_in5 : std_logic_vector(1 downto 0);
    signal VN2032_in0 : std_logic_vector(1 downto 0);
    signal VN2032_in1 : std_logic_vector(1 downto 0);
    signal VN2032_in2 : std_logic_vector(1 downto 0);
    signal VN2032_in3 : std_logic_vector(1 downto 0);
    signal VN2032_in4 : std_logic_vector(1 downto 0);
    signal VN2032_in5 : std_logic_vector(1 downto 0);
    signal VN2033_in0 : std_logic_vector(1 downto 0);
    signal VN2033_in1 : std_logic_vector(1 downto 0);
    signal VN2033_in2 : std_logic_vector(1 downto 0);
    signal VN2033_in3 : std_logic_vector(1 downto 0);
    signal VN2033_in4 : std_logic_vector(1 downto 0);
    signal VN2033_in5 : std_logic_vector(1 downto 0);
    signal VN2034_in0 : std_logic_vector(1 downto 0);
    signal VN2034_in1 : std_logic_vector(1 downto 0);
    signal VN2034_in2 : std_logic_vector(1 downto 0);
    signal VN2034_in3 : std_logic_vector(1 downto 0);
    signal VN2034_in4 : std_logic_vector(1 downto 0);
    signal VN2034_in5 : std_logic_vector(1 downto 0);
    signal VN2035_in0 : std_logic_vector(1 downto 0);
    signal VN2035_in1 : std_logic_vector(1 downto 0);
    signal VN2035_in2 : std_logic_vector(1 downto 0);
    signal VN2035_in3 : std_logic_vector(1 downto 0);
    signal VN2035_in4 : std_logic_vector(1 downto 0);
    signal VN2035_in5 : std_logic_vector(1 downto 0);
    signal VN2036_in0 : std_logic_vector(1 downto 0);
    signal VN2036_in1 : std_logic_vector(1 downto 0);
    signal VN2036_in2 : std_logic_vector(1 downto 0);
    signal VN2036_in3 : std_logic_vector(1 downto 0);
    signal VN2036_in4 : std_logic_vector(1 downto 0);
    signal VN2036_in5 : std_logic_vector(1 downto 0);
    signal VN2037_in0 : std_logic_vector(1 downto 0);
    signal VN2037_in1 : std_logic_vector(1 downto 0);
    signal VN2037_in2 : std_logic_vector(1 downto 0);
    signal VN2037_in3 : std_logic_vector(1 downto 0);
    signal VN2037_in4 : std_logic_vector(1 downto 0);
    signal VN2037_in5 : std_logic_vector(1 downto 0);
    signal VN2038_in0 : std_logic_vector(1 downto 0);
    signal VN2038_in1 : std_logic_vector(1 downto 0);
    signal VN2038_in2 : std_logic_vector(1 downto 0);
    signal VN2038_in3 : std_logic_vector(1 downto 0);
    signal VN2038_in4 : std_logic_vector(1 downto 0);
    signal VN2038_in5 : std_logic_vector(1 downto 0);
    signal VN2039_in0 : std_logic_vector(1 downto 0);
    signal VN2039_in1 : std_logic_vector(1 downto 0);
    signal VN2039_in2 : std_logic_vector(1 downto 0);
    signal VN2039_in3 : std_logic_vector(1 downto 0);
    signal VN2039_in4 : std_logic_vector(1 downto 0);
    signal VN2039_in5 : std_logic_vector(1 downto 0);
    signal VN2040_in0 : std_logic_vector(1 downto 0);
    signal VN2040_in1 : std_logic_vector(1 downto 0);
    signal VN2040_in2 : std_logic_vector(1 downto 0);
    signal VN2040_in3 : std_logic_vector(1 downto 0);
    signal VN2040_in4 : std_logic_vector(1 downto 0);
    signal VN2040_in5 : std_logic_vector(1 downto 0);
    signal VN2041_in0 : std_logic_vector(1 downto 0);
    signal VN2041_in1 : std_logic_vector(1 downto 0);
    signal VN2041_in2 : std_logic_vector(1 downto 0);
    signal VN2041_in3 : std_logic_vector(1 downto 0);
    signal VN2041_in4 : std_logic_vector(1 downto 0);
    signal VN2041_in5 : std_logic_vector(1 downto 0);
    signal VN2042_in0 : std_logic_vector(1 downto 0);
    signal VN2042_in1 : std_logic_vector(1 downto 0);
    signal VN2042_in2 : std_logic_vector(1 downto 0);
    signal VN2042_in3 : std_logic_vector(1 downto 0);
    signal VN2042_in4 : std_logic_vector(1 downto 0);
    signal VN2042_in5 : std_logic_vector(1 downto 0);
    signal VN2043_in0 : std_logic_vector(1 downto 0);
    signal VN2043_in1 : std_logic_vector(1 downto 0);
    signal VN2043_in2 : std_logic_vector(1 downto 0);
    signal VN2043_in3 : std_logic_vector(1 downto 0);
    signal VN2043_in4 : std_logic_vector(1 downto 0);
    signal VN2043_in5 : std_logic_vector(1 downto 0);
    signal VN2044_in0 : std_logic_vector(1 downto 0);
    signal VN2044_in1 : std_logic_vector(1 downto 0);
    signal VN2044_in2 : std_logic_vector(1 downto 0);
    signal VN2044_in3 : std_logic_vector(1 downto 0);
    signal VN2044_in4 : std_logic_vector(1 downto 0);
    signal VN2044_in5 : std_logic_vector(1 downto 0);
    signal VN2045_in0 : std_logic_vector(1 downto 0);
    signal VN2045_in1 : std_logic_vector(1 downto 0);
    signal VN2045_in2 : std_logic_vector(1 downto 0);
    signal VN2045_in3 : std_logic_vector(1 downto 0);
    signal VN2045_in4 : std_logic_vector(1 downto 0);
    signal VN2045_in5 : std_logic_vector(1 downto 0);
    signal VN2046_in0 : std_logic_vector(1 downto 0);
    signal VN2046_in1 : std_logic_vector(1 downto 0);
    signal VN2046_in2 : std_logic_vector(1 downto 0);
    signal VN2046_in3 : std_logic_vector(1 downto 0);
    signal VN2046_in4 : std_logic_vector(1 downto 0);
    signal VN2046_in5 : std_logic_vector(1 downto 0);
    signal VN2047_in0 : std_logic_vector(1 downto 0);
    signal VN2047_in1 : std_logic_vector(1 downto 0);
    signal VN2047_in2 : std_logic_vector(1 downto 0);
    signal VN2047_in3 : std_logic_vector(1 downto 0);
    signal VN2047_in4 : std_logic_vector(1 downto 0);
    signal VN2047_in5 : std_logic_vector(1 downto 0);
    

begin

  VN0_in0 <= VN_sign_in(0) & VN_data_in(0);
  VN0_in1 <= VN_sign_in(1) & VN_data_in(1);
  VN0_in2 <= VN_sign_in(2) & VN_data_in(2);
  VN0_in3 <= VN_sign_in(3) & VN_data_in(3);
  VN0_in4 <= VN_sign_in(4) & VN_data_in(4);
  VN0_in5 <= VN_sign_in(5) & VN_data_in(5);
  VN1_in0 <= VN_sign_in(6) & VN_data_in(6);
  VN1_in1 <= VN_sign_in(7) & VN_data_in(7);
  VN1_in2 <= VN_sign_in(8) & VN_data_in(8);
  VN1_in3 <= VN_sign_in(9) & VN_data_in(9);
  VN1_in4 <= VN_sign_in(10) & VN_data_in(10);
  VN1_in5 <= VN_sign_in(11) & VN_data_in(11);
  VN2_in0 <= VN_sign_in(12) & VN_data_in(12);
  VN2_in1 <= VN_sign_in(13) & VN_data_in(13);
  VN2_in2 <= VN_sign_in(14) & VN_data_in(14);
  VN2_in3 <= VN_sign_in(15) & VN_data_in(15);
  VN2_in4 <= VN_sign_in(16) & VN_data_in(16);
  VN2_in5 <= VN_sign_in(17) & VN_data_in(17);
  VN3_in0 <= VN_sign_in(18) & VN_data_in(18);
  VN3_in1 <= VN_sign_in(19) & VN_data_in(19);
  VN3_in2 <= VN_sign_in(20) & VN_data_in(20);
  VN3_in3 <= VN_sign_in(21) & VN_data_in(21);
  VN3_in4 <= VN_sign_in(22) & VN_data_in(22);
  VN3_in5 <= VN_sign_in(23) & VN_data_in(23);
  VN4_in0 <= VN_sign_in(24) & VN_data_in(24);
  VN4_in1 <= VN_sign_in(25) & VN_data_in(25);
  VN4_in2 <= VN_sign_in(26) & VN_data_in(26);
  VN4_in3 <= VN_sign_in(27) & VN_data_in(27);
  VN4_in4 <= VN_sign_in(28) & VN_data_in(28);
  VN4_in5 <= VN_sign_in(29) & VN_data_in(29);
  VN5_in0 <= VN_sign_in(30) & VN_data_in(30);
  VN5_in1 <= VN_sign_in(31) & VN_data_in(31);
  VN5_in2 <= VN_sign_in(32) & VN_data_in(32);
  VN5_in3 <= VN_sign_in(33) & VN_data_in(33);
  VN5_in4 <= VN_sign_in(34) & VN_data_in(34);
  VN5_in5 <= VN_sign_in(35) & VN_data_in(35);
  VN6_in0 <= VN_sign_in(36) & VN_data_in(36);
  VN6_in1 <= VN_sign_in(37) & VN_data_in(37);
  VN6_in2 <= VN_sign_in(38) & VN_data_in(38);
  VN6_in3 <= VN_sign_in(39) & VN_data_in(39);
  VN6_in4 <= VN_sign_in(40) & VN_data_in(40);
  VN6_in5 <= VN_sign_in(41) & VN_data_in(41);
  VN7_in0 <= VN_sign_in(42) & VN_data_in(42);
  VN7_in1 <= VN_sign_in(43) & VN_data_in(43);
  VN7_in2 <= VN_sign_in(44) & VN_data_in(44);
  VN7_in3 <= VN_sign_in(45) & VN_data_in(45);
  VN7_in4 <= VN_sign_in(46) & VN_data_in(46);
  VN7_in5 <= VN_sign_in(47) & VN_data_in(47);
  VN8_in0 <= VN_sign_in(48) & VN_data_in(48);
  VN8_in1 <= VN_sign_in(49) & VN_data_in(49);
  VN8_in2 <= VN_sign_in(50) & VN_data_in(50);
  VN8_in3 <= VN_sign_in(51) & VN_data_in(51);
  VN8_in4 <= VN_sign_in(52) & VN_data_in(52);
  VN8_in5 <= VN_sign_in(53) & VN_data_in(53);
  VN9_in0 <= VN_sign_in(54) & VN_data_in(54);
  VN9_in1 <= VN_sign_in(55) & VN_data_in(55);
  VN9_in2 <= VN_sign_in(56) & VN_data_in(56);
  VN9_in3 <= VN_sign_in(57) & VN_data_in(57);
  VN9_in4 <= VN_sign_in(58) & VN_data_in(58);
  VN9_in5 <= VN_sign_in(59) & VN_data_in(59);
  VN10_in0 <= VN_sign_in(60) & VN_data_in(60);
  VN10_in1 <= VN_sign_in(61) & VN_data_in(61);
  VN10_in2 <= VN_sign_in(62) & VN_data_in(62);
  VN10_in3 <= VN_sign_in(63) & VN_data_in(63);
  VN10_in4 <= VN_sign_in(64) & VN_data_in(64);
  VN10_in5 <= VN_sign_in(65) & VN_data_in(65);
  VN11_in0 <= VN_sign_in(66) & VN_data_in(66);
  VN11_in1 <= VN_sign_in(67) & VN_data_in(67);
  VN11_in2 <= VN_sign_in(68) & VN_data_in(68);
  VN11_in3 <= VN_sign_in(69) & VN_data_in(69);
  VN11_in4 <= VN_sign_in(70) & VN_data_in(70);
  VN11_in5 <= VN_sign_in(71) & VN_data_in(71);
  VN12_in0 <= VN_sign_in(72) & VN_data_in(72);
  VN12_in1 <= VN_sign_in(73) & VN_data_in(73);
  VN12_in2 <= VN_sign_in(74) & VN_data_in(74);
  VN12_in3 <= VN_sign_in(75) & VN_data_in(75);
  VN12_in4 <= VN_sign_in(76) & VN_data_in(76);
  VN12_in5 <= VN_sign_in(77) & VN_data_in(77);
  VN13_in0 <= VN_sign_in(78) & VN_data_in(78);
  VN13_in1 <= VN_sign_in(79) & VN_data_in(79);
  VN13_in2 <= VN_sign_in(80) & VN_data_in(80);
  VN13_in3 <= VN_sign_in(81) & VN_data_in(81);
  VN13_in4 <= VN_sign_in(82) & VN_data_in(82);
  VN13_in5 <= VN_sign_in(83) & VN_data_in(83);
  VN14_in0 <= VN_sign_in(84) & VN_data_in(84);
  VN14_in1 <= VN_sign_in(85) & VN_data_in(85);
  VN14_in2 <= VN_sign_in(86) & VN_data_in(86);
  VN14_in3 <= VN_sign_in(87) & VN_data_in(87);
  VN14_in4 <= VN_sign_in(88) & VN_data_in(88);
  VN14_in5 <= VN_sign_in(89) & VN_data_in(89);
  VN15_in0 <= VN_sign_in(90) & VN_data_in(90);
  VN15_in1 <= VN_sign_in(91) & VN_data_in(91);
  VN15_in2 <= VN_sign_in(92) & VN_data_in(92);
  VN15_in3 <= VN_sign_in(93) & VN_data_in(93);
  VN15_in4 <= VN_sign_in(94) & VN_data_in(94);
  VN15_in5 <= VN_sign_in(95) & VN_data_in(95);
  VN16_in0 <= VN_sign_in(96) & VN_data_in(96);
  VN16_in1 <= VN_sign_in(97) & VN_data_in(97);
  VN16_in2 <= VN_sign_in(98) & VN_data_in(98);
  VN16_in3 <= VN_sign_in(99) & VN_data_in(99);
  VN16_in4 <= VN_sign_in(100) & VN_data_in(100);
  VN16_in5 <= VN_sign_in(101) & VN_data_in(101);
  VN17_in0 <= VN_sign_in(102) & VN_data_in(102);
  VN17_in1 <= VN_sign_in(103) & VN_data_in(103);
  VN17_in2 <= VN_sign_in(104) & VN_data_in(104);
  VN17_in3 <= VN_sign_in(105) & VN_data_in(105);
  VN17_in4 <= VN_sign_in(106) & VN_data_in(106);
  VN17_in5 <= VN_sign_in(107) & VN_data_in(107);
  VN18_in0 <= VN_sign_in(108) & VN_data_in(108);
  VN18_in1 <= VN_sign_in(109) & VN_data_in(109);
  VN18_in2 <= VN_sign_in(110) & VN_data_in(110);
  VN18_in3 <= VN_sign_in(111) & VN_data_in(111);
  VN18_in4 <= VN_sign_in(112) & VN_data_in(112);
  VN18_in5 <= VN_sign_in(113) & VN_data_in(113);
  VN19_in0 <= VN_sign_in(114) & VN_data_in(114);
  VN19_in1 <= VN_sign_in(115) & VN_data_in(115);
  VN19_in2 <= VN_sign_in(116) & VN_data_in(116);
  VN19_in3 <= VN_sign_in(117) & VN_data_in(117);
  VN19_in4 <= VN_sign_in(118) & VN_data_in(118);
  VN19_in5 <= VN_sign_in(119) & VN_data_in(119);
  VN20_in0 <= VN_sign_in(120) & VN_data_in(120);
  VN20_in1 <= VN_sign_in(121) & VN_data_in(121);
  VN20_in2 <= VN_sign_in(122) & VN_data_in(122);
  VN20_in3 <= VN_sign_in(123) & VN_data_in(123);
  VN20_in4 <= VN_sign_in(124) & VN_data_in(124);
  VN20_in5 <= VN_sign_in(125) & VN_data_in(125);
  VN21_in0 <= VN_sign_in(126) & VN_data_in(126);
  VN21_in1 <= VN_sign_in(127) & VN_data_in(127);
  VN21_in2 <= VN_sign_in(128) & VN_data_in(128);
  VN21_in3 <= VN_sign_in(129) & VN_data_in(129);
  VN21_in4 <= VN_sign_in(130) & VN_data_in(130);
  VN21_in5 <= VN_sign_in(131) & VN_data_in(131);
  VN22_in0 <= VN_sign_in(132) & VN_data_in(132);
  VN22_in1 <= VN_sign_in(133) & VN_data_in(133);
  VN22_in2 <= VN_sign_in(134) & VN_data_in(134);
  VN22_in3 <= VN_sign_in(135) & VN_data_in(135);
  VN22_in4 <= VN_sign_in(136) & VN_data_in(136);
  VN22_in5 <= VN_sign_in(137) & VN_data_in(137);
  VN23_in0 <= VN_sign_in(138) & VN_data_in(138);
  VN23_in1 <= VN_sign_in(139) & VN_data_in(139);
  VN23_in2 <= VN_sign_in(140) & VN_data_in(140);
  VN23_in3 <= VN_sign_in(141) & VN_data_in(141);
  VN23_in4 <= VN_sign_in(142) & VN_data_in(142);
  VN23_in5 <= VN_sign_in(143) & VN_data_in(143);
  VN24_in0 <= VN_sign_in(144) & VN_data_in(144);
  VN24_in1 <= VN_sign_in(145) & VN_data_in(145);
  VN24_in2 <= VN_sign_in(146) & VN_data_in(146);
  VN24_in3 <= VN_sign_in(147) & VN_data_in(147);
  VN24_in4 <= VN_sign_in(148) & VN_data_in(148);
  VN24_in5 <= VN_sign_in(149) & VN_data_in(149);
  VN25_in0 <= VN_sign_in(150) & VN_data_in(150);
  VN25_in1 <= VN_sign_in(151) & VN_data_in(151);
  VN25_in2 <= VN_sign_in(152) & VN_data_in(152);
  VN25_in3 <= VN_sign_in(153) & VN_data_in(153);
  VN25_in4 <= VN_sign_in(154) & VN_data_in(154);
  VN25_in5 <= VN_sign_in(155) & VN_data_in(155);
  VN26_in0 <= VN_sign_in(156) & VN_data_in(156);
  VN26_in1 <= VN_sign_in(157) & VN_data_in(157);
  VN26_in2 <= VN_sign_in(158) & VN_data_in(158);
  VN26_in3 <= VN_sign_in(159) & VN_data_in(159);
  VN26_in4 <= VN_sign_in(160) & VN_data_in(160);
  VN26_in5 <= VN_sign_in(161) & VN_data_in(161);
  VN27_in0 <= VN_sign_in(162) & VN_data_in(162);
  VN27_in1 <= VN_sign_in(163) & VN_data_in(163);
  VN27_in2 <= VN_sign_in(164) & VN_data_in(164);
  VN27_in3 <= VN_sign_in(165) & VN_data_in(165);
  VN27_in4 <= VN_sign_in(166) & VN_data_in(166);
  VN27_in5 <= VN_sign_in(167) & VN_data_in(167);
  VN28_in0 <= VN_sign_in(168) & VN_data_in(168);
  VN28_in1 <= VN_sign_in(169) & VN_data_in(169);
  VN28_in2 <= VN_sign_in(170) & VN_data_in(170);
  VN28_in3 <= VN_sign_in(171) & VN_data_in(171);
  VN28_in4 <= VN_sign_in(172) & VN_data_in(172);
  VN28_in5 <= VN_sign_in(173) & VN_data_in(173);
  VN29_in0 <= VN_sign_in(174) & VN_data_in(174);
  VN29_in1 <= VN_sign_in(175) & VN_data_in(175);
  VN29_in2 <= VN_sign_in(176) & VN_data_in(176);
  VN29_in3 <= VN_sign_in(177) & VN_data_in(177);
  VN29_in4 <= VN_sign_in(178) & VN_data_in(178);
  VN29_in5 <= VN_sign_in(179) & VN_data_in(179);
  VN30_in0 <= VN_sign_in(180) & VN_data_in(180);
  VN30_in1 <= VN_sign_in(181) & VN_data_in(181);
  VN30_in2 <= VN_sign_in(182) & VN_data_in(182);
  VN30_in3 <= VN_sign_in(183) & VN_data_in(183);
  VN30_in4 <= VN_sign_in(184) & VN_data_in(184);
  VN30_in5 <= VN_sign_in(185) & VN_data_in(185);
  VN31_in0 <= VN_sign_in(186) & VN_data_in(186);
  VN31_in1 <= VN_sign_in(187) & VN_data_in(187);
  VN31_in2 <= VN_sign_in(188) & VN_data_in(188);
  VN31_in3 <= VN_sign_in(189) & VN_data_in(189);
  VN31_in4 <= VN_sign_in(190) & VN_data_in(190);
  VN31_in5 <= VN_sign_in(191) & VN_data_in(191);
  VN32_in0 <= VN_sign_in(192) & VN_data_in(192);
  VN32_in1 <= VN_sign_in(193) & VN_data_in(193);
  VN32_in2 <= VN_sign_in(194) & VN_data_in(194);
  VN32_in3 <= VN_sign_in(195) & VN_data_in(195);
  VN32_in4 <= VN_sign_in(196) & VN_data_in(196);
  VN32_in5 <= VN_sign_in(197) & VN_data_in(197);
  VN33_in0 <= VN_sign_in(198) & VN_data_in(198);
  VN33_in1 <= VN_sign_in(199) & VN_data_in(199);
  VN33_in2 <= VN_sign_in(200) & VN_data_in(200);
  VN33_in3 <= VN_sign_in(201) & VN_data_in(201);
  VN33_in4 <= VN_sign_in(202) & VN_data_in(202);
  VN33_in5 <= VN_sign_in(203) & VN_data_in(203);
  VN34_in0 <= VN_sign_in(204) & VN_data_in(204);
  VN34_in1 <= VN_sign_in(205) & VN_data_in(205);
  VN34_in2 <= VN_sign_in(206) & VN_data_in(206);
  VN34_in3 <= VN_sign_in(207) & VN_data_in(207);
  VN34_in4 <= VN_sign_in(208) & VN_data_in(208);
  VN34_in5 <= VN_sign_in(209) & VN_data_in(209);
  VN35_in0 <= VN_sign_in(210) & VN_data_in(210);
  VN35_in1 <= VN_sign_in(211) & VN_data_in(211);
  VN35_in2 <= VN_sign_in(212) & VN_data_in(212);
  VN35_in3 <= VN_sign_in(213) & VN_data_in(213);
  VN35_in4 <= VN_sign_in(214) & VN_data_in(214);
  VN35_in5 <= VN_sign_in(215) & VN_data_in(215);
  VN36_in0 <= VN_sign_in(216) & VN_data_in(216);
  VN36_in1 <= VN_sign_in(217) & VN_data_in(217);
  VN36_in2 <= VN_sign_in(218) & VN_data_in(218);
  VN36_in3 <= VN_sign_in(219) & VN_data_in(219);
  VN36_in4 <= VN_sign_in(220) & VN_data_in(220);
  VN36_in5 <= VN_sign_in(221) & VN_data_in(221);
  VN37_in0 <= VN_sign_in(222) & VN_data_in(222);
  VN37_in1 <= VN_sign_in(223) & VN_data_in(223);
  VN37_in2 <= VN_sign_in(224) & VN_data_in(224);
  VN37_in3 <= VN_sign_in(225) & VN_data_in(225);
  VN37_in4 <= VN_sign_in(226) & VN_data_in(226);
  VN37_in5 <= VN_sign_in(227) & VN_data_in(227);
  VN38_in0 <= VN_sign_in(228) & VN_data_in(228);
  VN38_in1 <= VN_sign_in(229) & VN_data_in(229);
  VN38_in2 <= VN_sign_in(230) & VN_data_in(230);
  VN38_in3 <= VN_sign_in(231) & VN_data_in(231);
  VN38_in4 <= VN_sign_in(232) & VN_data_in(232);
  VN38_in5 <= VN_sign_in(233) & VN_data_in(233);
  VN39_in0 <= VN_sign_in(234) & VN_data_in(234);
  VN39_in1 <= VN_sign_in(235) & VN_data_in(235);
  VN39_in2 <= VN_sign_in(236) & VN_data_in(236);
  VN39_in3 <= VN_sign_in(237) & VN_data_in(237);
  VN39_in4 <= VN_sign_in(238) & VN_data_in(238);
  VN39_in5 <= VN_sign_in(239) & VN_data_in(239);
  VN40_in0 <= VN_sign_in(240) & VN_data_in(240);
  VN40_in1 <= VN_sign_in(241) & VN_data_in(241);
  VN40_in2 <= VN_sign_in(242) & VN_data_in(242);
  VN40_in3 <= VN_sign_in(243) & VN_data_in(243);
  VN40_in4 <= VN_sign_in(244) & VN_data_in(244);
  VN40_in5 <= VN_sign_in(245) & VN_data_in(245);
  VN41_in0 <= VN_sign_in(246) & VN_data_in(246);
  VN41_in1 <= VN_sign_in(247) & VN_data_in(247);
  VN41_in2 <= VN_sign_in(248) & VN_data_in(248);
  VN41_in3 <= VN_sign_in(249) & VN_data_in(249);
  VN41_in4 <= VN_sign_in(250) & VN_data_in(250);
  VN41_in5 <= VN_sign_in(251) & VN_data_in(251);
  VN42_in0 <= VN_sign_in(252) & VN_data_in(252);
  VN42_in1 <= VN_sign_in(253) & VN_data_in(253);
  VN42_in2 <= VN_sign_in(254) & VN_data_in(254);
  VN42_in3 <= VN_sign_in(255) & VN_data_in(255);
  VN42_in4 <= VN_sign_in(256) & VN_data_in(256);
  VN42_in5 <= VN_sign_in(257) & VN_data_in(257);
  VN43_in0 <= VN_sign_in(258) & VN_data_in(258);
  VN43_in1 <= VN_sign_in(259) & VN_data_in(259);
  VN43_in2 <= VN_sign_in(260) & VN_data_in(260);
  VN43_in3 <= VN_sign_in(261) & VN_data_in(261);
  VN43_in4 <= VN_sign_in(262) & VN_data_in(262);
  VN43_in5 <= VN_sign_in(263) & VN_data_in(263);
  VN44_in0 <= VN_sign_in(264) & VN_data_in(264);
  VN44_in1 <= VN_sign_in(265) & VN_data_in(265);
  VN44_in2 <= VN_sign_in(266) & VN_data_in(266);
  VN44_in3 <= VN_sign_in(267) & VN_data_in(267);
  VN44_in4 <= VN_sign_in(268) & VN_data_in(268);
  VN44_in5 <= VN_sign_in(269) & VN_data_in(269);
  VN45_in0 <= VN_sign_in(270) & VN_data_in(270);
  VN45_in1 <= VN_sign_in(271) & VN_data_in(271);
  VN45_in2 <= VN_sign_in(272) & VN_data_in(272);
  VN45_in3 <= VN_sign_in(273) & VN_data_in(273);
  VN45_in4 <= VN_sign_in(274) & VN_data_in(274);
  VN45_in5 <= VN_sign_in(275) & VN_data_in(275);
  VN46_in0 <= VN_sign_in(276) & VN_data_in(276);
  VN46_in1 <= VN_sign_in(277) & VN_data_in(277);
  VN46_in2 <= VN_sign_in(278) & VN_data_in(278);
  VN46_in3 <= VN_sign_in(279) & VN_data_in(279);
  VN46_in4 <= VN_sign_in(280) & VN_data_in(280);
  VN46_in5 <= VN_sign_in(281) & VN_data_in(281);
  VN47_in0 <= VN_sign_in(282) & VN_data_in(282);
  VN47_in1 <= VN_sign_in(283) & VN_data_in(283);
  VN47_in2 <= VN_sign_in(284) & VN_data_in(284);
  VN47_in3 <= VN_sign_in(285) & VN_data_in(285);
  VN47_in4 <= VN_sign_in(286) & VN_data_in(286);
  VN47_in5 <= VN_sign_in(287) & VN_data_in(287);
  VN48_in0 <= VN_sign_in(288) & VN_data_in(288);
  VN48_in1 <= VN_sign_in(289) & VN_data_in(289);
  VN48_in2 <= VN_sign_in(290) & VN_data_in(290);
  VN48_in3 <= VN_sign_in(291) & VN_data_in(291);
  VN48_in4 <= VN_sign_in(292) & VN_data_in(292);
  VN48_in5 <= VN_sign_in(293) & VN_data_in(293);
  VN49_in0 <= VN_sign_in(294) & VN_data_in(294);
  VN49_in1 <= VN_sign_in(295) & VN_data_in(295);
  VN49_in2 <= VN_sign_in(296) & VN_data_in(296);
  VN49_in3 <= VN_sign_in(297) & VN_data_in(297);
  VN49_in4 <= VN_sign_in(298) & VN_data_in(298);
  VN49_in5 <= VN_sign_in(299) & VN_data_in(299);
  VN50_in0 <= VN_sign_in(300) & VN_data_in(300);
  VN50_in1 <= VN_sign_in(301) & VN_data_in(301);
  VN50_in2 <= VN_sign_in(302) & VN_data_in(302);
  VN50_in3 <= VN_sign_in(303) & VN_data_in(303);
  VN50_in4 <= VN_sign_in(304) & VN_data_in(304);
  VN50_in5 <= VN_sign_in(305) & VN_data_in(305);
  VN51_in0 <= VN_sign_in(306) & VN_data_in(306);
  VN51_in1 <= VN_sign_in(307) & VN_data_in(307);
  VN51_in2 <= VN_sign_in(308) & VN_data_in(308);
  VN51_in3 <= VN_sign_in(309) & VN_data_in(309);
  VN51_in4 <= VN_sign_in(310) & VN_data_in(310);
  VN51_in5 <= VN_sign_in(311) & VN_data_in(311);
  VN52_in0 <= VN_sign_in(312) & VN_data_in(312);
  VN52_in1 <= VN_sign_in(313) & VN_data_in(313);
  VN52_in2 <= VN_sign_in(314) & VN_data_in(314);
  VN52_in3 <= VN_sign_in(315) & VN_data_in(315);
  VN52_in4 <= VN_sign_in(316) & VN_data_in(316);
  VN52_in5 <= VN_sign_in(317) & VN_data_in(317);
  VN53_in0 <= VN_sign_in(318) & VN_data_in(318);
  VN53_in1 <= VN_sign_in(319) & VN_data_in(319);
  VN53_in2 <= VN_sign_in(320) & VN_data_in(320);
  VN53_in3 <= VN_sign_in(321) & VN_data_in(321);
  VN53_in4 <= VN_sign_in(322) & VN_data_in(322);
  VN53_in5 <= VN_sign_in(323) & VN_data_in(323);
  VN54_in0 <= VN_sign_in(324) & VN_data_in(324);
  VN54_in1 <= VN_sign_in(325) & VN_data_in(325);
  VN54_in2 <= VN_sign_in(326) & VN_data_in(326);
  VN54_in3 <= VN_sign_in(327) & VN_data_in(327);
  VN54_in4 <= VN_sign_in(328) & VN_data_in(328);
  VN54_in5 <= VN_sign_in(329) & VN_data_in(329);
  VN55_in0 <= VN_sign_in(330) & VN_data_in(330);
  VN55_in1 <= VN_sign_in(331) & VN_data_in(331);
  VN55_in2 <= VN_sign_in(332) & VN_data_in(332);
  VN55_in3 <= VN_sign_in(333) & VN_data_in(333);
  VN55_in4 <= VN_sign_in(334) & VN_data_in(334);
  VN55_in5 <= VN_sign_in(335) & VN_data_in(335);
  VN56_in0 <= VN_sign_in(336) & VN_data_in(336);
  VN56_in1 <= VN_sign_in(337) & VN_data_in(337);
  VN56_in2 <= VN_sign_in(338) & VN_data_in(338);
  VN56_in3 <= VN_sign_in(339) & VN_data_in(339);
  VN56_in4 <= VN_sign_in(340) & VN_data_in(340);
  VN56_in5 <= VN_sign_in(341) & VN_data_in(341);
  VN57_in0 <= VN_sign_in(342) & VN_data_in(342);
  VN57_in1 <= VN_sign_in(343) & VN_data_in(343);
  VN57_in2 <= VN_sign_in(344) & VN_data_in(344);
  VN57_in3 <= VN_sign_in(345) & VN_data_in(345);
  VN57_in4 <= VN_sign_in(346) & VN_data_in(346);
  VN57_in5 <= VN_sign_in(347) & VN_data_in(347);
  VN58_in0 <= VN_sign_in(348) & VN_data_in(348);
  VN58_in1 <= VN_sign_in(349) & VN_data_in(349);
  VN58_in2 <= VN_sign_in(350) & VN_data_in(350);
  VN58_in3 <= VN_sign_in(351) & VN_data_in(351);
  VN58_in4 <= VN_sign_in(352) & VN_data_in(352);
  VN58_in5 <= VN_sign_in(353) & VN_data_in(353);
  VN59_in0 <= VN_sign_in(354) & VN_data_in(354);
  VN59_in1 <= VN_sign_in(355) & VN_data_in(355);
  VN59_in2 <= VN_sign_in(356) & VN_data_in(356);
  VN59_in3 <= VN_sign_in(357) & VN_data_in(357);
  VN59_in4 <= VN_sign_in(358) & VN_data_in(358);
  VN59_in5 <= VN_sign_in(359) & VN_data_in(359);
  VN60_in0 <= VN_sign_in(360) & VN_data_in(360);
  VN60_in1 <= VN_sign_in(361) & VN_data_in(361);
  VN60_in2 <= VN_sign_in(362) & VN_data_in(362);
  VN60_in3 <= VN_sign_in(363) & VN_data_in(363);
  VN60_in4 <= VN_sign_in(364) & VN_data_in(364);
  VN60_in5 <= VN_sign_in(365) & VN_data_in(365);
  VN61_in0 <= VN_sign_in(366) & VN_data_in(366);
  VN61_in1 <= VN_sign_in(367) & VN_data_in(367);
  VN61_in2 <= VN_sign_in(368) & VN_data_in(368);
  VN61_in3 <= VN_sign_in(369) & VN_data_in(369);
  VN61_in4 <= VN_sign_in(370) & VN_data_in(370);
  VN61_in5 <= VN_sign_in(371) & VN_data_in(371);
  VN62_in0 <= VN_sign_in(372) & VN_data_in(372);
  VN62_in1 <= VN_sign_in(373) & VN_data_in(373);
  VN62_in2 <= VN_sign_in(374) & VN_data_in(374);
  VN62_in3 <= VN_sign_in(375) & VN_data_in(375);
  VN62_in4 <= VN_sign_in(376) & VN_data_in(376);
  VN62_in5 <= VN_sign_in(377) & VN_data_in(377);
  VN63_in0 <= VN_sign_in(378) & VN_data_in(378);
  VN63_in1 <= VN_sign_in(379) & VN_data_in(379);
  VN63_in2 <= VN_sign_in(380) & VN_data_in(380);
  VN63_in3 <= VN_sign_in(381) & VN_data_in(381);
  VN63_in4 <= VN_sign_in(382) & VN_data_in(382);
  VN63_in5 <= VN_sign_in(383) & VN_data_in(383);
  VN64_in0 <= VN_sign_in(384) & VN_data_in(384);
  VN64_in1 <= VN_sign_in(385) & VN_data_in(385);
  VN64_in2 <= VN_sign_in(386) & VN_data_in(386);
  VN64_in3 <= VN_sign_in(387) & VN_data_in(387);
  VN64_in4 <= VN_sign_in(388) & VN_data_in(388);
  VN64_in5 <= VN_sign_in(389) & VN_data_in(389);
  VN65_in0 <= VN_sign_in(390) & VN_data_in(390);
  VN65_in1 <= VN_sign_in(391) & VN_data_in(391);
  VN65_in2 <= VN_sign_in(392) & VN_data_in(392);
  VN65_in3 <= VN_sign_in(393) & VN_data_in(393);
  VN65_in4 <= VN_sign_in(394) & VN_data_in(394);
  VN65_in5 <= VN_sign_in(395) & VN_data_in(395);
  VN66_in0 <= VN_sign_in(396) & VN_data_in(396);
  VN66_in1 <= VN_sign_in(397) & VN_data_in(397);
  VN66_in2 <= VN_sign_in(398) & VN_data_in(398);
  VN66_in3 <= VN_sign_in(399) & VN_data_in(399);
  VN66_in4 <= VN_sign_in(400) & VN_data_in(400);
  VN66_in5 <= VN_sign_in(401) & VN_data_in(401);
  VN67_in0 <= VN_sign_in(402) & VN_data_in(402);
  VN67_in1 <= VN_sign_in(403) & VN_data_in(403);
  VN67_in2 <= VN_sign_in(404) & VN_data_in(404);
  VN67_in3 <= VN_sign_in(405) & VN_data_in(405);
  VN67_in4 <= VN_sign_in(406) & VN_data_in(406);
  VN67_in5 <= VN_sign_in(407) & VN_data_in(407);
  VN68_in0 <= VN_sign_in(408) & VN_data_in(408);
  VN68_in1 <= VN_sign_in(409) & VN_data_in(409);
  VN68_in2 <= VN_sign_in(410) & VN_data_in(410);
  VN68_in3 <= VN_sign_in(411) & VN_data_in(411);
  VN68_in4 <= VN_sign_in(412) & VN_data_in(412);
  VN68_in5 <= VN_sign_in(413) & VN_data_in(413);
  VN69_in0 <= VN_sign_in(414) & VN_data_in(414);
  VN69_in1 <= VN_sign_in(415) & VN_data_in(415);
  VN69_in2 <= VN_sign_in(416) & VN_data_in(416);
  VN69_in3 <= VN_sign_in(417) & VN_data_in(417);
  VN69_in4 <= VN_sign_in(418) & VN_data_in(418);
  VN69_in5 <= VN_sign_in(419) & VN_data_in(419);
  VN70_in0 <= VN_sign_in(420) & VN_data_in(420);
  VN70_in1 <= VN_sign_in(421) & VN_data_in(421);
  VN70_in2 <= VN_sign_in(422) & VN_data_in(422);
  VN70_in3 <= VN_sign_in(423) & VN_data_in(423);
  VN70_in4 <= VN_sign_in(424) & VN_data_in(424);
  VN70_in5 <= VN_sign_in(425) & VN_data_in(425);
  VN71_in0 <= VN_sign_in(426) & VN_data_in(426);
  VN71_in1 <= VN_sign_in(427) & VN_data_in(427);
  VN71_in2 <= VN_sign_in(428) & VN_data_in(428);
  VN71_in3 <= VN_sign_in(429) & VN_data_in(429);
  VN71_in4 <= VN_sign_in(430) & VN_data_in(430);
  VN71_in5 <= VN_sign_in(431) & VN_data_in(431);
  VN72_in0 <= VN_sign_in(432) & VN_data_in(432);
  VN72_in1 <= VN_sign_in(433) & VN_data_in(433);
  VN72_in2 <= VN_sign_in(434) & VN_data_in(434);
  VN72_in3 <= VN_sign_in(435) & VN_data_in(435);
  VN72_in4 <= VN_sign_in(436) & VN_data_in(436);
  VN72_in5 <= VN_sign_in(437) & VN_data_in(437);
  VN73_in0 <= VN_sign_in(438) & VN_data_in(438);
  VN73_in1 <= VN_sign_in(439) & VN_data_in(439);
  VN73_in2 <= VN_sign_in(440) & VN_data_in(440);
  VN73_in3 <= VN_sign_in(441) & VN_data_in(441);
  VN73_in4 <= VN_sign_in(442) & VN_data_in(442);
  VN73_in5 <= VN_sign_in(443) & VN_data_in(443);
  VN74_in0 <= VN_sign_in(444) & VN_data_in(444);
  VN74_in1 <= VN_sign_in(445) & VN_data_in(445);
  VN74_in2 <= VN_sign_in(446) & VN_data_in(446);
  VN74_in3 <= VN_sign_in(447) & VN_data_in(447);
  VN74_in4 <= VN_sign_in(448) & VN_data_in(448);
  VN74_in5 <= VN_sign_in(449) & VN_data_in(449);
  VN75_in0 <= VN_sign_in(450) & VN_data_in(450);
  VN75_in1 <= VN_sign_in(451) & VN_data_in(451);
  VN75_in2 <= VN_sign_in(452) & VN_data_in(452);
  VN75_in3 <= VN_sign_in(453) & VN_data_in(453);
  VN75_in4 <= VN_sign_in(454) & VN_data_in(454);
  VN75_in5 <= VN_sign_in(455) & VN_data_in(455);
  VN76_in0 <= VN_sign_in(456) & VN_data_in(456);
  VN76_in1 <= VN_sign_in(457) & VN_data_in(457);
  VN76_in2 <= VN_sign_in(458) & VN_data_in(458);
  VN76_in3 <= VN_sign_in(459) & VN_data_in(459);
  VN76_in4 <= VN_sign_in(460) & VN_data_in(460);
  VN76_in5 <= VN_sign_in(461) & VN_data_in(461);
  VN77_in0 <= VN_sign_in(462) & VN_data_in(462);
  VN77_in1 <= VN_sign_in(463) & VN_data_in(463);
  VN77_in2 <= VN_sign_in(464) & VN_data_in(464);
  VN77_in3 <= VN_sign_in(465) & VN_data_in(465);
  VN77_in4 <= VN_sign_in(466) & VN_data_in(466);
  VN77_in5 <= VN_sign_in(467) & VN_data_in(467);
  VN78_in0 <= VN_sign_in(468) & VN_data_in(468);
  VN78_in1 <= VN_sign_in(469) & VN_data_in(469);
  VN78_in2 <= VN_sign_in(470) & VN_data_in(470);
  VN78_in3 <= VN_sign_in(471) & VN_data_in(471);
  VN78_in4 <= VN_sign_in(472) & VN_data_in(472);
  VN78_in5 <= VN_sign_in(473) & VN_data_in(473);
  VN79_in0 <= VN_sign_in(474) & VN_data_in(474);
  VN79_in1 <= VN_sign_in(475) & VN_data_in(475);
  VN79_in2 <= VN_sign_in(476) & VN_data_in(476);
  VN79_in3 <= VN_sign_in(477) & VN_data_in(477);
  VN79_in4 <= VN_sign_in(478) & VN_data_in(478);
  VN79_in5 <= VN_sign_in(479) & VN_data_in(479);
  VN80_in0 <= VN_sign_in(480) & VN_data_in(480);
  VN80_in1 <= VN_sign_in(481) & VN_data_in(481);
  VN80_in2 <= VN_sign_in(482) & VN_data_in(482);
  VN80_in3 <= VN_sign_in(483) & VN_data_in(483);
  VN80_in4 <= VN_sign_in(484) & VN_data_in(484);
  VN80_in5 <= VN_sign_in(485) & VN_data_in(485);
  VN81_in0 <= VN_sign_in(486) & VN_data_in(486);
  VN81_in1 <= VN_sign_in(487) & VN_data_in(487);
  VN81_in2 <= VN_sign_in(488) & VN_data_in(488);
  VN81_in3 <= VN_sign_in(489) & VN_data_in(489);
  VN81_in4 <= VN_sign_in(490) & VN_data_in(490);
  VN81_in5 <= VN_sign_in(491) & VN_data_in(491);
  VN82_in0 <= VN_sign_in(492) & VN_data_in(492);
  VN82_in1 <= VN_sign_in(493) & VN_data_in(493);
  VN82_in2 <= VN_sign_in(494) & VN_data_in(494);
  VN82_in3 <= VN_sign_in(495) & VN_data_in(495);
  VN82_in4 <= VN_sign_in(496) & VN_data_in(496);
  VN82_in5 <= VN_sign_in(497) & VN_data_in(497);
  VN83_in0 <= VN_sign_in(498) & VN_data_in(498);
  VN83_in1 <= VN_sign_in(499) & VN_data_in(499);
  VN83_in2 <= VN_sign_in(500) & VN_data_in(500);
  VN83_in3 <= VN_sign_in(501) & VN_data_in(501);
  VN83_in4 <= VN_sign_in(502) & VN_data_in(502);
  VN83_in5 <= VN_sign_in(503) & VN_data_in(503);
  VN84_in0 <= VN_sign_in(504) & VN_data_in(504);
  VN84_in1 <= VN_sign_in(505) & VN_data_in(505);
  VN84_in2 <= VN_sign_in(506) & VN_data_in(506);
  VN84_in3 <= VN_sign_in(507) & VN_data_in(507);
  VN84_in4 <= VN_sign_in(508) & VN_data_in(508);
  VN84_in5 <= VN_sign_in(509) & VN_data_in(509);
  VN85_in0 <= VN_sign_in(510) & VN_data_in(510);
  VN85_in1 <= VN_sign_in(511) & VN_data_in(511);
  VN85_in2 <= VN_sign_in(512) & VN_data_in(512);
  VN85_in3 <= VN_sign_in(513) & VN_data_in(513);
  VN85_in4 <= VN_sign_in(514) & VN_data_in(514);
  VN85_in5 <= VN_sign_in(515) & VN_data_in(515);
  VN86_in0 <= VN_sign_in(516) & VN_data_in(516);
  VN86_in1 <= VN_sign_in(517) & VN_data_in(517);
  VN86_in2 <= VN_sign_in(518) & VN_data_in(518);
  VN86_in3 <= VN_sign_in(519) & VN_data_in(519);
  VN86_in4 <= VN_sign_in(520) & VN_data_in(520);
  VN86_in5 <= VN_sign_in(521) & VN_data_in(521);
  VN87_in0 <= VN_sign_in(522) & VN_data_in(522);
  VN87_in1 <= VN_sign_in(523) & VN_data_in(523);
  VN87_in2 <= VN_sign_in(524) & VN_data_in(524);
  VN87_in3 <= VN_sign_in(525) & VN_data_in(525);
  VN87_in4 <= VN_sign_in(526) & VN_data_in(526);
  VN87_in5 <= VN_sign_in(527) & VN_data_in(527);
  VN88_in0 <= VN_sign_in(528) & VN_data_in(528);
  VN88_in1 <= VN_sign_in(529) & VN_data_in(529);
  VN88_in2 <= VN_sign_in(530) & VN_data_in(530);
  VN88_in3 <= VN_sign_in(531) & VN_data_in(531);
  VN88_in4 <= VN_sign_in(532) & VN_data_in(532);
  VN88_in5 <= VN_sign_in(533) & VN_data_in(533);
  VN89_in0 <= VN_sign_in(534) & VN_data_in(534);
  VN89_in1 <= VN_sign_in(535) & VN_data_in(535);
  VN89_in2 <= VN_sign_in(536) & VN_data_in(536);
  VN89_in3 <= VN_sign_in(537) & VN_data_in(537);
  VN89_in4 <= VN_sign_in(538) & VN_data_in(538);
  VN89_in5 <= VN_sign_in(539) & VN_data_in(539);
  VN90_in0 <= VN_sign_in(540) & VN_data_in(540);
  VN90_in1 <= VN_sign_in(541) & VN_data_in(541);
  VN90_in2 <= VN_sign_in(542) & VN_data_in(542);
  VN90_in3 <= VN_sign_in(543) & VN_data_in(543);
  VN90_in4 <= VN_sign_in(544) & VN_data_in(544);
  VN90_in5 <= VN_sign_in(545) & VN_data_in(545);
  VN91_in0 <= VN_sign_in(546) & VN_data_in(546);
  VN91_in1 <= VN_sign_in(547) & VN_data_in(547);
  VN91_in2 <= VN_sign_in(548) & VN_data_in(548);
  VN91_in3 <= VN_sign_in(549) & VN_data_in(549);
  VN91_in4 <= VN_sign_in(550) & VN_data_in(550);
  VN91_in5 <= VN_sign_in(551) & VN_data_in(551);
  VN92_in0 <= VN_sign_in(552) & VN_data_in(552);
  VN92_in1 <= VN_sign_in(553) & VN_data_in(553);
  VN92_in2 <= VN_sign_in(554) & VN_data_in(554);
  VN92_in3 <= VN_sign_in(555) & VN_data_in(555);
  VN92_in4 <= VN_sign_in(556) & VN_data_in(556);
  VN92_in5 <= VN_sign_in(557) & VN_data_in(557);
  VN93_in0 <= VN_sign_in(558) & VN_data_in(558);
  VN93_in1 <= VN_sign_in(559) & VN_data_in(559);
  VN93_in2 <= VN_sign_in(560) & VN_data_in(560);
  VN93_in3 <= VN_sign_in(561) & VN_data_in(561);
  VN93_in4 <= VN_sign_in(562) & VN_data_in(562);
  VN93_in5 <= VN_sign_in(563) & VN_data_in(563);
  VN94_in0 <= VN_sign_in(564) & VN_data_in(564);
  VN94_in1 <= VN_sign_in(565) & VN_data_in(565);
  VN94_in2 <= VN_sign_in(566) & VN_data_in(566);
  VN94_in3 <= VN_sign_in(567) & VN_data_in(567);
  VN94_in4 <= VN_sign_in(568) & VN_data_in(568);
  VN94_in5 <= VN_sign_in(569) & VN_data_in(569);
  VN95_in0 <= VN_sign_in(570) & VN_data_in(570);
  VN95_in1 <= VN_sign_in(571) & VN_data_in(571);
  VN95_in2 <= VN_sign_in(572) & VN_data_in(572);
  VN95_in3 <= VN_sign_in(573) & VN_data_in(573);
  VN95_in4 <= VN_sign_in(574) & VN_data_in(574);
  VN95_in5 <= VN_sign_in(575) & VN_data_in(575);
  VN96_in0 <= VN_sign_in(576) & VN_data_in(576);
  VN96_in1 <= VN_sign_in(577) & VN_data_in(577);
  VN96_in2 <= VN_sign_in(578) & VN_data_in(578);
  VN96_in3 <= VN_sign_in(579) & VN_data_in(579);
  VN96_in4 <= VN_sign_in(580) & VN_data_in(580);
  VN96_in5 <= VN_sign_in(581) & VN_data_in(581);
  VN97_in0 <= VN_sign_in(582) & VN_data_in(582);
  VN97_in1 <= VN_sign_in(583) & VN_data_in(583);
  VN97_in2 <= VN_sign_in(584) & VN_data_in(584);
  VN97_in3 <= VN_sign_in(585) & VN_data_in(585);
  VN97_in4 <= VN_sign_in(586) & VN_data_in(586);
  VN97_in5 <= VN_sign_in(587) & VN_data_in(587);
  VN98_in0 <= VN_sign_in(588) & VN_data_in(588);
  VN98_in1 <= VN_sign_in(589) & VN_data_in(589);
  VN98_in2 <= VN_sign_in(590) & VN_data_in(590);
  VN98_in3 <= VN_sign_in(591) & VN_data_in(591);
  VN98_in4 <= VN_sign_in(592) & VN_data_in(592);
  VN98_in5 <= VN_sign_in(593) & VN_data_in(593);
  VN99_in0 <= VN_sign_in(594) & VN_data_in(594);
  VN99_in1 <= VN_sign_in(595) & VN_data_in(595);
  VN99_in2 <= VN_sign_in(596) & VN_data_in(596);
  VN99_in3 <= VN_sign_in(597) & VN_data_in(597);
  VN99_in4 <= VN_sign_in(598) & VN_data_in(598);
  VN99_in5 <= VN_sign_in(599) & VN_data_in(599);
  VN100_in0 <= VN_sign_in(600) & VN_data_in(600);
  VN100_in1 <= VN_sign_in(601) & VN_data_in(601);
  VN100_in2 <= VN_sign_in(602) & VN_data_in(602);
  VN100_in3 <= VN_sign_in(603) & VN_data_in(603);
  VN100_in4 <= VN_sign_in(604) & VN_data_in(604);
  VN100_in5 <= VN_sign_in(605) & VN_data_in(605);
  VN101_in0 <= VN_sign_in(606) & VN_data_in(606);
  VN101_in1 <= VN_sign_in(607) & VN_data_in(607);
  VN101_in2 <= VN_sign_in(608) & VN_data_in(608);
  VN101_in3 <= VN_sign_in(609) & VN_data_in(609);
  VN101_in4 <= VN_sign_in(610) & VN_data_in(610);
  VN101_in5 <= VN_sign_in(611) & VN_data_in(611);
  VN102_in0 <= VN_sign_in(612) & VN_data_in(612);
  VN102_in1 <= VN_sign_in(613) & VN_data_in(613);
  VN102_in2 <= VN_sign_in(614) & VN_data_in(614);
  VN102_in3 <= VN_sign_in(615) & VN_data_in(615);
  VN102_in4 <= VN_sign_in(616) & VN_data_in(616);
  VN102_in5 <= VN_sign_in(617) & VN_data_in(617);
  VN103_in0 <= VN_sign_in(618) & VN_data_in(618);
  VN103_in1 <= VN_sign_in(619) & VN_data_in(619);
  VN103_in2 <= VN_sign_in(620) & VN_data_in(620);
  VN103_in3 <= VN_sign_in(621) & VN_data_in(621);
  VN103_in4 <= VN_sign_in(622) & VN_data_in(622);
  VN103_in5 <= VN_sign_in(623) & VN_data_in(623);
  VN104_in0 <= VN_sign_in(624) & VN_data_in(624);
  VN104_in1 <= VN_sign_in(625) & VN_data_in(625);
  VN104_in2 <= VN_sign_in(626) & VN_data_in(626);
  VN104_in3 <= VN_sign_in(627) & VN_data_in(627);
  VN104_in4 <= VN_sign_in(628) & VN_data_in(628);
  VN104_in5 <= VN_sign_in(629) & VN_data_in(629);
  VN105_in0 <= VN_sign_in(630) & VN_data_in(630);
  VN105_in1 <= VN_sign_in(631) & VN_data_in(631);
  VN105_in2 <= VN_sign_in(632) & VN_data_in(632);
  VN105_in3 <= VN_sign_in(633) & VN_data_in(633);
  VN105_in4 <= VN_sign_in(634) & VN_data_in(634);
  VN105_in5 <= VN_sign_in(635) & VN_data_in(635);
  VN106_in0 <= VN_sign_in(636) & VN_data_in(636);
  VN106_in1 <= VN_sign_in(637) & VN_data_in(637);
  VN106_in2 <= VN_sign_in(638) & VN_data_in(638);
  VN106_in3 <= VN_sign_in(639) & VN_data_in(639);
  VN106_in4 <= VN_sign_in(640) & VN_data_in(640);
  VN106_in5 <= VN_sign_in(641) & VN_data_in(641);
  VN107_in0 <= VN_sign_in(642) & VN_data_in(642);
  VN107_in1 <= VN_sign_in(643) & VN_data_in(643);
  VN107_in2 <= VN_sign_in(644) & VN_data_in(644);
  VN107_in3 <= VN_sign_in(645) & VN_data_in(645);
  VN107_in4 <= VN_sign_in(646) & VN_data_in(646);
  VN107_in5 <= VN_sign_in(647) & VN_data_in(647);
  VN108_in0 <= VN_sign_in(648) & VN_data_in(648);
  VN108_in1 <= VN_sign_in(649) & VN_data_in(649);
  VN108_in2 <= VN_sign_in(650) & VN_data_in(650);
  VN108_in3 <= VN_sign_in(651) & VN_data_in(651);
  VN108_in4 <= VN_sign_in(652) & VN_data_in(652);
  VN108_in5 <= VN_sign_in(653) & VN_data_in(653);
  VN109_in0 <= VN_sign_in(654) & VN_data_in(654);
  VN109_in1 <= VN_sign_in(655) & VN_data_in(655);
  VN109_in2 <= VN_sign_in(656) & VN_data_in(656);
  VN109_in3 <= VN_sign_in(657) & VN_data_in(657);
  VN109_in4 <= VN_sign_in(658) & VN_data_in(658);
  VN109_in5 <= VN_sign_in(659) & VN_data_in(659);
  VN110_in0 <= VN_sign_in(660) & VN_data_in(660);
  VN110_in1 <= VN_sign_in(661) & VN_data_in(661);
  VN110_in2 <= VN_sign_in(662) & VN_data_in(662);
  VN110_in3 <= VN_sign_in(663) & VN_data_in(663);
  VN110_in4 <= VN_sign_in(664) & VN_data_in(664);
  VN110_in5 <= VN_sign_in(665) & VN_data_in(665);
  VN111_in0 <= VN_sign_in(666) & VN_data_in(666);
  VN111_in1 <= VN_sign_in(667) & VN_data_in(667);
  VN111_in2 <= VN_sign_in(668) & VN_data_in(668);
  VN111_in3 <= VN_sign_in(669) & VN_data_in(669);
  VN111_in4 <= VN_sign_in(670) & VN_data_in(670);
  VN111_in5 <= VN_sign_in(671) & VN_data_in(671);
  VN112_in0 <= VN_sign_in(672) & VN_data_in(672);
  VN112_in1 <= VN_sign_in(673) & VN_data_in(673);
  VN112_in2 <= VN_sign_in(674) & VN_data_in(674);
  VN112_in3 <= VN_sign_in(675) & VN_data_in(675);
  VN112_in4 <= VN_sign_in(676) & VN_data_in(676);
  VN112_in5 <= VN_sign_in(677) & VN_data_in(677);
  VN113_in0 <= VN_sign_in(678) & VN_data_in(678);
  VN113_in1 <= VN_sign_in(679) & VN_data_in(679);
  VN113_in2 <= VN_sign_in(680) & VN_data_in(680);
  VN113_in3 <= VN_sign_in(681) & VN_data_in(681);
  VN113_in4 <= VN_sign_in(682) & VN_data_in(682);
  VN113_in5 <= VN_sign_in(683) & VN_data_in(683);
  VN114_in0 <= VN_sign_in(684) & VN_data_in(684);
  VN114_in1 <= VN_sign_in(685) & VN_data_in(685);
  VN114_in2 <= VN_sign_in(686) & VN_data_in(686);
  VN114_in3 <= VN_sign_in(687) & VN_data_in(687);
  VN114_in4 <= VN_sign_in(688) & VN_data_in(688);
  VN114_in5 <= VN_sign_in(689) & VN_data_in(689);
  VN115_in0 <= VN_sign_in(690) & VN_data_in(690);
  VN115_in1 <= VN_sign_in(691) & VN_data_in(691);
  VN115_in2 <= VN_sign_in(692) & VN_data_in(692);
  VN115_in3 <= VN_sign_in(693) & VN_data_in(693);
  VN115_in4 <= VN_sign_in(694) & VN_data_in(694);
  VN115_in5 <= VN_sign_in(695) & VN_data_in(695);
  VN116_in0 <= VN_sign_in(696) & VN_data_in(696);
  VN116_in1 <= VN_sign_in(697) & VN_data_in(697);
  VN116_in2 <= VN_sign_in(698) & VN_data_in(698);
  VN116_in3 <= VN_sign_in(699) & VN_data_in(699);
  VN116_in4 <= VN_sign_in(700) & VN_data_in(700);
  VN116_in5 <= VN_sign_in(701) & VN_data_in(701);
  VN117_in0 <= VN_sign_in(702) & VN_data_in(702);
  VN117_in1 <= VN_sign_in(703) & VN_data_in(703);
  VN117_in2 <= VN_sign_in(704) & VN_data_in(704);
  VN117_in3 <= VN_sign_in(705) & VN_data_in(705);
  VN117_in4 <= VN_sign_in(706) & VN_data_in(706);
  VN117_in5 <= VN_sign_in(707) & VN_data_in(707);
  VN118_in0 <= VN_sign_in(708) & VN_data_in(708);
  VN118_in1 <= VN_sign_in(709) & VN_data_in(709);
  VN118_in2 <= VN_sign_in(710) & VN_data_in(710);
  VN118_in3 <= VN_sign_in(711) & VN_data_in(711);
  VN118_in4 <= VN_sign_in(712) & VN_data_in(712);
  VN118_in5 <= VN_sign_in(713) & VN_data_in(713);
  VN119_in0 <= VN_sign_in(714) & VN_data_in(714);
  VN119_in1 <= VN_sign_in(715) & VN_data_in(715);
  VN119_in2 <= VN_sign_in(716) & VN_data_in(716);
  VN119_in3 <= VN_sign_in(717) & VN_data_in(717);
  VN119_in4 <= VN_sign_in(718) & VN_data_in(718);
  VN119_in5 <= VN_sign_in(719) & VN_data_in(719);
  VN120_in0 <= VN_sign_in(720) & VN_data_in(720);
  VN120_in1 <= VN_sign_in(721) & VN_data_in(721);
  VN120_in2 <= VN_sign_in(722) & VN_data_in(722);
  VN120_in3 <= VN_sign_in(723) & VN_data_in(723);
  VN120_in4 <= VN_sign_in(724) & VN_data_in(724);
  VN120_in5 <= VN_sign_in(725) & VN_data_in(725);
  VN121_in0 <= VN_sign_in(726) & VN_data_in(726);
  VN121_in1 <= VN_sign_in(727) & VN_data_in(727);
  VN121_in2 <= VN_sign_in(728) & VN_data_in(728);
  VN121_in3 <= VN_sign_in(729) & VN_data_in(729);
  VN121_in4 <= VN_sign_in(730) & VN_data_in(730);
  VN121_in5 <= VN_sign_in(731) & VN_data_in(731);
  VN122_in0 <= VN_sign_in(732) & VN_data_in(732);
  VN122_in1 <= VN_sign_in(733) & VN_data_in(733);
  VN122_in2 <= VN_sign_in(734) & VN_data_in(734);
  VN122_in3 <= VN_sign_in(735) & VN_data_in(735);
  VN122_in4 <= VN_sign_in(736) & VN_data_in(736);
  VN122_in5 <= VN_sign_in(737) & VN_data_in(737);
  VN123_in0 <= VN_sign_in(738) & VN_data_in(738);
  VN123_in1 <= VN_sign_in(739) & VN_data_in(739);
  VN123_in2 <= VN_sign_in(740) & VN_data_in(740);
  VN123_in3 <= VN_sign_in(741) & VN_data_in(741);
  VN123_in4 <= VN_sign_in(742) & VN_data_in(742);
  VN123_in5 <= VN_sign_in(743) & VN_data_in(743);
  VN124_in0 <= VN_sign_in(744) & VN_data_in(744);
  VN124_in1 <= VN_sign_in(745) & VN_data_in(745);
  VN124_in2 <= VN_sign_in(746) & VN_data_in(746);
  VN124_in3 <= VN_sign_in(747) & VN_data_in(747);
  VN124_in4 <= VN_sign_in(748) & VN_data_in(748);
  VN124_in5 <= VN_sign_in(749) & VN_data_in(749);
  VN125_in0 <= VN_sign_in(750) & VN_data_in(750);
  VN125_in1 <= VN_sign_in(751) & VN_data_in(751);
  VN125_in2 <= VN_sign_in(752) & VN_data_in(752);
  VN125_in3 <= VN_sign_in(753) & VN_data_in(753);
  VN125_in4 <= VN_sign_in(754) & VN_data_in(754);
  VN125_in5 <= VN_sign_in(755) & VN_data_in(755);
  VN126_in0 <= VN_sign_in(756) & VN_data_in(756);
  VN126_in1 <= VN_sign_in(757) & VN_data_in(757);
  VN126_in2 <= VN_sign_in(758) & VN_data_in(758);
  VN126_in3 <= VN_sign_in(759) & VN_data_in(759);
  VN126_in4 <= VN_sign_in(760) & VN_data_in(760);
  VN126_in5 <= VN_sign_in(761) & VN_data_in(761);
  VN127_in0 <= VN_sign_in(762) & VN_data_in(762);
  VN127_in1 <= VN_sign_in(763) & VN_data_in(763);
  VN127_in2 <= VN_sign_in(764) & VN_data_in(764);
  VN127_in3 <= VN_sign_in(765) & VN_data_in(765);
  VN127_in4 <= VN_sign_in(766) & VN_data_in(766);
  VN127_in5 <= VN_sign_in(767) & VN_data_in(767);
  VN128_in0 <= VN_sign_in(768) & VN_data_in(768);
  VN128_in1 <= VN_sign_in(769) & VN_data_in(769);
  VN128_in2 <= VN_sign_in(770) & VN_data_in(770);
  VN128_in3 <= VN_sign_in(771) & VN_data_in(771);
  VN128_in4 <= VN_sign_in(772) & VN_data_in(772);
  VN128_in5 <= VN_sign_in(773) & VN_data_in(773);
  VN129_in0 <= VN_sign_in(774) & VN_data_in(774);
  VN129_in1 <= VN_sign_in(775) & VN_data_in(775);
  VN129_in2 <= VN_sign_in(776) & VN_data_in(776);
  VN129_in3 <= VN_sign_in(777) & VN_data_in(777);
  VN129_in4 <= VN_sign_in(778) & VN_data_in(778);
  VN129_in5 <= VN_sign_in(779) & VN_data_in(779);
  VN130_in0 <= VN_sign_in(780) & VN_data_in(780);
  VN130_in1 <= VN_sign_in(781) & VN_data_in(781);
  VN130_in2 <= VN_sign_in(782) & VN_data_in(782);
  VN130_in3 <= VN_sign_in(783) & VN_data_in(783);
  VN130_in4 <= VN_sign_in(784) & VN_data_in(784);
  VN130_in5 <= VN_sign_in(785) & VN_data_in(785);
  VN131_in0 <= VN_sign_in(786) & VN_data_in(786);
  VN131_in1 <= VN_sign_in(787) & VN_data_in(787);
  VN131_in2 <= VN_sign_in(788) & VN_data_in(788);
  VN131_in3 <= VN_sign_in(789) & VN_data_in(789);
  VN131_in4 <= VN_sign_in(790) & VN_data_in(790);
  VN131_in5 <= VN_sign_in(791) & VN_data_in(791);
  VN132_in0 <= VN_sign_in(792) & VN_data_in(792);
  VN132_in1 <= VN_sign_in(793) & VN_data_in(793);
  VN132_in2 <= VN_sign_in(794) & VN_data_in(794);
  VN132_in3 <= VN_sign_in(795) & VN_data_in(795);
  VN132_in4 <= VN_sign_in(796) & VN_data_in(796);
  VN132_in5 <= VN_sign_in(797) & VN_data_in(797);
  VN133_in0 <= VN_sign_in(798) & VN_data_in(798);
  VN133_in1 <= VN_sign_in(799) & VN_data_in(799);
  VN133_in2 <= VN_sign_in(800) & VN_data_in(800);
  VN133_in3 <= VN_sign_in(801) & VN_data_in(801);
  VN133_in4 <= VN_sign_in(802) & VN_data_in(802);
  VN133_in5 <= VN_sign_in(803) & VN_data_in(803);
  VN134_in0 <= VN_sign_in(804) & VN_data_in(804);
  VN134_in1 <= VN_sign_in(805) & VN_data_in(805);
  VN134_in2 <= VN_sign_in(806) & VN_data_in(806);
  VN134_in3 <= VN_sign_in(807) & VN_data_in(807);
  VN134_in4 <= VN_sign_in(808) & VN_data_in(808);
  VN134_in5 <= VN_sign_in(809) & VN_data_in(809);
  VN135_in0 <= VN_sign_in(810) & VN_data_in(810);
  VN135_in1 <= VN_sign_in(811) & VN_data_in(811);
  VN135_in2 <= VN_sign_in(812) & VN_data_in(812);
  VN135_in3 <= VN_sign_in(813) & VN_data_in(813);
  VN135_in4 <= VN_sign_in(814) & VN_data_in(814);
  VN135_in5 <= VN_sign_in(815) & VN_data_in(815);
  VN136_in0 <= VN_sign_in(816) & VN_data_in(816);
  VN136_in1 <= VN_sign_in(817) & VN_data_in(817);
  VN136_in2 <= VN_sign_in(818) & VN_data_in(818);
  VN136_in3 <= VN_sign_in(819) & VN_data_in(819);
  VN136_in4 <= VN_sign_in(820) & VN_data_in(820);
  VN136_in5 <= VN_sign_in(821) & VN_data_in(821);
  VN137_in0 <= VN_sign_in(822) & VN_data_in(822);
  VN137_in1 <= VN_sign_in(823) & VN_data_in(823);
  VN137_in2 <= VN_sign_in(824) & VN_data_in(824);
  VN137_in3 <= VN_sign_in(825) & VN_data_in(825);
  VN137_in4 <= VN_sign_in(826) & VN_data_in(826);
  VN137_in5 <= VN_sign_in(827) & VN_data_in(827);
  VN138_in0 <= VN_sign_in(828) & VN_data_in(828);
  VN138_in1 <= VN_sign_in(829) & VN_data_in(829);
  VN138_in2 <= VN_sign_in(830) & VN_data_in(830);
  VN138_in3 <= VN_sign_in(831) & VN_data_in(831);
  VN138_in4 <= VN_sign_in(832) & VN_data_in(832);
  VN138_in5 <= VN_sign_in(833) & VN_data_in(833);
  VN139_in0 <= VN_sign_in(834) & VN_data_in(834);
  VN139_in1 <= VN_sign_in(835) & VN_data_in(835);
  VN139_in2 <= VN_sign_in(836) & VN_data_in(836);
  VN139_in3 <= VN_sign_in(837) & VN_data_in(837);
  VN139_in4 <= VN_sign_in(838) & VN_data_in(838);
  VN139_in5 <= VN_sign_in(839) & VN_data_in(839);
  VN140_in0 <= VN_sign_in(840) & VN_data_in(840);
  VN140_in1 <= VN_sign_in(841) & VN_data_in(841);
  VN140_in2 <= VN_sign_in(842) & VN_data_in(842);
  VN140_in3 <= VN_sign_in(843) & VN_data_in(843);
  VN140_in4 <= VN_sign_in(844) & VN_data_in(844);
  VN140_in5 <= VN_sign_in(845) & VN_data_in(845);
  VN141_in0 <= VN_sign_in(846) & VN_data_in(846);
  VN141_in1 <= VN_sign_in(847) & VN_data_in(847);
  VN141_in2 <= VN_sign_in(848) & VN_data_in(848);
  VN141_in3 <= VN_sign_in(849) & VN_data_in(849);
  VN141_in4 <= VN_sign_in(850) & VN_data_in(850);
  VN141_in5 <= VN_sign_in(851) & VN_data_in(851);
  VN142_in0 <= VN_sign_in(852) & VN_data_in(852);
  VN142_in1 <= VN_sign_in(853) & VN_data_in(853);
  VN142_in2 <= VN_sign_in(854) & VN_data_in(854);
  VN142_in3 <= VN_sign_in(855) & VN_data_in(855);
  VN142_in4 <= VN_sign_in(856) & VN_data_in(856);
  VN142_in5 <= VN_sign_in(857) & VN_data_in(857);
  VN143_in0 <= VN_sign_in(858) & VN_data_in(858);
  VN143_in1 <= VN_sign_in(859) & VN_data_in(859);
  VN143_in2 <= VN_sign_in(860) & VN_data_in(860);
  VN143_in3 <= VN_sign_in(861) & VN_data_in(861);
  VN143_in4 <= VN_sign_in(862) & VN_data_in(862);
  VN143_in5 <= VN_sign_in(863) & VN_data_in(863);
  VN144_in0 <= VN_sign_in(864) & VN_data_in(864);
  VN144_in1 <= VN_sign_in(865) & VN_data_in(865);
  VN144_in2 <= VN_sign_in(866) & VN_data_in(866);
  VN144_in3 <= VN_sign_in(867) & VN_data_in(867);
  VN144_in4 <= VN_sign_in(868) & VN_data_in(868);
  VN144_in5 <= VN_sign_in(869) & VN_data_in(869);
  VN145_in0 <= VN_sign_in(870) & VN_data_in(870);
  VN145_in1 <= VN_sign_in(871) & VN_data_in(871);
  VN145_in2 <= VN_sign_in(872) & VN_data_in(872);
  VN145_in3 <= VN_sign_in(873) & VN_data_in(873);
  VN145_in4 <= VN_sign_in(874) & VN_data_in(874);
  VN145_in5 <= VN_sign_in(875) & VN_data_in(875);
  VN146_in0 <= VN_sign_in(876) & VN_data_in(876);
  VN146_in1 <= VN_sign_in(877) & VN_data_in(877);
  VN146_in2 <= VN_sign_in(878) & VN_data_in(878);
  VN146_in3 <= VN_sign_in(879) & VN_data_in(879);
  VN146_in4 <= VN_sign_in(880) & VN_data_in(880);
  VN146_in5 <= VN_sign_in(881) & VN_data_in(881);
  VN147_in0 <= VN_sign_in(882) & VN_data_in(882);
  VN147_in1 <= VN_sign_in(883) & VN_data_in(883);
  VN147_in2 <= VN_sign_in(884) & VN_data_in(884);
  VN147_in3 <= VN_sign_in(885) & VN_data_in(885);
  VN147_in4 <= VN_sign_in(886) & VN_data_in(886);
  VN147_in5 <= VN_sign_in(887) & VN_data_in(887);
  VN148_in0 <= VN_sign_in(888) & VN_data_in(888);
  VN148_in1 <= VN_sign_in(889) & VN_data_in(889);
  VN148_in2 <= VN_sign_in(890) & VN_data_in(890);
  VN148_in3 <= VN_sign_in(891) & VN_data_in(891);
  VN148_in4 <= VN_sign_in(892) & VN_data_in(892);
  VN148_in5 <= VN_sign_in(893) & VN_data_in(893);
  VN149_in0 <= VN_sign_in(894) & VN_data_in(894);
  VN149_in1 <= VN_sign_in(895) & VN_data_in(895);
  VN149_in2 <= VN_sign_in(896) & VN_data_in(896);
  VN149_in3 <= VN_sign_in(897) & VN_data_in(897);
  VN149_in4 <= VN_sign_in(898) & VN_data_in(898);
  VN149_in5 <= VN_sign_in(899) & VN_data_in(899);
  VN150_in0 <= VN_sign_in(900) & VN_data_in(900);
  VN150_in1 <= VN_sign_in(901) & VN_data_in(901);
  VN150_in2 <= VN_sign_in(902) & VN_data_in(902);
  VN150_in3 <= VN_sign_in(903) & VN_data_in(903);
  VN150_in4 <= VN_sign_in(904) & VN_data_in(904);
  VN150_in5 <= VN_sign_in(905) & VN_data_in(905);
  VN151_in0 <= VN_sign_in(906) & VN_data_in(906);
  VN151_in1 <= VN_sign_in(907) & VN_data_in(907);
  VN151_in2 <= VN_sign_in(908) & VN_data_in(908);
  VN151_in3 <= VN_sign_in(909) & VN_data_in(909);
  VN151_in4 <= VN_sign_in(910) & VN_data_in(910);
  VN151_in5 <= VN_sign_in(911) & VN_data_in(911);
  VN152_in0 <= VN_sign_in(912) & VN_data_in(912);
  VN152_in1 <= VN_sign_in(913) & VN_data_in(913);
  VN152_in2 <= VN_sign_in(914) & VN_data_in(914);
  VN152_in3 <= VN_sign_in(915) & VN_data_in(915);
  VN152_in4 <= VN_sign_in(916) & VN_data_in(916);
  VN152_in5 <= VN_sign_in(917) & VN_data_in(917);
  VN153_in0 <= VN_sign_in(918) & VN_data_in(918);
  VN153_in1 <= VN_sign_in(919) & VN_data_in(919);
  VN153_in2 <= VN_sign_in(920) & VN_data_in(920);
  VN153_in3 <= VN_sign_in(921) & VN_data_in(921);
  VN153_in4 <= VN_sign_in(922) & VN_data_in(922);
  VN153_in5 <= VN_sign_in(923) & VN_data_in(923);
  VN154_in0 <= VN_sign_in(924) & VN_data_in(924);
  VN154_in1 <= VN_sign_in(925) & VN_data_in(925);
  VN154_in2 <= VN_sign_in(926) & VN_data_in(926);
  VN154_in3 <= VN_sign_in(927) & VN_data_in(927);
  VN154_in4 <= VN_sign_in(928) & VN_data_in(928);
  VN154_in5 <= VN_sign_in(929) & VN_data_in(929);
  VN155_in0 <= VN_sign_in(930) & VN_data_in(930);
  VN155_in1 <= VN_sign_in(931) & VN_data_in(931);
  VN155_in2 <= VN_sign_in(932) & VN_data_in(932);
  VN155_in3 <= VN_sign_in(933) & VN_data_in(933);
  VN155_in4 <= VN_sign_in(934) & VN_data_in(934);
  VN155_in5 <= VN_sign_in(935) & VN_data_in(935);
  VN156_in0 <= VN_sign_in(936) & VN_data_in(936);
  VN156_in1 <= VN_sign_in(937) & VN_data_in(937);
  VN156_in2 <= VN_sign_in(938) & VN_data_in(938);
  VN156_in3 <= VN_sign_in(939) & VN_data_in(939);
  VN156_in4 <= VN_sign_in(940) & VN_data_in(940);
  VN156_in5 <= VN_sign_in(941) & VN_data_in(941);
  VN157_in0 <= VN_sign_in(942) & VN_data_in(942);
  VN157_in1 <= VN_sign_in(943) & VN_data_in(943);
  VN157_in2 <= VN_sign_in(944) & VN_data_in(944);
  VN157_in3 <= VN_sign_in(945) & VN_data_in(945);
  VN157_in4 <= VN_sign_in(946) & VN_data_in(946);
  VN157_in5 <= VN_sign_in(947) & VN_data_in(947);
  VN158_in0 <= VN_sign_in(948) & VN_data_in(948);
  VN158_in1 <= VN_sign_in(949) & VN_data_in(949);
  VN158_in2 <= VN_sign_in(950) & VN_data_in(950);
  VN158_in3 <= VN_sign_in(951) & VN_data_in(951);
  VN158_in4 <= VN_sign_in(952) & VN_data_in(952);
  VN158_in5 <= VN_sign_in(953) & VN_data_in(953);
  VN159_in0 <= VN_sign_in(954) & VN_data_in(954);
  VN159_in1 <= VN_sign_in(955) & VN_data_in(955);
  VN159_in2 <= VN_sign_in(956) & VN_data_in(956);
  VN159_in3 <= VN_sign_in(957) & VN_data_in(957);
  VN159_in4 <= VN_sign_in(958) & VN_data_in(958);
  VN159_in5 <= VN_sign_in(959) & VN_data_in(959);
  VN160_in0 <= VN_sign_in(960) & VN_data_in(960);
  VN160_in1 <= VN_sign_in(961) & VN_data_in(961);
  VN160_in2 <= VN_sign_in(962) & VN_data_in(962);
  VN160_in3 <= VN_sign_in(963) & VN_data_in(963);
  VN160_in4 <= VN_sign_in(964) & VN_data_in(964);
  VN160_in5 <= VN_sign_in(965) & VN_data_in(965);
  VN161_in0 <= VN_sign_in(966) & VN_data_in(966);
  VN161_in1 <= VN_sign_in(967) & VN_data_in(967);
  VN161_in2 <= VN_sign_in(968) & VN_data_in(968);
  VN161_in3 <= VN_sign_in(969) & VN_data_in(969);
  VN161_in4 <= VN_sign_in(970) & VN_data_in(970);
  VN161_in5 <= VN_sign_in(971) & VN_data_in(971);
  VN162_in0 <= VN_sign_in(972) & VN_data_in(972);
  VN162_in1 <= VN_sign_in(973) & VN_data_in(973);
  VN162_in2 <= VN_sign_in(974) & VN_data_in(974);
  VN162_in3 <= VN_sign_in(975) & VN_data_in(975);
  VN162_in4 <= VN_sign_in(976) & VN_data_in(976);
  VN162_in5 <= VN_sign_in(977) & VN_data_in(977);
  VN163_in0 <= VN_sign_in(978) & VN_data_in(978);
  VN163_in1 <= VN_sign_in(979) & VN_data_in(979);
  VN163_in2 <= VN_sign_in(980) & VN_data_in(980);
  VN163_in3 <= VN_sign_in(981) & VN_data_in(981);
  VN163_in4 <= VN_sign_in(982) & VN_data_in(982);
  VN163_in5 <= VN_sign_in(983) & VN_data_in(983);
  VN164_in0 <= VN_sign_in(984) & VN_data_in(984);
  VN164_in1 <= VN_sign_in(985) & VN_data_in(985);
  VN164_in2 <= VN_sign_in(986) & VN_data_in(986);
  VN164_in3 <= VN_sign_in(987) & VN_data_in(987);
  VN164_in4 <= VN_sign_in(988) & VN_data_in(988);
  VN164_in5 <= VN_sign_in(989) & VN_data_in(989);
  VN165_in0 <= VN_sign_in(990) & VN_data_in(990);
  VN165_in1 <= VN_sign_in(991) & VN_data_in(991);
  VN165_in2 <= VN_sign_in(992) & VN_data_in(992);
  VN165_in3 <= VN_sign_in(993) & VN_data_in(993);
  VN165_in4 <= VN_sign_in(994) & VN_data_in(994);
  VN165_in5 <= VN_sign_in(995) & VN_data_in(995);
  VN166_in0 <= VN_sign_in(996) & VN_data_in(996);
  VN166_in1 <= VN_sign_in(997) & VN_data_in(997);
  VN166_in2 <= VN_sign_in(998) & VN_data_in(998);
  VN166_in3 <= VN_sign_in(999) & VN_data_in(999);
  VN166_in4 <= VN_sign_in(1000) & VN_data_in(1000);
  VN166_in5 <= VN_sign_in(1001) & VN_data_in(1001);
  VN167_in0 <= VN_sign_in(1002) & VN_data_in(1002);
  VN167_in1 <= VN_sign_in(1003) & VN_data_in(1003);
  VN167_in2 <= VN_sign_in(1004) & VN_data_in(1004);
  VN167_in3 <= VN_sign_in(1005) & VN_data_in(1005);
  VN167_in4 <= VN_sign_in(1006) & VN_data_in(1006);
  VN167_in5 <= VN_sign_in(1007) & VN_data_in(1007);
  VN168_in0 <= VN_sign_in(1008) & VN_data_in(1008);
  VN168_in1 <= VN_sign_in(1009) & VN_data_in(1009);
  VN168_in2 <= VN_sign_in(1010) & VN_data_in(1010);
  VN168_in3 <= VN_sign_in(1011) & VN_data_in(1011);
  VN168_in4 <= VN_sign_in(1012) & VN_data_in(1012);
  VN168_in5 <= VN_sign_in(1013) & VN_data_in(1013);
  VN169_in0 <= VN_sign_in(1014) & VN_data_in(1014);
  VN169_in1 <= VN_sign_in(1015) & VN_data_in(1015);
  VN169_in2 <= VN_sign_in(1016) & VN_data_in(1016);
  VN169_in3 <= VN_sign_in(1017) & VN_data_in(1017);
  VN169_in4 <= VN_sign_in(1018) & VN_data_in(1018);
  VN169_in5 <= VN_sign_in(1019) & VN_data_in(1019);
  VN170_in0 <= VN_sign_in(1020) & VN_data_in(1020);
  VN170_in1 <= VN_sign_in(1021) & VN_data_in(1021);
  VN170_in2 <= VN_sign_in(1022) & VN_data_in(1022);
  VN170_in3 <= VN_sign_in(1023) & VN_data_in(1023);
  VN170_in4 <= VN_sign_in(1024) & VN_data_in(1024);
  VN170_in5 <= VN_sign_in(1025) & VN_data_in(1025);
  VN171_in0 <= VN_sign_in(1026) & VN_data_in(1026);
  VN171_in1 <= VN_sign_in(1027) & VN_data_in(1027);
  VN171_in2 <= VN_sign_in(1028) & VN_data_in(1028);
  VN171_in3 <= VN_sign_in(1029) & VN_data_in(1029);
  VN171_in4 <= VN_sign_in(1030) & VN_data_in(1030);
  VN171_in5 <= VN_sign_in(1031) & VN_data_in(1031);
  VN172_in0 <= VN_sign_in(1032) & VN_data_in(1032);
  VN172_in1 <= VN_sign_in(1033) & VN_data_in(1033);
  VN172_in2 <= VN_sign_in(1034) & VN_data_in(1034);
  VN172_in3 <= VN_sign_in(1035) & VN_data_in(1035);
  VN172_in4 <= VN_sign_in(1036) & VN_data_in(1036);
  VN172_in5 <= VN_sign_in(1037) & VN_data_in(1037);
  VN173_in0 <= VN_sign_in(1038) & VN_data_in(1038);
  VN173_in1 <= VN_sign_in(1039) & VN_data_in(1039);
  VN173_in2 <= VN_sign_in(1040) & VN_data_in(1040);
  VN173_in3 <= VN_sign_in(1041) & VN_data_in(1041);
  VN173_in4 <= VN_sign_in(1042) & VN_data_in(1042);
  VN173_in5 <= VN_sign_in(1043) & VN_data_in(1043);
  VN174_in0 <= VN_sign_in(1044) & VN_data_in(1044);
  VN174_in1 <= VN_sign_in(1045) & VN_data_in(1045);
  VN174_in2 <= VN_sign_in(1046) & VN_data_in(1046);
  VN174_in3 <= VN_sign_in(1047) & VN_data_in(1047);
  VN174_in4 <= VN_sign_in(1048) & VN_data_in(1048);
  VN174_in5 <= VN_sign_in(1049) & VN_data_in(1049);
  VN175_in0 <= VN_sign_in(1050) & VN_data_in(1050);
  VN175_in1 <= VN_sign_in(1051) & VN_data_in(1051);
  VN175_in2 <= VN_sign_in(1052) & VN_data_in(1052);
  VN175_in3 <= VN_sign_in(1053) & VN_data_in(1053);
  VN175_in4 <= VN_sign_in(1054) & VN_data_in(1054);
  VN175_in5 <= VN_sign_in(1055) & VN_data_in(1055);
  VN176_in0 <= VN_sign_in(1056) & VN_data_in(1056);
  VN176_in1 <= VN_sign_in(1057) & VN_data_in(1057);
  VN176_in2 <= VN_sign_in(1058) & VN_data_in(1058);
  VN176_in3 <= VN_sign_in(1059) & VN_data_in(1059);
  VN176_in4 <= VN_sign_in(1060) & VN_data_in(1060);
  VN176_in5 <= VN_sign_in(1061) & VN_data_in(1061);
  VN177_in0 <= VN_sign_in(1062) & VN_data_in(1062);
  VN177_in1 <= VN_sign_in(1063) & VN_data_in(1063);
  VN177_in2 <= VN_sign_in(1064) & VN_data_in(1064);
  VN177_in3 <= VN_sign_in(1065) & VN_data_in(1065);
  VN177_in4 <= VN_sign_in(1066) & VN_data_in(1066);
  VN177_in5 <= VN_sign_in(1067) & VN_data_in(1067);
  VN178_in0 <= VN_sign_in(1068) & VN_data_in(1068);
  VN178_in1 <= VN_sign_in(1069) & VN_data_in(1069);
  VN178_in2 <= VN_sign_in(1070) & VN_data_in(1070);
  VN178_in3 <= VN_sign_in(1071) & VN_data_in(1071);
  VN178_in4 <= VN_sign_in(1072) & VN_data_in(1072);
  VN178_in5 <= VN_sign_in(1073) & VN_data_in(1073);
  VN179_in0 <= VN_sign_in(1074) & VN_data_in(1074);
  VN179_in1 <= VN_sign_in(1075) & VN_data_in(1075);
  VN179_in2 <= VN_sign_in(1076) & VN_data_in(1076);
  VN179_in3 <= VN_sign_in(1077) & VN_data_in(1077);
  VN179_in4 <= VN_sign_in(1078) & VN_data_in(1078);
  VN179_in5 <= VN_sign_in(1079) & VN_data_in(1079);
  VN180_in0 <= VN_sign_in(1080) & VN_data_in(1080);
  VN180_in1 <= VN_sign_in(1081) & VN_data_in(1081);
  VN180_in2 <= VN_sign_in(1082) & VN_data_in(1082);
  VN180_in3 <= VN_sign_in(1083) & VN_data_in(1083);
  VN180_in4 <= VN_sign_in(1084) & VN_data_in(1084);
  VN180_in5 <= VN_sign_in(1085) & VN_data_in(1085);
  VN181_in0 <= VN_sign_in(1086) & VN_data_in(1086);
  VN181_in1 <= VN_sign_in(1087) & VN_data_in(1087);
  VN181_in2 <= VN_sign_in(1088) & VN_data_in(1088);
  VN181_in3 <= VN_sign_in(1089) & VN_data_in(1089);
  VN181_in4 <= VN_sign_in(1090) & VN_data_in(1090);
  VN181_in5 <= VN_sign_in(1091) & VN_data_in(1091);
  VN182_in0 <= VN_sign_in(1092) & VN_data_in(1092);
  VN182_in1 <= VN_sign_in(1093) & VN_data_in(1093);
  VN182_in2 <= VN_sign_in(1094) & VN_data_in(1094);
  VN182_in3 <= VN_sign_in(1095) & VN_data_in(1095);
  VN182_in4 <= VN_sign_in(1096) & VN_data_in(1096);
  VN182_in5 <= VN_sign_in(1097) & VN_data_in(1097);
  VN183_in0 <= VN_sign_in(1098) & VN_data_in(1098);
  VN183_in1 <= VN_sign_in(1099) & VN_data_in(1099);
  VN183_in2 <= VN_sign_in(1100) & VN_data_in(1100);
  VN183_in3 <= VN_sign_in(1101) & VN_data_in(1101);
  VN183_in4 <= VN_sign_in(1102) & VN_data_in(1102);
  VN183_in5 <= VN_sign_in(1103) & VN_data_in(1103);
  VN184_in0 <= VN_sign_in(1104) & VN_data_in(1104);
  VN184_in1 <= VN_sign_in(1105) & VN_data_in(1105);
  VN184_in2 <= VN_sign_in(1106) & VN_data_in(1106);
  VN184_in3 <= VN_sign_in(1107) & VN_data_in(1107);
  VN184_in4 <= VN_sign_in(1108) & VN_data_in(1108);
  VN184_in5 <= VN_sign_in(1109) & VN_data_in(1109);
  VN185_in0 <= VN_sign_in(1110) & VN_data_in(1110);
  VN185_in1 <= VN_sign_in(1111) & VN_data_in(1111);
  VN185_in2 <= VN_sign_in(1112) & VN_data_in(1112);
  VN185_in3 <= VN_sign_in(1113) & VN_data_in(1113);
  VN185_in4 <= VN_sign_in(1114) & VN_data_in(1114);
  VN185_in5 <= VN_sign_in(1115) & VN_data_in(1115);
  VN186_in0 <= VN_sign_in(1116) & VN_data_in(1116);
  VN186_in1 <= VN_sign_in(1117) & VN_data_in(1117);
  VN186_in2 <= VN_sign_in(1118) & VN_data_in(1118);
  VN186_in3 <= VN_sign_in(1119) & VN_data_in(1119);
  VN186_in4 <= VN_sign_in(1120) & VN_data_in(1120);
  VN186_in5 <= VN_sign_in(1121) & VN_data_in(1121);
  VN187_in0 <= VN_sign_in(1122) & VN_data_in(1122);
  VN187_in1 <= VN_sign_in(1123) & VN_data_in(1123);
  VN187_in2 <= VN_sign_in(1124) & VN_data_in(1124);
  VN187_in3 <= VN_sign_in(1125) & VN_data_in(1125);
  VN187_in4 <= VN_sign_in(1126) & VN_data_in(1126);
  VN187_in5 <= VN_sign_in(1127) & VN_data_in(1127);
  VN188_in0 <= VN_sign_in(1128) & VN_data_in(1128);
  VN188_in1 <= VN_sign_in(1129) & VN_data_in(1129);
  VN188_in2 <= VN_sign_in(1130) & VN_data_in(1130);
  VN188_in3 <= VN_sign_in(1131) & VN_data_in(1131);
  VN188_in4 <= VN_sign_in(1132) & VN_data_in(1132);
  VN188_in5 <= VN_sign_in(1133) & VN_data_in(1133);
  VN189_in0 <= VN_sign_in(1134) & VN_data_in(1134);
  VN189_in1 <= VN_sign_in(1135) & VN_data_in(1135);
  VN189_in2 <= VN_sign_in(1136) & VN_data_in(1136);
  VN189_in3 <= VN_sign_in(1137) & VN_data_in(1137);
  VN189_in4 <= VN_sign_in(1138) & VN_data_in(1138);
  VN189_in5 <= VN_sign_in(1139) & VN_data_in(1139);
  VN190_in0 <= VN_sign_in(1140) & VN_data_in(1140);
  VN190_in1 <= VN_sign_in(1141) & VN_data_in(1141);
  VN190_in2 <= VN_sign_in(1142) & VN_data_in(1142);
  VN190_in3 <= VN_sign_in(1143) & VN_data_in(1143);
  VN190_in4 <= VN_sign_in(1144) & VN_data_in(1144);
  VN190_in5 <= VN_sign_in(1145) & VN_data_in(1145);
  VN191_in0 <= VN_sign_in(1146) & VN_data_in(1146);
  VN191_in1 <= VN_sign_in(1147) & VN_data_in(1147);
  VN191_in2 <= VN_sign_in(1148) & VN_data_in(1148);
  VN191_in3 <= VN_sign_in(1149) & VN_data_in(1149);
  VN191_in4 <= VN_sign_in(1150) & VN_data_in(1150);
  VN191_in5 <= VN_sign_in(1151) & VN_data_in(1151);
  VN192_in0 <= VN_sign_in(1152) & VN_data_in(1152);
  VN192_in1 <= VN_sign_in(1153) & VN_data_in(1153);
  VN192_in2 <= VN_sign_in(1154) & VN_data_in(1154);
  VN192_in3 <= VN_sign_in(1155) & VN_data_in(1155);
  VN192_in4 <= VN_sign_in(1156) & VN_data_in(1156);
  VN192_in5 <= VN_sign_in(1157) & VN_data_in(1157);
  VN193_in0 <= VN_sign_in(1158) & VN_data_in(1158);
  VN193_in1 <= VN_sign_in(1159) & VN_data_in(1159);
  VN193_in2 <= VN_sign_in(1160) & VN_data_in(1160);
  VN193_in3 <= VN_sign_in(1161) & VN_data_in(1161);
  VN193_in4 <= VN_sign_in(1162) & VN_data_in(1162);
  VN193_in5 <= VN_sign_in(1163) & VN_data_in(1163);
  VN194_in0 <= VN_sign_in(1164) & VN_data_in(1164);
  VN194_in1 <= VN_sign_in(1165) & VN_data_in(1165);
  VN194_in2 <= VN_sign_in(1166) & VN_data_in(1166);
  VN194_in3 <= VN_sign_in(1167) & VN_data_in(1167);
  VN194_in4 <= VN_sign_in(1168) & VN_data_in(1168);
  VN194_in5 <= VN_sign_in(1169) & VN_data_in(1169);
  VN195_in0 <= VN_sign_in(1170) & VN_data_in(1170);
  VN195_in1 <= VN_sign_in(1171) & VN_data_in(1171);
  VN195_in2 <= VN_sign_in(1172) & VN_data_in(1172);
  VN195_in3 <= VN_sign_in(1173) & VN_data_in(1173);
  VN195_in4 <= VN_sign_in(1174) & VN_data_in(1174);
  VN195_in5 <= VN_sign_in(1175) & VN_data_in(1175);
  VN196_in0 <= VN_sign_in(1176) & VN_data_in(1176);
  VN196_in1 <= VN_sign_in(1177) & VN_data_in(1177);
  VN196_in2 <= VN_sign_in(1178) & VN_data_in(1178);
  VN196_in3 <= VN_sign_in(1179) & VN_data_in(1179);
  VN196_in4 <= VN_sign_in(1180) & VN_data_in(1180);
  VN196_in5 <= VN_sign_in(1181) & VN_data_in(1181);
  VN197_in0 <= VN_sign_in(1182) & VN_data_in(1182);
  VN197_in1 <= VN_sign_in(1183) & VN_data_in(1183);
  VN197_in2 <= VN_sign_in(1184) & VN_data_in(1184);
  VN197_in3 <= VN_sign_in(1185) & VN_data_in(1185);
  VN197_in4 <= VN_sign_in(1186) & VN_data_in(1186);
  VN197_in5 <= VN_sign_in(1187) & VN_data_in(1187);
  VN198_in0 <= VN_sign_in(1188) & VN_data_in(1188);
  VN198_in1 <= VN_sign_in(1189) & VN_data_in(1189);
  VN198_in2 <= VN_sign_in(1190) & VN_data_in(1190);
  VN198_in3 <= VN_sign_in(1191) & VN_data_in(1191);
  VN198_in4 <= VN_sign_in(1192) & VN_data_in(1192);
  VN198_in5 <= VN_sign_in(1193) & VN_data_in(1193);
  VN199_in0 <= VN_sign_in(1194) & VN_data_in(1194);
  VN199_in1 <= VN_sign_in(1195) & VN_data_in(1195);
  VN199_in2 <= VN_sign_in(1196) & VN_data_in(1196);
  VN199_in3 <= VN_sign_in(1197) & VN_data_in(1197);
  VN199_in4 <= VN_sign_in(1198) & VN_data_in(1198);
  VN199_in5 <= VN_sign_in(1199) & VN_data_in(1199);
  VN200_in0 <= VN_sign_in(1200) & VN_data_in(1200);
  VN200_in1 <= VN_sign_in(1201) & VN_data_in(1201);
  VN200_in2 <= VN_sign_in(1202) & VN_data_in(1202);
  VN200_in3 <= VN_sign_in(1203) & VN_data_in(1203);
  VN200_in4 <= VN_sign_in(1204) & VN_data_in(1204);
  VN200_in5 <= VN_sign_in(1205) & VN_data_in(1205);
  VN201_in0 <= VN_sign_in(1206) & VN_data_in(1206);
  VN201_in1 <= VN_sign_in(1207) & VN_data_in(1207);
  VN201_in2 <= VN_sign_in(1208) & VN_data_in(1208);
  VN201_in3 <= VN_sign_in(1209) & VN_data_in(1209);
  VN201_in4 <= VN_sign_in(1210) & VN_data_in(1210);
  VN201_in5 <= VN_sign_in(1211) & VN_data_in(1211);
  VN202_in0 <= VN_sign_in(1212) & VN_data_in(1212);
  VN202_in1 <= VN_sign_in(1213) & VN_data_in(1213);
  VN202_in2 <= VN_sign_in(1214) & VN_data_in(1214);
  VN202_in3 <= VN_sign_in(1215) & VN_data_in(1215);
  VN202_in4 <= VN_sign_in(1216) & VN_data_in(1216);
  VN202_in5 <= VN_sign_in(1217) & VN_data_in(1217);
  VN203_in0 <= VN_sign_in(1218) & VN_data_in(1218);
  VN203_in1 <= VN_sign_in(1219) & VN_data_in(1219);
  VN203_in2 <= VN_sign_in(1220) & VN_data_in(1220);
  VN203_in3 <= VN_sign_in(1221) & VN_data_in(1221);
  VN203_in4 <= VN_sign_in(1222) & VN_data_in(1222);
  VN203_in5 <= VN_sign_in(1223) & VN_data_in(1223);
  VN204_in0 <= VN_sign_in(1224) & VN_data_in(1224);
  VN204_in1 <= VN_sign_in(1225) & VN_data_in(1225);
  VN204_in2 <= VN_sign_in(1226) & VN_data_in(1226);
  VN204_in3 <= VN_sign_in(1227) & VN_data_in(1227);
  VN204_in4 <= VN_sign_in(1228) & VN_data_in(1228);
  VN204_in5 <= VN_sign_in(1229) & VN_data_in(1229);
  VN205_in0 <= VN_sign_in(1230) & VN_data_in(1230);
  VN205_in1 <= VN_sign_in(1231) & VN_data_in(1231);
  VN205_in2 <= VN_sign_in(1232) & VN_data_in(1232);
  VN205_in3 <= VN_sign_in(1233) & VN_data_in(1233);
  VN205_in4 <= VN_sign_in(1234) & VN_data_in(1234);
  VN205_in5 <= VN_sign_in(1235) & VN_data_in(1235);
  VN206_in0 <= VN_sign_in(1236) & VN_data_in(1236);
  VN206_in1 <= VN_sign_in(1237) & VN_data_in(1237);
  VN206_in2 <= VN_sign_in(1238) & VN_data_in(1238);
  VN206_in3 <= VN_sign_in(1239) & VN_data_in(1239);
  VN206_in4 <= VN_sign_in(1240) & VN_data_in(1240);
  VN206_in5 <= VN_sign_in(1241) & VN_data_in(1241);
  VN207_in0 <= VN_sign_in(1242) & VN_data_in(1242);
  VN207_in1 <= VN_sign_in(1243) & VN_data_in(1243);
  VN207_in2 <= VN_sign_in(1244) & VN_data_in(1244);
  VN207_in3 <= VN_sign_in(1245) & VN_data_in(1245);
  VN207_in4 <= VN_sign_in(1246) & VN_data_in(1246);
  VN207_in5 <= VN_sign_in(1247) & VN_data_in(1247);
  VN208_in0 <= VN_sign_in(1248) & VN_data_in(1248);
  VN208_in1 <= VN_sign_in(1249) & VN_data_in(1249);
  VN208_in2 <= VN_sign_in(1250) & VN_data_in(1250);
  VN208_in3 <= VN_sign_in(1251) & VN_data_in(1251);
  VN208_in4 <= VN_sign_in(1252) & VN_data_in(1252);
  VN208_in5 <= VN_sign_in(1253) & VN_data_in(1253);
  VN209_in0 <= VN_sign_in(1254) & VN_data_in(1254);
  VN209_in1 <= VN_sign_in(1255) & VN_data_in(1255);
  VN209_in2 <= VN_sign_in(1256) & VN_data_in(1256);
  VN209_in3 <= VN_sign_in(1257) & VN_data_in(1257);
  VN209_in4 <= VN_sign_in(1258) & VN_data_in(1258);
  VN209_in5 <= VN_sign_in(1259) & VN_data_in(1259);
  VN210_in0 <= VN_sign_in(1260) & VN_data_in(1260);
  VN210_in1 <= VN_sign_in(1261) & VN_data_in(1261);
  VN210_in2 <= VN_sign_in(1262) & VN_data_in(1262);
  VN210_in3 <= VN_sign_in(1263) & VN_data_in(1263);
  VN210_in4 <= VN_sign_in(1264) & VN_data_in(1264);
  VN210_in5 <= VN_sign_in(1265) & VN_data_in(1265);
  VN211_in0 <= VN_sign_in(1266) & VN_data_in(1266);
  VN211_in1 <= VN_sign_in(1267) & VN_data_in(1267);
  VN211_in2 <= VN_sign_in(1268) & VN_data_in(1268);
  VN211_in3 <= VN_sign_in(1269) & VN_data_in(1269);
  VN211_in4 <= VN_sign_in(1270) & VN_data_in(1270);
  VN211_in5 <= VN_sign_in(1271) & VN_data_in(1271);
  VN212_in0 <= VN_sign_in(1272) & VN_data_in(1272);
  VN212_in1 <= VN_sign_in(1273) & VN_data_in(1273);
  VN212_in2 <= VN_sign_in(1274) & VN_data_in(1274);
  VN212_in3 <= VN_sign_in(1275) & VN_data_in(1275);
  VN212_in4 <= VN_sign_in(1276) & VN_data_in(1276);
  VN212_in5 <= VN_sign_in(1277) & VN_data_in(1277);
  VN213_in0 <= VN_sign_in(1278) & VN_data_in(1278);
  VN213_in1 <= VN_sign_in(1279) & VN_data_in(1279);
  VN213_in2 <= VN_sign_in(1280) & VN_data_in(1280);
  VN213_in3 <= VN_sign_in(1281) & VN_data_in(1281);
  VN213_in4 <= VN_sign_in(1282) & VN_data_in(1282);
  VN213_in5 <= VN_sign_in(1283) & VN_data_in(1283);
  VN214_in0 <= VN_sign_in(1284) & VN_data_in(1284);
  VN214_in1 <= VN_sign_in(1285) & VN_data_in(1285);
  VN214_in2 <= VN_sign_in(1286) & VN_data_in(1286);
  VN214_in3 <= VN_sign_in(1287) & VN_data_in(1287);
  VN214_in4 <= VN_sign_in(1288) & VN_data_in(1288);
  VN214_in5 <= VN_sign_in(1289) & VN_data_in(1289);
  VN215_in0 <= VN_sign_in(1290) & VN_data_in(1290);
  VN215_in1 <= VN_sign_in(1291) & VN_data_in(1291);
  VN215_in2 <= VN_sign_in(1292) & VN_data_in(1292);
  VN215_in3 <= VN_sign_in(1293) & VN_data_in(1293);
  VN215_in4 <= VN_sign_in(1294) & VN_data_in(1294);
  VN215_in5 <= VN_sign_in(1295) & VN_data_in(1295);
  VN216_in0 <= VN_sign_in(1296) & VN_data_in(1296);
  VN216_in1 <= VN_sign_in(1297) & VN_data_in(1297);
  VN216_in2 <= VN_sign_in(1298) & VN_data_in(1298);
  VN216_in3 <= VN_sign_in(1299) & VN_data_in(1299);
  VN216_in4 <= VN_sign_in(1300) & VN_data_in(1300);
  VN216_in5 <= VN_sign_in(1301) & VN_data_in(1301);
  VN217_in0 <= VN_sign_in(1302) & VN_data_in(1302);
  VN217_in1 <= VN_sign_in(1303) & VN_data_in(1303);
  VN217_in2 <= VN_sign_in(1304) & VN_data_in(1304);
  VN217_in3 <= VN_sign_in(1305) & VN_data_in(1305);
  VN217_in4 <= VN_sign_in(1306) & VN_data_in(1306);
  VN217_in5 <= VN_sign_in(1307) & VN_data_in(1307);
  VN218_in0 <= VN_sign_in(1308) & VN_data_in(1308);
  VN218_in1 <= VN_sign_in(1309) & VN_data_in(1309);
  VN218_in2 <= VN_sign_in(1310) & VN_data_in(1310);
  VN218_in3 <= VN_sign_in(1311) & VN_data_in(1311);
  VN218_in4 <= VN_sign_in(1312) & VN_data_in(1312);
  VN218_in5 <= VN_sign_in(1313) & VN_data_in(1313);
  VN219_in0 <= VN_sign_in(1314) & VN_data_in(1314);
  VN219_in1 <= VN_sign_in(1315) & VN_data_in(1315);
  VN219_in2 <= VN_sign_in(1316) & VN_data_in(1316);
  VN219_in3 <= VN_sign_in(1317) & VN_data_in(1317);
  VN219_in4 <= VN_sign_in(1318) & VN_data_in(1318);
  VN219_in5 <= VN_sign_in(1319) & VN_data_in(1319);
  VN220_in0 <= VN_sign_in(1320) & VN_data_in(1320);
  VN220_in1 <= VN_sign_in(1321) & VN_data_in(1321);
  VN220_in2 <= VN_sign_in(1322) & VN_data_in(1322);
  VN220_in3 <= VN_sign_in(1323) & VN_data_in(1323);
  VN220_in4 <= VN_sign_in(1324) & VN_data_in(1324);
  VN220_in5 <= VN_sign_in(1325) & VN_data_in(1325);
  VN221_in0 <= VN_sign_in(1326) & VN_data_in(1326);
  VN221_in1 <= VN_sign_in(1327) & VN_data_in(1327);
  VN221_in2 <= VN_sign_in(1328) & VN_data_in(1328);
  VN221_in3 <= VN_sign_in(1329) & VN_data_in(1329);
  VN221_in4 <= VN_sign_in(1330) & VN_data_in(1330);
  VN221_in5 <= VN_sign_in(1331) & VN_data_in(1331);
  VN222_in0 <= VN_sign_in(1332) & VN_data_in(1332);
  VN222_in1 <= VN_sign_in(1333) & VN_data_in(1333);
  VN222_in2 <= VN_sign_in(1334) & VN_data_in(1334);
  VN222_in3 <= VN_sign_in(1335) & VN_data_in(1335);
  VN222_in4 <= VN_sign_in(1336) & VN_data_in(1336);
  VN222_in5 <= VN_sign_in(1337) & VN_data_in(1337);
  VN223_in0 <= VN_sign_in(1338) & VN_data_in(1338);
  VN223_in1 <= VN_sign_in(1339) & VN_data_in(1339);
  VN223_in2 <= VN_sign_in(1340) & VN_data_in(1340);
  VN223_in3 <= VN_sign_in(1341) & VN_data_in(1341);
  VN223_in4 <= VN_sign_in(1342) & VN_data_in(1342);
  VN223_in5 <= VN_sign_in(1343) & VN_data_in(1343);
  VN224_in0 <= VN_sign_in(1344) & VN_data_in(1344);
  VN224_in1 <= VN_sign_in(1345) & VN_data_in(1345);
  VN224_in2 <= VN_sign_in(1346) & VN_data_in(1346);
  VN224_in3 <= VN_sign_in(1347) & VN_data_in(1347);
  VN224_in4 <= VN_sign_in(1348) & VN_data_in(1348);
  VN224_in5 <= VN_sign_in(1349) & VN_data_in(1349);
  VN225_in0 <= VN_sign_in(1350) & VN_data_in(1350);
  VN225_in1 <= VN_sign_in(1351) & VN_data_in(1351);
  VN225_in2 <= VN_sign_in(1352) & VN_data_in(1352);
  VN225_in3 <= VN_sign_in(1353) & VN_data_in(1353);
  VN225_in4 <= VN_sign_in(1354) & VN_data_in(1354);
  VN225_in5 <= VN_sign_in(1355) & VN_data_in(1355);
  VN226_in0 <= VN_sign_in(1356) & VN_data_in(1356);
  VN226_in1 <= VN_sign_in(1357) & VN_data_in(1357);
  VN226_in2 <= VN_sign_in(1358) & VN_data_in(1358);
  VN226_in3 <= VN_sign_in(1359) & VN_data_in(1359);
  VN226_in4 <= VN_sign_in(1360) & VN_data_in(1360);
  VN226_in5 <= VN_sign_in(1361) & VN_data_in(1361);
  VN227_in0 <= VN_sign_in(1362) & VN_data_in(1362);
  VN227_in1 <= VN_sign_in(1363) & VN_data_in(1363);
  VN227_in2 <= VN_sign_in(1364) & VN_data_in(1364);
  VN227_in3 <= VN_sign_in(1365) & VN_data_in(1365);
  VN227_in4 <= VN_sign_in(1366) & VN_data_in(1366);
  VN227_in5 <= VN_sign_in(1367) & VN_data_in(1367);
  VN228_in0 <= VN_sign_in(1368) & VN_data_in(1368);
  VN228_in1 <= VN_sign_in(1369) & VN_data_in(1369);
  VN228_in2 <= VN_sign_in(1370) & VN_data_in(1370);
  VN228_in3 <= VN_sign_in(1371) & VN_data_in(1371);
  VN228_in4 <= VN_sign_in(1372) & VN_data_in(1372);
  VN228_in5 <= VN_sign_in(1373) & VN_data_in(1373);
  VN229_in0 <= VN_sign_in(1374) & VN_data_in(1374);
  VN229_in1 <= VN_sign_in(1375) & VN_data_in(1375);
  VN229_in2 <= VN_sign_in(1376) & VN_data_in(1376);
  VN229_in3 <= VN_sign_in(1377) & VN_data_in(1377);
  VN229_in4 <= VN_sign_in(1378) & VN_data_in(1378);
  VN229_in5 <= VN_sign_in(1379) & VN_data_in(1379);
  VN230_in0 <= VN_sign_in(1380) & VN_data_in(1380);
  VN230_in1 <= VN_sign_in(1381) & VN_data_in(1381);
  VN230_in2 <= VN_sign_in(1382) & VN_data_in(1382);
  VN230_in3 <= VN_sign_in(1383) & VN_data_in(1383);
  VN230_in4 <= VN_sign_in(1384) & VN_data_in(1384);
  VN230_in5 <= VN_sign_in(1385) & VN_data_in(1385);
  VN231_in0 <= VN_sign_in(1386) & VN_data_in(1386);
  VN231_in1 <= VN_sign_in(1387) & VN_data_in(1387);
  VN231_in2 <= VN_sign_in(1388) & VN_data_in(1388);
  VN231_in3 <= VN_sign_in(1389) & VN_data_in(1389);
  VN231_in4 <= VN_sign_in(1390) & VN_data_in(1390);
  VN231_in5 <= VN_sign_in(1391) & VN_data_in(1391);
  VN232_in0 <= VN_sign_in(1392) & VN_data_in(1392);
  VN232_in1 <= VN_sign_in(1393) & VN_data_in(1393);
  VN232_in2 <= VN_sign_in(1394) & VN_data_in(1394);
  VN232_in3 <= VN_sign_in(1395) & VN_data_in(1395);
  VN232_in4 <= VN_sign_in(1396) & VN_data_in(1396);
  VN232_in5 <= VN_sign_in(1397) & VN_data_in(1397);
  VN233_in0 <= VN_sign_in(1398) & VN_data_in(1398);
  VN233_in1 <= VN_sign_in(1399) & VN_data_in(1399);
  VN233_in2 <= VN_sign_in(1400) & VN_data_in(1400);
  VN233_in3 <= VN_sign_in(1401) & VN_data_in(1401);
  VN233_in4 <= VN_sign_in(1402) & VN_data_in(1402);
  VN233_in5 <= VN_sign_in(1403) & VN_data_in(1403);
  VN234_in0 <= VN_sign_in(1404) & VN_data_in(1404);
  VN234_in1 <= VN_sign_in(1405) & VN_data_in(1405);
  VN234_in2 <= VN_sign_in(1406) & VN_data_in(1406);
  VN234_in3 <= VN_sign_in(1407) & VN_data_in(1407);
  VN234_in4 <= VN_sign_in(1408) & VN_data_in(1408);
  VN234_in5 <= VN_sign_in(1409) & VN_data_in(1409);
  VN235_in0 <= VN_sign_in(1410) & VN_data_in(1410);
  VN235_in1 <= VN_sign_in(1411) & VN_data_in(1411);
  VN235_in2 <= VN_sign_in(1412) & VN_data_in(1412);
  VN235_in3 <= VN_sign_in(1413) & VN_data_in(1413);
  VN235_in4 <= VN_sign_in(1414) & VN_data_in(1414);
  VN235_in5 <= VN_sign_in(1415) & VN_data_in(1415);
  VN236_in0 <= VN_sign_in(1416) & VN_data_in(1416);
  VN236_in1 <= VN_sign_in(1417) & VN_data_in(1417);
  VN236_in2 <= VN_sign_in(1418) & VN_data_in(1418);
  VN236_in3 <= VN_sign_in(1419) & VN_data_in(1419);
  VN236_in4 <= VN_sign_in(1420) & VN_data_in(1420);
  VN236_in5 <= VN_sign_in(1421) & VN_data_in(1421);
  VN237_in0 <= VN_sign_in(1422) & VN_data_in(1422);
  VN237_in1 <= VN_sign_in(1423) & VN_data_in(1423);
  VN237_in2 <= VN_sign_in(1424) & VN_data_in(1424);
  VN237_in3 <= VN_sign_in(1425) & VN_data_in(1425);
  VN237_in4 <= VN_sign_in(1426) & VN_data_in(1426);
  VN237_in5 <= VN_sign_in(1427) & VN_data_in(1427);
  VN238_in0 <= VN_sign_in(1428) & VN_data_in(1428);
  VN238_in1 <= VN_sign_in(1429) & VN_data_in(1429);
  VN238_in2 <= VN_sign_in(1430) & VN_data_in(1430);
  VN238_in3 <= VN_sign_in(1431) & VN_data_in(1431);
  VN238_in4 <= VN_sign_in(1432) & VN_data_in(1432);
  VN238_in5 <= VN_sign_in(1433) & VN_data_in(1433);
  VN239_in0 <= VN_sign_in(1434) & VN_data_in(1434);
  VN239_in1 <= VN_sign_in(1435) & VN_data_in(1435);
  VN239_in2 <= VN_sign_in(1436) & VN_data_in(1436);
  VN239_in3 <= VN_sign_in(1437) & VN_data_in(1437);
  VN239_in4 <= VN_sign_in(1438) & VN_data_in(1438);
  VN239_in5 <= VN_sign_in(1439) & VN_data_in(1439);
  VN240_in0 <= VN_sign_in(1440) & VN_data_in(1440);
  VN240_in1 <= VN_sign_in(1441) & VN_data_in(1441);
  VN240_in2 <= VN_sign_in(1442) & VN_data_in(1442);
  VN240_in3 <= VN_sign_in(1443) & VN_data_in(1443);
  VN240_in4 <= VN_sign_in(1444) & VN_data_in(1444);
  VN240_in5 <= VN_sign_in(1445) & VN_data_in(1445);
  VN241_in0 <= VN_sign_in(1446) & VN_data_in(1446);
  VN241_in1 <= VN_sign_in(1447) & VN_data_in(1447);
  VN241_in2 <= VN_sign_in(1448) & VN_data_in(1448);
  VN241_in3 <= VN_sign_in(1449) & VN_data_in(1449);
  VN241_in4 <= VN_sign_in(1450) & VN_data_in(1450);
  VN241_in5 <= VN_sign_in(1451) & VN_data_in(1451);
  VN242_in0 <= VN_sign_in(1452) & VN_data_in(1452);
  VN242_in1 <= VN_sign_in(1453) & VN_data_in(1453);
  VN242_in2 <= VN_sign_in(1454) & VN_data_in(1454);
  VN242_in3 <= VN_sign_in(1455) & VN_data_in(1455);
  VN242_in4 <= VN_sign_in(1456) & VN_data_in(1456);
  VN242_in5 <= VN_sign_in(1457) & VN_data_in(1457);
  VN243_in0 <= VN_sign_in(1458) & VN_data_in(1458);
  VN243_in1 <= VN_sign_in(1459) & VN_data_in(1459);
  VN243_in2 <= VN_sign_in(1460) & VN_data_in(1460);
  VN243_in3 <= VN_sign_in(1461) & VN_data_in(1461);
  VN243_in4 <= VN_sign_in(1462) & VN_data_in(1462);
  VN243_in5 <= VN_sign_in(1463) & VN_data_in(1463);
  VN244_in0 <= VN_sign_in(1464) & VN_data_in(1464);
  VN244_in1 <= VN_sign_in(1465) & VN_data_in(1465);
  VN244_in2 <= VN_sign_in(1466) & VN_data_in(1466);
  VN244_in3 <= VN_sign_in(1467) & VN_data_in(1467);
  VN244_in4 <= VN_sign_in(1468) & VN_data_in(1468);
  VN244_in5 <= VN_sign_in(1469) & VN_data_in(1469);
  VN245_in0 <= VN_sign_in(1470) & VN_data_in(1470);
  VN245_in1 <= VN_sign_in(1471) & VN_data_in(1471);
  VN245_in2 <= VN_sign_in(1472) & VN_data_in(1472);
  VN245_in3 <= VN_sign_in(1473) & VN_data_in(1473);
  VN245_in4 <= VN_sign_in(1474) & VN_data_in(1474);
  VN245_in5 <= VN_sign_in(1475) & VN_data_in(1475);
  VN246_in0 <= VN_sign_in(1476) & VN_data_in(1476);
  VN246_in1 <= VN_sign_in(1477) & VN_data_in(1477);
  VN246_in2 <= VN_sign_in(1478) & VN_data_in(1478);
  VN246_in3 <= VN_sign_in(1479) & VN_data_in(1479);
  VN246_in4 <= VN_sign_in(1480) & VN_data_in(1480);
  VN246_in5 <= VN_sign_in(1481) & VN_data_in(1481);
  VN247_in0 <= VN_sign_in(1482) & VN_data_in(1482);
  VN247_in1 <= VN_sign_in(1483) & VN_data_in(1483);
  VN247_in2 <= VN_sign_in(1484) & VN_data_in(1484);
  VN247_in3 <= VN_sign_in(1485) & VN_data_in(1485);
  VN247_in4 <= VN_sign_in(1486) & VN_data_in(1486);
  VN247_in5 <= VN_sign_in(1487) & VN_data_in(1487);
  VN248_in0 <= VN_sign_in(1488) & VN_data_in(1488);
  VN248_in1 <= VN_sign_in(1489) & VN_data_in(1489);
  VN248_in2 <= VN_sign_in(1490) & VN_data_in(1490);
  VN248_in3 <= VN_sign_in(1491) & VN_data_in(1491);
  VN248_in4 <= VN_sign_in(1492) & VN_data_in(1492);
  VN248_in5 <= VN_sign_in(1493) & VN_data_in(1493);
  VN249_in0 <= VN_sign_in(1494) & VN_data_in(1494);
  VN249_in1 <= VN_sign_in(1495) & VN_data_in(1495);
  VN249_in2 <= VN_sign_in(1496) & VN_data_in(1496);
  VN249_in3 <= VN_sign_in(1497) & VN_data_in(1497);
  VN249_in4 <= VN_sign_in(1498) & VN_data_in(1498);
  VN249_in5 <= VN_sign_in(1499) & VN_data_in(1499);
  VN250_in0 <= VN_sign_in(1500) & VN_data_in(1500);
  VN250_in1 <= VN_sign_in(1501) & VN_data_in(1501);
  VN250_in2 <= VN_sign_in(1502) & VN_data_in(1502);
  VN250_in3 <= VN_sign_in(1503) & VN_data_in(1503);
  VN250_in4 <= VN_sign_in(1504) & VN_data_in(1504);
  VN250_in5 <= VN_sign_in(1505) & VN_data_in(1505);
  VN251_in0 <= VN_sign_in(1506) & VN_data_in(1506);
  VN251_in1 <= VN_sign_in(1507) & VN_data_in(1507);
  VN251_in2 <= VN_sign_in(1508) & VN_data_in(1508);
  VN251_in3 <= VN_sign_in(1509) & VN_data_in(1509);
  VN251_in4 <= VN_sign_in(1510) & VN_data_in(1510);
  VN251_in5 <= VN_sign_in(1511) & VN_data_in(1511);
  VN252_in0 <= VN_sign_in(1512) & VN_data_in(1512);
  VN252_in1 <= VN_sign_in(1513) & VN_data_in(1513);
  VN252_in2 <= VN_sign_in(1514) & VN_data_in(1514);
  VN252_in3 <= VN_sign_in(1515) & VN_data_in(1515);
  VN252_in4 <= VN_sign_in(1516) & VN_data_in(1516);
  VN252_in5 <= VN_sign_in(1517) & VN_data_in(1517);
  VN253_in0 <= VN_sign_in(1518) & VN_data_in(1518);
  VN253_in1 <= VN_sign_in(1519) & VN_data_in(1519);
  VN253_in2 <= VN_sign_in(1520) & VN_data_in(1520);
  VN253_in3 <= VN_sign_in(1521) & VN_data_in(1521);
  VN253_in4 <= VN_sign_in(1522) & VN_data_in(1522);
  VN253_in5 <= VN_sign_in(1523) & VN_data_in(1523);
  VN254_in0 <= VN_sign_in(1524) & VN_data_in(1524);
  VN254_in1 <= VN_sign_in(1525) & VN_data_in(1525);
  VN254_in2 <= VN_sign_in(1526) & VN_data_in(1526);
  VN254_in3 <= VN_sign_in(1527) & VN_data_in(1527);
  VN254_in4 <= VN_sign_in(1528) & VN_data_in(1528);
  VN254_in5 <= VN_sign_in(1529) & VN_data_in(1529);
  VN255_in0 <= VN_sign_in(1530) & VN_data_in(1530);
  VN255_in1 <= VN_sign_in(1531) & VN_data_in(1531);
  VN255_in2 <= VN_sign_in(1532) & VN_data_in(1532);
  VN255_in3 <= VN_sign_in(1533) & VN_data_in(1533);
  VN255_in4 <= VN_sign_in(1534) & VN_data_in(1534);
  VN255_in5 <= VN_sign_in(1535) & VN_data_in(1535);
  VN256_in0 <= VN_sign_in(1536) & VN_data_in(1536);
  VN256_in1 <= VN_sign_in(1537) & VN_data_in(1537);
  VN256_in2 <= VN_sign_in(1538) & VN_data_in(1538);
  VN256_in3 <= VN_sign_in(1539) & VN_data_in(1539);
  VN256_in4 <= VN_sign_in(1540) & VN_data_in(1540);
  VN256_in5 <= VN_sign_in(1541) & VN_data_in(1541);
  VN257_in0 <= VN_sign_in(1542) & VN_data_in(1542);
  VN257_in1 <= VN_sign_in(1543) & VN_data_in(1543);
  VN257_in2 <= VN_sign_in(1544) & VN_data_in(1544);
  VN257_in3 <= VN_sign_in(1545) & VN_data_in(1545);
  VN257_in4 <= VN_sign_in(1546) & VN_data_in(1546);
  VN257_in5 <= VN_sign_in(1547) & VN_data_in(1547);
  VN258_in0 <= VN_sign_in(1548) & VN_data_in(1548);
  VN258_in1 <= VN_sign_in(1549) & VN_data_in(1549);
  VN258_in2 <= VN_sign_in(1550) & VN_data_in(1550);
  VN258_in3 <= VN_sign_in(1551) & VN_data_in(1551);
  VN258_in4 <= VN_sign_in(1552) & VN_data_in(1552);
  VN258_in5 <= VN_sign_in(1553) & VN_data_in(1553);
  VN259_in0 <= VN_sign_in(1554) & VN_data_in(1554);
  VN259_in1 <= VN_sign_in(1555) & VN_data_in(1555);
  VN259_in2 <= VN_sign_in(1556) & VN_data_in(1556);
  VN259_in3 <= VN_sign_in(1557) & VN_data_in(1557);
  VN259_in4 <= VN_sign_in(1558) & VN_data_in(1558);
  VN259_in5 <= VN_sign_in(1559) & VN_data_in(1559);
  VN260_in0 <= VN_sign_in(1560) & VN_data_in(1560);
  VN260_in1 <= VN_sign_in(1561) & VN_data_in(1561);
  VN260_in2 <= VN_sign_in(1562) & VN_data_in(1562);
  VN260_in3 <= VN_sign_in(1563) & VN_data_in(1563);
  VN260_in4 <= VN_sign_in(1564) & VN_data_in(1564);
  VN260_in5 <= VN_sign_in(1565) & VN_data_in(1565);
  VN261_in0 <= VN_sign_in(1566) & VN_data_in(1566);
  VN261_in1 <= VN_sign_in(1567) & VN_data_in(1567);
  VN261_in2 <= VN_sign_in(1568) & VN_data_in(1568);
  VN261_in3 <= VN_sign_in(1569) & VN_data_in(1569);
  VN261_in4 <= VN_sign_in(1570) & VN_data_in(1570);
  VN261_in5 <= VN_sign_in(1571) & VN_data_in(1571);
  VN262_in0 <= VN_sign_in(1572) & VN_data_in(1572);
  VN262_in1 <= VN_sign_in(1573) & VN_data_in(1573);
  VN262_in2 <= VN_sign_in(1574) & VN_data_in(1574);
  VN262_in3 <= VN_sign_in(1575) & VN_data_in(1575);
  VN262_in4 <= VN_sign_in(1576) & VN_data_in(1576);
  VN262_in5 <= VN_sign_in(1577) & VN_data_in(1577);
  VN263_in0 <= VN_sign_in(1578) & VN_data_in(1578);
  VN263_in1 <= VN_sign_in(1579) & VN_data_in(1579);
  VN263_in2 <= VN_sign_in(1580) & VN_data_in(1580);
  VN263_in3 <= VN_sign_in(1581) & VN_data_in(1581);
  VN263_in4 <= VN_sign_in(1582) & VN_data_in(1582);
  VN263_in5 <= VN_sign_in(1583) & VN_data_in(1583);
  VN264_in0 <= VN_sign_in(1584) & VN_data_in(1584);
  VN264_in1 <= VN_sign_in(1585) & VN_data_in(1585);
  VN264_in2 <= VN_sign_in(1586) & VN_data_in(1586);
  VN264_in3 <= VN_sign_in(1587) & VN_data_in(1587);
  VN264_in4 <= VN_sign_in(1588) & VN_data_in(1588);
  VN264_in5 <= VN_sign_in(1589) & VN_data_in(1589);
  VN265_in0 <= VN_sign_in(1590) & VN_data_in(1590);
  VN265_in1 <= VN_sign_in(1591) & VN_data_in(1591);
  VN265_in2 <= VN_sign_in(1592) & VN_data_in(1592);
  VN265_in3 <= VN_sign_in(1593) & VN_data_in(1593);
  VN265_in4 <= VN_sign_in(1594) & VN_data_in(1594);
  VN265_in5 <= VN_sign_in(1595) & VN_data_in(1595);
  VN266_in0 <= VN_sign_in(1596) & VN_data_in(1596);
  VN266_in1 <= VN_sign_in(1597) & VN_data_in(1597);
  VN266_in2 <= VN_sign_in(1598) & VN_data_in(1598);
  VN266_in3 <= VN_sign_in(1599) & VN_data_in(1599);
  VN266_in4 <= VN_sign_in(1600) & VN_data_in(1600);
  VN266_in5 <= VN_sign_in(1601) & VN_data_in(1601);
  VN267_in0 <= VN_sign_in(1602) & VN_data_in(1602);
  VN267_in1 <= VN_sign_in(1603) & VN_data_in(1603);
  VN267_in2 <= VN_sign_in(1604) & VN_data_in(1604);
  VN267_in3 <= VN_sign_in(1605) & VN_data_in(1605);
  VN267_in4 <= VN_sign_in(1606) & VN_data_in(1606);
  VN267_in5 <= VN_sign_in(1607) & VN_data_in(1607);
  VN268_in0 <= VN_sign_in(1608) & VN_data_in(1608);
  VN268_in1 <= VN_sign_in(1609) & VN_data_in(1609);
  VN268_in2 <= VN_sign_in(1610) & VN_data_in(1610);
  VN268_in3 <= VN_sign_in(1611) & VN_data_in(1611);
  VN268_in4 <= VN_sign_in(1612) & VN_data_in(1612);
  VN268_in5 <= VN_sign_in(1613) & VN_data_in(1613);
  VN269_in0 <= VN_sign_in(1614) & VN_data_in(1614);
  VN269_in1 <= VN_sign_in(1615) & VN_data_in(1615);
  VN269_in2 <= VN_sign_in(1616) & VN_data_in(1616);
  VN269_in3 <= VN_sign_in(1617) & VN_data_in(1617);
  VN269_in4 <= VN_sign_in(1618) & VN_data_in(1618);
  VN269_in5 <= VN_sign_in(1619) & VN_data_in(1619);
  VN270_in0 <= VN_sign_in(1620) & VN_data_in(1620);
  VN270_in1 <= VN_sign_in(1621) & VN_data_in(1621);
  VN270_in2 <= VN_sign_in(1622) & VN_data_in(1622);
  VN270_in3 <= VN_sign_in(1623) & VN_data_in(1623);
  VN270_in4 <= VN_sign_in(1624) & VN_data_in(1624);
  VN270_in5 <= VN_sign_in(1625) & VN_data_in(1625);
  VN271_in0 <= VN_sign_in(1626) & VN_data_in(1626);
  VN271_in1 <= VN_sign_in(1627) & VN_data_in(1627);
  VN271_in2 <= VN_sign_in(1628) & VN_data_in(1628);
  VN271_in3 <= VN_sign_in(1629) & VN_data_in(1629);
  VN271_in4 <= VN_sign_in(1630) & VN_data_in(1630);
  VN271_in5 <= VN_sign_in(1631) & VN_data_in(1631);
  VN272_in0 <= VN_sign_in(1632) & VN_data_in(1632);
  VN272_in1 <= VN_sign_in(1633) & VN_data_in(1633);
  VN272_in2 <= VN_sign_in(1634) & VN_data_in(1634);
  VN272_in3 <= VN_sign_in(1635) & VN_data_in(1635);
  VN272_in4 <= VN_sign_in(1636) & VN_data_in(1636);
  VN272_in5 <= VN_sign_in(1637) & VN_data_in(1637);
  VN273_in0 <= VN_sign_in(1638) & VN_data_in(1638);
  VN273_in1 <= VN_sign_in(1639) & VN_data_in(1639);
  VN273_in2 <= VN_sign_in(1640) & VN_data_in(1640);
  VN273_in3 <= VN_sign_in(1641) & VN_data_in(1641);
  VN273_in4 <= VN_sign_in(1642) & VN_data_in(1642);
  VN273_in5 <= VN_sign_in(1643) & VN_data_in(1643);
  VN274_in0 <= VN_sign_in(1644) & VN_data_in(1644);
  VN274_in1 <= VN_sign_in(1645) & VN_data_in(1645);
  VN274_in2 <= VN_sign_in(1646) & VN_data_in(1646);
  VN274_in3 <= VN_sign_in(1647) & VN_data_in(1647);
  VN274_in4 <= VN_sign_in(1648) & VN_data_in(1648);
  VN274_in5 <= VN_sign_in(1649) & VN_data_in(1649);
  VN275_in0 <= VN_sign_in(1650) & VN_data_in(1650);
  VN275_in1 <= VN_sign_in(1651) & VN_data_in(1651);
  VN275_in2 <= VN_sign_in(1652) & VN_data_in(1652);
  VN275_in3 <= VN_sign_in(1653) & VN_data_in(1653);
  VN275_in4 <= VN_sign_in(1654) & VN_data_in(1654);
  VN275_in5 <= VN_sign_in(1655) & VN_data_in(1655);
  VN276_in0 <= VN_sign_in(1656) & VN_data_in(1656);
  VN276_in1 <= VN_sign_in(1657) & VN_data_in(1657);
  VN276_in2 <= VN_sign_in(1658) & VN_data_in(1658);
  VN276_in3 <= VN_sign_in(1659) & VN_data_in(1659);
  VN276_in4 <= VN_sign_in(1660) & VN_data_in(1660);
  VN276_in5 <= VN_sign_in(1661) & VN_data_in(1661);
  VN277_in0 <= VN_sign_in(1662) & VN_data_in(1662);
  VN277_in1 <= VN_sign_in(1663) & VN_data_in(1663);
  VN277_in2 <= VN_sign_in(1664) & VN_data_in(1664);
  VN277_in3 <= VN_sign_in(1665) & VN_data_in(1665);
  VN277_in4 <= VN_sign_in(1666) & VN_data_in(1666);
  VN277_in5 <= VN_sign_in(1667) & VN_data_in(1667);
  VN278_in0 <= VN_sign_in(1668) & VN_data_in(1668);
  VN278_in1 <= VN_sign_in(1669) & VN_data_in(1669);
  VN278_in2 <= VN_sign_in(1670) & VN_data_in(1670);
  VN278_in3 <= VN_sign_in(1671) & VN_data_in(1671);
  VN278_in4 <= VN_sign_in(1672) & VN_data_in(1672);
  VN278_in5 <= VN_sign_in(1673) & VN_data_in(1673);
  VN279_in0 <= VN_sign_in(1674) & VN_data_in(1674);
  VN279_in1 <= VN_sign_in(1675) & VN_data_in(1675);
  VN279_in2 <= VN_sign_in(1676) & VN_data_in(1676);
  VN279_in3 <= VN_sign_in(1677) & VN_data_in(1677);
  VN279_in4 <= VN_sign_in(1678) & VN_data_in(1678);
  VN279_in5 <= VN_sign_in(1679) & VN_data_in(1679);
  VN280_in0 <= VN_sign_in(1680) & VN_data_in(1680);
  VN280_in1 <= VN_sign_in(1681) & VN_data_in(1681);
  VN280_in2 <= VN_sign_in(1682) & VN_data_in(1682);
  VN280_in3 <= VN_sign_in(1683) & VN_data_in(1683);
  VN280_in4 <= VN_sign_in(1684) & VN_data_in(1684);
  VN280_in5 <= VN_sign_in(1685) & VN_data_in(1685);
  VN281_in0 <= VN_sign_in(1686) & VN_data_in(1686);
  VN281_in1 <= VN_sign_in(1687) & VN_data_in(1687);
  VN281_in2 <= VN_sign_in(1688) & VN_data_in(1688);
  VN281_in3 <= VN_sign_in(1689) & VN_data_in(1689);
  VN281_in4 <= VN_sign_in(1690) & VN_data_in(1690);
  VN281_in5 <= VN_sign_in(1691) & VN_data_in(1691);
  VN282_in0 <= VN_sign_in(1692) & VN_data_in(1692);
  VN282_in1 <= VN_sign_in(1693) & VN_data_in(1693);
  VN282_in2 <= VN_sign_in(1694) & VN_data_in(1694);
  VN282_in3 <= VN_sign_in(1695) & VN_data_in(1695);
  VN282_in4 <= VN_sign_in(1696) & VN_data_in(1696);
  VN282_in5 <= VN_sign_in(1697) & VN_data_in(1697);
  VN283_in0 <= VN_sign_in(1698) & VN_data_in(1698);
  VN283_in1 <= VN_sign_in(1699) & VN_data_in(1699);
  VN283_in2 <= VN_sign_in(1700) & VN_data_in(1700);
  VN283_in3 <= VN_sign_in(1701) & VN_data_in(1701);
  VN283_in4 <= VN_sign_in(1702) & VN_data_in(1702);
  VN283_in5 <= VN_sign_in(1703) & VN_data_in(1703);
  VN284_in0 <= VN_sign_in(1704) & VN_data_in(1704);
  VN284_in1 <= VN_sign_in(1705) & VN_data_in(1705);
  VN284_in2 <= VN_sign_in(1706) & VN_data_in(1706);
  VN284_in3 <= VN_sign_in(1707) & VN_data_in(1707);
  VN284_in4 <= VN_sign_in(1708) & VN_data_in(1708);
  VN284_in5 <= VN_sign_in(1709) & VN_data_in(1709);
  VN285_in0 <= VN_sign_in(1710) & VN_data_in(1710);
  VN285_in1 <= VN_sign_in(1711) & VN_data_in(1711);
  VN285_in2 <= VN_sign_in(1712) & VN_data_in(1712);
  VN285_in3 <= VN_sign_in(1713) & VN_data_in(1713);
  VN285_in4 <= VN_sign_in(1714) & VN_data_in(1714);
  VN285_in5 <= VN_sign_in(1715) & VN_data_in(1715);
  VN286_in0 <= VN_sign_in(1716) & VN_data_in(1716);
  VN286_in1 <= VN_sign_in(1717) & VN_data_in(1717);
  VN286_in2 <= VN_sign_in(1718) & VN_data_in(1718);
  VN286_in3 <= VN_sign_in(1719) & VN_data_in(1719);
  VN286_in4 <= VN_sign_in(1720) & VN_data_in(1720);
  VN286_in5 <= VN_sign_in(1721) & VN_data_in(1721);
  VN287_in0 <= VN_sign_in(1722) & VN_data_in(1722);
  VN287_in1 <= VN_sign_in(1723) & VN_data_in(1723);
  VN287_in2 <= VN_sign_in(1724) & VN_data_in(1724);
  VN287_in3 <= VN_sign_in(1725) & VN_data_in(1725);
  VN287_in4 <= VN_sign_in(1726) & VN_data_in(1726);
  VN287_in5 <= VN_sign_in(1727) & VN_data_in(1727);
  VN288_in0 <= VN_sign_in(1728) & VN_data_in(1728);
  VN288_in1 <= VN_sign_in(1729) & VN_data_in(1729);
  VN288_in2 <= VN_sign_in(1730) & VN_data_in(1730);
  VN288_in3 <= VN_sign_in(1731) & VN_data_in(1731);
  VN288_in4 <= VN_sign_in(1732) & VN_data_in(1732);
  VN288_in5 <= VN_sign_in(1733) & VN_data_in(1733);
  VN289_in0 <= VN_sign_in(1734) & VN_data_in(1734);
  VN289_in1 <= VN_sign_in(1735) & VN_data_in(1735);
  VN289_in2 <= VN_sign_in(1736) & VN_data_in(1736);
  VN289_in3 <= VN_sign_in(1737) & VN_data_in(1737);
  VN289_in4 <= VN_sign_in(1738) & VN_data_in(1738);
  VN289_in5 <= VN_sign_in(1739) & VN_data_in(1739);
  VN290_in0 <= VN_sign_in(1740) & VN_data_in(1740);
  VN290_in1 <= VN_sign_in(1741) & VN_data_in(1741);
  VN290_in2 <= VN_sign_in(1742) & VN_data_in(1742);
  VN290_in3 <= VN_sign_in(1743) & VN_data_in(1743);
  VN290_in4 <= VN_sign_in(1744) & VN_data_in(1744);
  VN290_in5 <= VN_sign_in(1745) & VN_data_in(1745);
  VN291_in0 <= VN_sign_in(1746) & VN_data_in(1746);
  VN291_in1 <= VN_sign_in(1747) & VN_data_in(1747);
  VN291_in2 <= VN_sign_in(1748) & VN_data_in(1748);
  VN291_in3 <= VN_sign_in(1749) & VN_data_in(1749);
  VN291_in4 <= VN_sign_in(1750) & VN_data_in(1750);
  VN291_in5 <= VN_sign_in(1751) & VN_data_in(1751);
  VN292_in0 <= VN_sign_in(1752) & VN_data_in(1752);
  VN292_in1 <= VN_sign_in(1753) & VN_data_in(1753);
  VN292_in2 <= VN_sign_in(1754) & VN_data_in(1754);
  VN292_in3 <= VN_sign_in(1755) & VN_data_in(1755);
  VN292_in4 <= VN_sign_in(1756) & VN_data_in(1756);
  VN292_in5 <= VN_sign_in(1757) & VN_data_in(1757);
  VN293_in0 <= VN_sign_in(1758) & VN_data_in(1758);
  VN293_in1 <= VN_sign_in(1759) & VN_data_in(1759);
  VN293_in2 <= VN_sign_in(1760) & VN_data_in(1760);
  VN293_in3 <= VN_sign_in(1761) & VN_data_in(1761);
  VN293_in4 <= VN_sign_in(1762) & VN_data_in(1762);
  VN293_in5 <= VN_sign_in(1763) & VN_data_in(1763);
  VN294_in0 <= VN_sign_in(1764) & VN_data_in(1764);
  VN294_in1 <= VN_sign_in(1765) & VN_data_in(1765);
  VN294_in2 <= VN_sign_in(1766) & VN_data_in(1766);
  VN294_in3 <= VN_sign_in(1767) & VN_data_in(1767);
  VN294_in4 <= VN_sign_in(1768) & VN_data_in(1768);
  VN294_in5 <= VN_sign_in(1769) & VN_data_in(1769);
  VN295_in0 <= VN_sign_in(1770) & VN_data_in(1770);
  VN295_in1 <= VN_sign_in(1771) & VN_data_in(1771);
  VN295_in2 <= VN_sign_in(1772) & VN_data_in(1772);
  VN295_in3 <= VN_sign_in(1773) & VN_data_in(1773);
  VN295_in4 <= VN_sign_in(1774) & VN_data_in(1774);
  VN295_in5 <= VN_sign_in(1775) & VN_data_in(1775);
  VN296_in0 <= VN_sign_in(1776) & VN_data_in(1776);
  VN296_in1 <= VN_sign_in(1777) & VN_data_in(1777);
  VN296_in2 <= VN_sign_in(1778) & VN_data_in(1778);
  VN296_in3 <= VN_sign_in(1779) & VN_data_in(1779);
  VN296_in4 <= VN_sign_in(1780) & VN_data_in(1780);
  VN296_in5 <= VN_sign_in(1781) & VN_data_in(1781);
  VN297_in0 <= VN_sign_in(1782) & VN_data_in(1782);
  VN297_in1 <= VN_sign_in(1783) & VN_data_in(1783);
  VN297_in2 <= VN_sign_in(1784) & VN_data_in(1784);
  VN297_in3 <= VN_sign_in(1785) & VN_data_in(1785);
  VN297_in4 <= VN_sign_in(1786) & VN_data_in(1786);
  VN297_in5 <= VN_sign_in(1787) & VN_data_in(1787);
  VN298_in0 <= VN_sign_in(1788) & VN_data_in(1788);
  VN298_in1 <= VN_sign_in(1789) & VN_data_in(1789);
  VN298_in2 <= VN_sign_in(1790) & VN_data_in(1790);
  VN298_in3 <= VN_sign_in(1791) & VN_data_in(1791);
  VN298_in4 <= VN_sign_in(1792) & VN_data_in(1792);
  VN298_in5 <= VN_sign_in(1793) & VN_data_in(1793);
  VN299_in0 <= VN_sign_in(1794) & VN_data_in(1794);
  VN299_in1 <= VN_sign_in(1795) & VN_data_in(1795);
  VN299_in2 <= VN_sign_in(1796) & VN_data_in(1796);
  VN299_in3 <= VN_sign_in(1797) & VN_data_in(1797);
  VN299_in4 <= VN_sign_in(1798) & VN_data_in(1798);
  VN299_in5 <= VN_sign_in(1799) & VN_data_in(1799);
  VN300_in0 <= VN_sign_in(1800) & VN_data_in(1800);
  VN300_in1 <= VN_sign_in(1801) & VN_data_in(1801);
  VN300_in2 <= VN_sign_in(1802) & VN_data_in(1802);
  VN300_in3 <= VN_sign_in(1803) & VN_data_in(1803);
  VN300_in4 <= VN_sign_in(1804) & VN_data_in(1804);
  VN300_in5 <= VN_sign_in(1805) & VN_data_in(1805);
  VN301_in0 <= VN_sign_in(1806) & VN_data_in(1806);
  VN301_in1 <= VN_sign_in(1807) & VN_data_in(1807);
  VN301_in2 <= VN_sign_in(1808) & VN_data_in(1808);
  VN301_in3 <= VN_sign_in(1809) & VN_data_in(1809);
  VN301_in4 <= VN_sign_in(1810) & VN_data_in(1810);
  VN301_in5 <= VN_sign_in(1811) & VN_data_in(1811);
  VN302_in0 <= VN_sign_in(1812) & VN_data_in(1812);
  VN302_in1 <= VN_sign_in(1813) & VN_data_in(1813);
  VN302_in2 <= VN_sign_in(1814) & VN_data_in(1814);
  VN302_in3 <= VN_sign_in(1815) & VN_data_in(1815);
  VN302_in4 <= VN_sign_in(1816) & VN_data_in(1816);
  VN302_in5 <= VN_sign_in(1817) & VN_data_in(1817);
  VN303_in0 <= VN_sign_in(1818) & VN_data_in(1818);
  VN303_in1 <= VN_sign_in(1819) & VN_data_in(1819);
  VN303_in2 <= VN_sign_in(1820) & VN_data_in(1820);
  VN303_in3 <= VN_sign_in(1821) & VN_data_in(1821);
  VN303_in4 <= VN_sign_in(1822) & VN_data_in(1822);
  VN303_in5 <= VN_sign_in(1823) & VN_data_in(1823);
  VN304_in0 <= VN_sign_in(1824) & VN_data_in(1824);
  VN304_in1 <= VN_sign_in(1825) & VN_data_in(1825);
  VN304_in2 <= VN_sign_in(1826) & VN_data_in(1826);
  VN304_in3 <= VN_sign_in(1827) & VN_data_in(1827);
  VN304_in4 <= VN_sign_in(1828) & VN_data_in(1828);
  VN304_in5 <= VN_sign_in(1829) & VN_data_in(1829);
  VN305_in0 <= VN_sign_in(1830) & VN_data_in(1830);
  VN305_in1 <= VN_sign_in(1831) & VN_data_in(1831);
  VN305_in2 <= VN_sign_in(1832) & VN_data_in(1832);
  VN305_in3 <= VN_sign_in(1833) & VN_data_in(1833);
  VN305_in4 <= VN_sign_in(1834) & VN_data_in(1834);
  VN305_in5 <= VN_sign_in(1835) & VN_data_in(1835);
  VN306_in0 <= VN_sign_in(1836) & VN_data_in(1836);
  VN306_in1 <= VN_sign_in(1837) & VN_data_in(1837);
  VN306_in2 <= VN_sign_in(1838) & VN_data_in(1838);
  VN306_in3 <= VN_sign_in(1839) & VN_data_in(1839);
  VN306_in4 <= VN_sign_in(1840) & VN_data_in(1840);
  VN306_in5 <= VN_sign_in(1841) & VN_data_in(1841);
  VN307_in0 <= VN_sign_in(1842) & VN_data_in(1842);
  VN307_in1 <= VN_sign_in(1843) & VN_data_in(1843);
  VN307_in2 <= VN_sign_in(1844) & VN_data_in(1844);
  VN307_in3 <= VN_sign_in(1845) & VN_data_in(1845);
  VN307_in4 <= VN_sign_in(1846) & VN_data_in(1846);
  VN307_in5 <= VN_sign_in(1847) & VN_data_in(1847);
  VN308_in0 <= VN_sign_in(1848) & VN_data_in(1848);
  VN308_in1 <= VN_sign_in(1849) & VN_data_in(1849);
  VN308_in2 <= VN_sign_in(1850) & VN_data_in(1850);
  VN308_in3 <= VN_sign_in(1851) & VN_data_in(1851);
  VN308_in4 <= VN_sign_in(1852) & VN_data_in(1852);
  VN308_in5 <= VN_sign_in(1853) & VN_data_in(1853);
  VN309_in0 <= VN_sign_in(1854) & VN_data_in(1854);
  VN309_in1 <= VN_sign_in(1855) & VN_data_in(1855);
  VN309_in2 <= VN_sign_in(1856) & VN_data_in(1856);
  VN309_in3 <= VN_sign_in(1857) & VN_data_in(1857);
  VN309_in4 <= VN_sign_in(1858) & VN_data_in(1858);
  VN309_in5 <= VN_sign_in(1859) & VN_data_in(1859);
  VN310_in0 <= VN_sign_in(1860) & VN_data_in(1860);
  VN310_in1 <= VN_sign_in(1861) & VN_data_in(1861);
  VN310_in2 <= VN_sign_in(1862) & VN_data_in(1862);
  VN310_in3 <= VN_sign_in(1863) & VN_data_in(1863);
  VN310_in4 <= VN_sign_in(1864) & VN_data_in(1864);
  VN310_in5 <= VN_sign_in(1865) & VN_data_in(1865);
  VN311_in0 <= VN_sign_in(1866) & VN_data_in(1866);
  VN311_in1 <= VN_sign_in(1867) & VN_data_in(1867);
  VN311_in2 <= VN_sign_in(1868) & VN_data_in(1868);
  VN311_in3 <= VN_sign_in(1869) & VN_data_in(1869);
  VN311_in4 <= VN_sign_in(1870) & VN_data_in(1870);
  VN311_in5 <= VN_sign_in(1871) & VN_data_in(1871);
  VN312_in0 <= VN_sign_in(1872) & VN_data_in(1872);
  VN312_in1 <= VN_sign_in(1873) & VN_data_in(1873);
  VN312_in2 <= VN_sign_in(1874) & VN_data_in(1874);
  VN312_in3 <= VN_sign_in(1875) & VN_data_in(1875);
  VN312_in4 <= VN_sign_in(1876) & VN_data_in(1876);
  VN312_in5 <= VN_sign_in(1877) & VN_data_in(1877);
  VN313_in0 <= VN_sign_in(1878) & VN_data_in(1878);
  VN313_in1 <= VN_sign_in(1879) & VN_data_in(1879);
  VN313_in2 <= VN_sign_in(1880) & VN_data_in(1880);
  VN313_in3 <= VN_sign_in(1881) & VN_data_in(1881);
  VN313_in4 <= VN_sign_in(1882) & VN_data_in(1882);
  VN313_in5 <= VN_sign_in(1883) & VN_data_in(1883);
  VN314_in0 <= VN_sign_in(1884) & VN_data_in(1884);
  VN314_in1 <= VN_sign_in(1885) & VN_data_in(1885);
  VN314_in2 <= VN_sign_in(1886) & VN_data_in(1886);
  VN314_in3 <= VN_sign_in(1887) & VN_data_in(1887);
  VN314_in4 <= VN_sign_in(1888) & VN_data_in(1888);
  VN314_in5 <= VN_sign_in(1889) & VN_data_in(1889);
  VN315_in0 <= VN_sign_in(1890) & VN_data_in(1890);
  VN315_in1 <= VN_sign_in(1891) & VN_data_in(1891);
  VN315_in2 <= VN_sign_in(1892) & VN_data_in(1892);
  VN315_in3 <= VN_sign_in(1893) & VN_data_in(1893);
  VN315_in4 <= VN_sign_in(1894) & VN_data_in(1894);
  VN315_in5 <= VN_sign_in(1895) & VN_data_in(1895);
  VN316_in0 <= VN_sign_in(1896) & VN_data_in(1896);
  VN316_in1 <= VN_sign_in(1897) & VN_data_in(1897);
  VN316_in2 <= VN_sign_in(1898) & VN_data_in(1898);
  VN316_in3 <= VN_sign_in(1899) & VN_data_in(1899);
  VN316_in4 <= VN_sign_in(1900) & VN_data_in(1900);
  VN316_in5 <= VN_sign_in(1901) & VN_data_in(1901);
  VN317_in0 <= VN_sign_in(1902) & VN_data_in(1902);
  VN317_in1 <= VN_sign_in(1903) & VN_data_in(1903);
  VN317_in2 <= VN_sign_in(1904) & VN_data_in(1904);
  VN317_in3 <= VN_sign_in(1905) & VN_data_in(1905);
  VN317_in4 <= VN_sign_in(1906) & VN_data_in(1906);
  VN317_in5 <= VN_sign_in(1907) & VN_data_in(1907);
  VN318_in0 <= VN_sign_in(1908) & VN_data_in(1908);
  VN318_in1 <= VN_sign_in(1909) & VN_data_in(1909);
  VN318_in2 <= VN_sign_in(1910) & VN_data_in(1910);
  VN318_in3 <= VN_sign_in(1911) & VN_data_in(1911);
  VN318_in4 <= VN_sign_in(1912) & VN_data_in(1912);
  VN318_in5 <= VN_sign_in(1913) & VN_data_in(1913);
  VN319_in0 <= VN_sign_in(1914) & VN_data_in(1914);
  VN319_in1 <= VN_sign_in(1915) & VN_data_in(1915);
  VN319_in2 <= VN_sign_in(1916) & VN_data_in(1916);
  VN319_in3 <= VN_sign_in(1917) & VN_data_in(1917);
  VN319_in4 <= VN_sign_in(1918) & VN_data_in(1918);
  VN319_in5 <= VN_sign_in(1919) & VN_data_in(1919);
  VN320_in0 <= VN_sign_in(1920) & VN_data_in(1920);
  VN320_in1 <= VN_sign_in(1921) & VN_data_in(1921);
  VN320_in2 <= VN_sign_in(1922) & VN_data_in(1922);
  VN320_in3 <= VN_sign_in(1923) & VN_data_in(1923);
  VN320_in4 <= VN_sign_in(1924) & VN_data_in(1924);
  VN320_in5 <= VN_sign_in(1925) & VN_data_in(1925);
  VN321_in0 <= VN_sign_in(1926) & VN_data_in(1926);
  VN321_in1 <= VN_sign_in(1927) & VN_data_in(1927);
  VN321_in2 <= VN_sign_in(1928) & VN_data_in(1928);
  VN321_in3 <= VN_sign_in(1929) & VN_data_in(1929);
  VN321_in4 <= VN_sign_in(1930) & VN_data_in(1930);
  VN321_in5 <= VN_sign_in(1931) & VN_data_in(1931);
  VN322_in0 <= VN_sign_in(1932) & VN_data_in(1932);
  VN322_in1 <= VN_sign_in(1933) & VN_data_in(1933);
  VN322_in2 <= VN_sign_in(1934) & VN_data_in(1934);
  VN322_in3 <= VN_sign_in(1935) & VN_data_in(1935);
  VN322_in4 <= VN_sign_in(1936) & VN_data_in(1936);
  VN322_in5 <= VN_sign_in(1937) & VN_data_in(1937);
  VN323_in0 <= VN_sign_in(1938) & VN_data_in(1938);
  VN323_in1 <= VN_sign_in(1939) & VN_data_in(1939);
  VN323_in2 <= VN_sign_in(1940) & VN_data_in(1940);
  VN323_in3 <= VN_sign_in(1941) & VN_data_in(1941);
  VN323_in4 <= VN_sign_in(1942) & VN_data_in(1942);
  VN323_in5 <= VN_sign_in(1943) & VN_data_in(1943);
  VN324_in0 <= VN_sign_in(1944) & VN_data_in(1944);
  VN324_in1 <= VN_sign_in(1945) & VN_data_in(1945);
  VN324_in2 <= VN_sign_in(1946) & VN_data_in(1946);
  VN324_in3 <= VN_sign_in(1947) & VN_data_in(1947);
  VN324_in4 <= VN_sign_in(1948) & VN_data_in(1948);
  VN324_in5 <= VN_sign_in(1949) & VN_data_in(1949);
  VN325_in0 <= VN_sign_in(1950) & VN_data_in(1950);
  VN325_in1 <= VN_sign_in(1951) & VN_data_in(1951);
  VN325_in2 <= VN_sign_in(1952) & VN_data_in(1952);
  VN325_in3 <= VN_sign_in(1953) & VN_data_in(1953);
  VN325_in4 <= VN_sign_in(1954) & VN_data_in(1954);
  VN325_in5 <= VN_sign_in(1955) & VN_data_in(1955);
  VN326_in0 <= VN_sign_in(1956) & VN_data_in(1956);
  VN326_in1 <= VN_sign_in(1957) & VN_data_in(1957);
  VN326_in2 <= VN_sign_in(1958) & VN_data_in(1958);
  VN326_in3 <= VN_sign_in(1959) & VN_data_in(1959);
  VN326_in4 <= VN_sign_in(1960) & VN_data_in(1960);
  VN326_in5 <= VN_sign_in(1961) & VN_data_in(1961);
  VN327_in0 <= VN_sign_in(1962) & VN_data_in(1962);
  VN327_in1 <= VN_sign_in(1963) & VN_data_in(1963);
  VN327_in2 <= VN_sign_in(1964) & VN_data_in(1964);
  VN327_in3 <= VN_sign_in(1965) & VN_data_in(1965);
  VN327_in4 <= VN_sign_in(1966) & VN_data_in(1966);
  VN327_in5 <= VN_sign_in(1967) & VN_data_in(1967);
  VN328_in0 <= VN_sign_in(1968) & VN_data_in(1968);
  VN328_in1 <= VN_sign_in(1969) & VN_data_in(1969);
  VN328_in2 <= VN_sign_in(1970) & VN_data_in(1970);
  VN328_in3 <= VN_sign_in(1971) & VN_data_in(1971);
  VN328_in4 <= VN_sign_in(1972) & VN_data_in(1972);
  VN328_in5 <= VN_sign_in(1973) & VN_data_in(1973);
  VN329_in0 <= VN_sign_in(1974) & VN_data_in(1974);
  VN329_in1 <= VN_sign_in(1975) & VN_data_in(1975);
  VN329_in2 <= VN_sign_in(1976) & VN_data_in(1976);
  VN329_in3 <= VN_sign_in(1977) & VN_data_in(1977);
  VN329_in4 <= VN_sign_in(1978) & VN_data_in(1978);
  VN329_in5 <= VN_sign_in(1979) & VN_data_in(1979);
  VN330_in0 <= VN_sign_in(1980) & VN_data_in(1980);
  VN330_in1 <= VN_sign_in(1981) & VN_data_in(1981);
  VN330_in2 <= VN_sign_in(1982) & VN_data_in(1982);
  VN330_in3 <= VN_sign_in(1983) & VN_data_in(1983);
  VN330_in4 <= VN_sign_in(1984) & VN_data_in(1984);
  VN330_in5 <= VN_sign_in(1985) & VN_data_in(1985);
  VN331_in0 <= VN_sign_in(1986) & VN_data_in(1986);
  VN331_in1 <= VN_sign_in(1987) & VN_data_in(1987);
  VN331_in2 <= VN_sign_in(1988) & VN_data_in(1988);
  VN331_in3 <= VN_sign_in(1989) & VN_data_in(1989);
  VN331_in4 <= VN_sign_in(1990) & VN_data_in(1990);
  VN331_in5 <= VN_sign_in(1991) & VN_data_in(1991);
  VN332_in0 <= VN_sign_in(1992) & VN_data_in(1992);
  VN332_in1 <= VN_sign_in(1993) & VN_data_in(1993);
  VN332_in2 <= VN_sign_in(1994) & VN_data_in(1994);
  VN332_in3 <= VN_sign_in(1995) & VN_data_in(1995);
  VN332_in4 <= VN_sign_in(1996) & VN_data_in(1996);
  VN332_in5 <= VN_sign_in(1997) & VN_data_in(1997);
  VN333_in0 <= VN_sign_in(1998) & VN_data_in(1998);
  VN333_in1 <= VN_sign_in(1999) & VN_data_in(1999);
  VN333_in2 <= VN_sign_in(2000) & VN_data_in(2000);
  VN333_in3 <= VN_sign_in(2001) & VN_data_in(2001);
  VN333_in4 <= VN_sign_in(2002) & VN_data_in(2002);
  VN333_in5 <= VN_sign_in(2003) & VN_data_in(2003);
  VN334_in0 <= VN_sign_in(2004) & VN_data_in(2004);
  VN334_in1 <= VN_sign_in(2005) & VN_data_in(2005);
  VN334_in2 <= VN_sign_in(2006) & VN_data_in(2006);
  VN334_in3 <= VN_sign_in(2007) & VN_data_in(2007);
  VN334_in4 <= VN_sign_in(2008) & VN_data_in(2008);
  VN334_in5 <= VN_sign_in(2009) & VN_data_in(2009);
  VN335_in0 <= VN_sign_in(2010) & VN_data_in(2010);
  VN335_in1 <= VN_sign_in(2011) & VN_data_in(2011);
  VN335_in2 <= VN_sign_in(2012) & VN_data_in(2012);
  VN335_in3 <= VN_sign_in(2013) & VN_data_in(2013);
  VN335_in4 <= VN_sign_in(2014) & VN_data_in(2014);
  VN335_in5 <= VN_sign_in(2015) & VN_data_in(2015);
  VN336_in0 <= VN_sign_in(2016) & VN_data_in(2016);
  VN336_in1 <= VN_sign_in(2017) & VN_data_in(2017);
  VN336_in2 <= VN_sign_in(2018) & VN_data_in(2018);
  VN336_in3 <= VN_sign_in(2019) & VN_data_in(2019);
  VN336_in4 <= VN_sign_in(2020) & VN_data_in(2020);
  VN336_in5 <= VN_sign_in(2021) & VN_data_in(2021);
  VN337_in0 <= VN_sign_in(2022) & VN_data_in(2022);
  VN337_in1 <= VN_sign_in(2023) & VN_data_in(2023);
  VN337_in2 <= VN_sign_in(2024) & VN_data_in(2024);
  VN337_in3 <= VN_sign_in(2025) & VN_data_in(2025);
  VN337_in4 <= VN_sign_in(2026) & VN_data_in(2026);
  VN337_in5 <= VN_sign_in(2027) & VN_data_in(2027);
  VN338_in0 <= VN_sign_in(2028) & VN_data_in(2028);
  VN338_in1 <= VN_sign_in(2029) & VN_data_in(2029);
  VN338_in2 <= VN_sign_in(2030) & VN_data_in(2030);
  VN338_in3 <= VN_sign_in(2031) & VN_data_in(2031);
  VN338_in4 <= VN_sign_in(2032) & VN_data_in(2032);
  VN338_in5 <= VN_sign_in(2033) & VN_data_in(2033);
  VN339_in0 <= VN_sign_in(2034) & VN_data_in(2034);
  VN339_in1 <= VN_sign_in(2035) & VN_data_in(2035);
  VN339_in2 <= VN_sign_in(2036) & VN_data_in(2036);
  VN339_in3 <= VN_sign_in(2037) & VN_data_in(2037);
  VN339_in4 <= VN_sign_in(2038) & VN_data_in(2038);
  VN339_in5 <= VN_sign_in(2039) & VN_data_in(2039);
  VN340_in0 <= VN_sign_in(2040) & VN_data_in(2040);
  VN340_in1 <= VN_sign_in(2041) & VN_data_in(2041);
  VN340_in2 <= VN_sign_in(2042) & VN_data_in(2042);
  VN340_in3 <= VN_sign_in(2043) & VN_data_in(2043);
  VN340_in4 <= VN_sign_in(2044) & VN_data_in(2044);
  VN340_in5 <= VN_sign_in(2045) & VN_data_in(2045);
  VN341_in0 <= VN_sign_in(2046) & VN_data_in(2046);
  VN341_in1 <= VN_sign_in(2047) & VN_data_in(2047);
  VN341_in2 <= VN_sign_in(2048) & VN_data_in(2048);
  VN341_in3 <= VN_sign_in(2049) & VN_data_in(2049);
  VN341_in4 <= VN_sign_in(2050) & VN_data_in(2050);
  VN341_in5 <= VN_sign_in(2051) & VN_data_in(2051);
  VN342_in0 <= VN_sign_in(2052) & VN_data_in(2052);
  VN342_in1 <= VN_sign_in(2053) & VN_data_in(2053);
  VN342_in2 <= VN_sign_in(2054) & VN_data_in(2054);
  VN342_in3 <= VN_sign_in(2055) & VN_data_in(2055);
  VN342_in4 <= VN_sign_in(2056) & VN_data_in(2056);
  VN342_in5 <= VN_sign_in(2057) & VN_data_in(2057);
  VN343_in0 <= VN_sign_in(2058) & VN_data_in(2058);
  VN343_in1 <= VN_sign_in(2059) & VN_data_in(2059);
  VN343_in2 <= VN_sign_in(2060) & VN_data_in(2060);
  VN343_in3 <= VN_sign_in(2061) & VN_data_in(2061);
  VN343_in4 <= VN_sign_in(2062) & VN_data_in(2062);
  VN343_in5 <= VN_sign_in(2063) & VN_data_in(2063);
  VN344_in0 <= VN_sign_in(2064) & VN_data_in(2064);
  VN344_in1 <= VN_sign_in(2065) & VN_data_in(2065);
  VN344_in2 <= VN_sign_in(2066) & VN_data_in(2066);
  VN344_in3 <= VN_sign_in(2067) & VN_data_in(2067);
  VN344_in4 <= VN_sign_in(2068) & VN_data_in(2068);
  VN344_in5 <= VN_sign_in(2069) & VN_data_in(2069);
  VN345_in0 <= VN_sign_in(2070) & VN_data_in(2070);
  VN345_in1 <= VN_sign_in(2071) & VN_data_in(2071);
  VN345_in2 <= VN_sign_in(2072) & VN_data_in(2072);
  VN345_in3 <= VN_sign_in(2073) & VN_data_in(2073);
  VN345_in4 <= VN_sign_in(2074) & VN_data_in(2074);
  VN345_in5 <= VN_sign_in(2075) & VN_data_in(2075);
  VN346_in0 <= VN_sign_in(2076) & VN_data_in(2076);
  VN346_in1 <= VN_sign_in(2077) & VN_data_in(2077);
  VN346_in2 <= VN_sign_in(2078) & VN_data_in(2078);
  VN346_in3 <= VN_sign_in(2079) & VN_data_in(2079);
  VN346_in4 <= VN_sign_in(2080) & VN_data_in(2080);
  VN346_in5 <= VN_sign_in(2081) & VN_data_in(2081);
  VN347_in0 <= VN_sign_in(2082) & VN_data_in(2082);
  VN347_in1 <= VN_sign_in(2083) & VN_data_in(2083);
  VN347_in2 <= VN_sign_in(2084) & VN_data_in(2084);
  VN347_in3 <= VN_sign_in(2085) & VN_data_in(2085);
  VN347_in4 <= VN_sign_in(2086) & VN_data_in(2086);
  VN347_in5 <= VN_sign_in(2087) & VN_data_in(2087);
  VN348_in0 <= VN_sign_in(2088) & VN_data_in(2088);
  VN348_in1 <= VN_sign_in(2089) & VN_data_in(2089);
  VN348_in2 <= VN_sign_in(2090) & VN_data_in(2090);
  VN348_in3 <= VN_sign_in(2091) & VN_data_in(2091);
  VN348_in4 <= VN_sign_in(2092) & VN_data_in(2092);
  VN348_in5 <= VN_sign_in(2093) & VN_data_in(2093);
  VN349_in0 <= VN_sign_in(2094) & VN_data_in(2094);
  VN349_in1 <= VN_sign_in(2095) & VN_data_in(2095);
  VN349_in2 <= VN_sign_in(2096) & VN_data_in(2096);
  VN349_in3 <= VN_sign_in(2097) & VN_data_in(2097);
  VN349_in4 <= VN_sign_in(2098) & VN_data_in(2098);
  VN349_in5 <= VN_sign_in(2099) & VN_data_in(2099);
  VN350_in0 <= VN_sign_in(2100) & VN_data_in(2100);
  VN350_in1 <= VN_sign_in(2101) & VN_data_in(2101);
  VN350_in2 <= VN_sign_in(2102) & VN_data_in(2102);
  VN350_in3 <= VN_sign_in(2103) & VN_data_in(2103);
  VN350_in4 <= VN_sign_in(2104) & VN_data_in(2104);
  VN350_in5 <= VN_sign_in(2105) & VN_data_in(2105);
  VN351_in0 <= VN_sign_in(2106) & VN_data_in(2106);
  VN351_in1 <= VN_sign_in(2107) & VN_data_in(2107);
  VN351_in2 <= VN_sign_in(2108) & VN_data_in(2108);
  VN351_in3 <= VN_sign_in(2109) & VN_data_in(2109);
  VN351_in4 <= VN_sign_in(2110) & VN_data_in(2110);
  VN351_in5 <= VN_sign_in(2111) & VN_data_in(2111);
  VN352_in0 <= VN_sign_in(2112) & VN_data_in(2112);
  VN352_in1 <= VN_sign_in(2113) & VN_data_in(2113);
  VN352_in2 <= VN_sign_in(2114) & VN_data_in(2114);
  VN352_in3 <= VN_sign_in(2115) & VN_data_in(2115);
  VN352_in4 <= VN_sign_in(2116) & VN_data_in(2116);
  VN352_in5 <= VN_sign_in(2117) & VN_data_in(2117);
  VN353_in0 <= VN_sign_in(2118) & VN_data_in(2118);
  VN353_in1 <= VN_sign_in(2119) & VN_data_in(2119);
  VN353_in2 <= VN_sign_in(2120) & VN_data_in(2120);
  VN353_in3 <= VN_sign_in(2121) & VN_data_in(2121);
  VN353_in4 <= VN_sign_in(2122) & VN_data_in(2122);
  VN353_in5 <= VN_sign_in(2123) & VN_data_in(2123);
  VN354_in0 <= VN_sign_in(2124) & VN_data_in(2124);
  VN354_in1 <= VN_sign_in(2125) & VN_data_in(2125);
  VN354_in2 <= VN_sign_in(2126) & VN_data_in(2126);
  VN354_in3 <= VN_sign_in(2127) & VN_data_in(2127);
  VN354_in4 <= VN_sign_in(2128) & VN_data_in(2128);
  VN354_in5 <= VN_sign_in(2129) & VN_data_in(2129);
  VN355_in0 <= VN_sign_in(2130) & VN_data_in(2130);
  VN355_in1 <= VN_sign_in(2131) & VN_data_in(2131);
  VN355_in2 <= VN_sign_in(2132) & VN_data_in(2132);
  VN355_in3 <= VN_sign_in(2133) & VN_data_in(2133);
  VN355_in4 <= VN_sign_in(2134) & VN_data_in(2134);
  VN355_in5 <= VN_sign_in(2135) & VN_data_in(2135);
  VN356_in0 <= VN_sign_in(2136) & VN_data_in(2136);
  VN356_in1 <= VN_sign_in(2137) & VN_data_in(2137);
  VN356_in2 <= VN_sign_in(2138) & VN_data_in(2138);
  VN356_in3 <= VN_sign_in(2139) & VN_data_in(2139);
  VN356_in4 <= VN_sign_in(2140) & VN_data_in(2140);
  VN356_in5 <= VN_sign_in(2141) & VN_data_in(2141);
  VN357_in0 <= VN_sign_in(2142) & VN_data_in(2142);
  VN357_in1 <= VN_sign_in(2143) & VN_data_in(2143);
  VN357_in2 <= VN_sign_in(2144) & VN_data_in(2144);
  VN357_in3 <= VN_sign_in(2145) & VN_data_in(2145);
  VN357_in4 <= VN_sign_in(2146) & VN_data_in(2146);
  VN357_in5 <= VN_sign_in(2147) & VN_data_in(2147);
  VN358_in0 <= VN_sign_in(2148) & VN_data_in(2148);
  VN358_in1 <= VN_sign_in(2149) & VN_data_in(2149);
  VN358_in2 <= VN_sign_in(2150) & VN_data_in(2150);
  VN358_in3 <= VN_sign_in(2151) & VN_data_in(2151);
  VN358_in4 <= VN_sign_in(2152) & VN_data_in(2152);
  VN358_in5 <= VN_sign_in(2153) & VN_data_in(2153);
  VN359_in0 <= VN_sign_in(2154) & VN_data_in(2154);
  VN359_in1 <= VN_sign_in(2155) & VN_data_in(2155);
  VN359_in2 <= VN_sign_in(2156) & VN_data_in(2156);
  VN359_in3 <= VN_sign_in(2157) & VN_data_in(2157);
  VN359_in4 <= VN_sign_in(2158) & VN_data_in(2158);
  VN359_in5 <= VN_sign_in(2159) & VN_data_in(2159);
  VN360_in0 <= VN_sign_in(2160) & VN_data_in(2160);
  VN360_in1 <= VN_sign_in(2161) & VN_data_in(2161);
  VN360_in2 <= VN_sign_in(2162) & VN_data_in(2162);
  VN360_in3 <= VN_sign_in(2163) & VN_data_in(2163);
  VN360_in4 <= VN_sign_in(2164) & VN_data_in(2164);
  VN360_in5 <= VN_sign_in(2165) & VN_data_in(2165);
  VN361_in0 <= VN_sign_in(2166) & VN_data_in(2166);
  VN361_in1 <= VN_sign_in(2167) & VN_data_in(2167);
  VN361_in2 <= VN_sign_in(2168) & VN_data_in(2168);
  VN361_in3 <= VN_sign_in(2169) & VN_data_in(2169);
  VN361_in4 <= VN_sign_in(2170) & VN_data_in(2170);
  VN361_in5 <= VN_sign_in(2171) & VN_data_in(2171);
  VN362_in0 <= VN_sign_in(2172) & VN_data_in(2172);
  VN362_in1 <= VN_sign_in(2173) & VN_data_in(2173);
  VN362_in2 <= VN_sign_in(2174) & VN_data_in(2174);
  VN362_in3 <= VN_sign_in(2175) & VN_data_in(2175);
  VN362_in4 <= VN_sign_in(2176) & VN_data_in(2176);
  VN362_in5 <= VN_sign_in(2177) & VN_data_in(2177);
  VN363_in0 <= VN_sign_in(2178) & VN_data_in(2178);
  VN363_in1 <= VN_sign_in(2179) & VN_data_in(2179);
  VN363_in2 <= VN_sign_in(2180) & VN_data_in(2180);
  VN363_in3 <= VN_sign_in(2181) & VN_data_in(2181);
  VN363_in4 <= VN_sign_in(2182) & VN_data_in(2182);
  VN363_in5 <= VN_sign_in(2183) & VN_data_in(2183);
  VN364_in0 <= VN_sign_in(2184) & VN_data_in(2184);
  VN364_in1 <= VN_sign_in(2185) & VN_data_in(2185);
  VN364_in2 <= VN_sign_in(2186) & VN_data_in(2186);
  VN364_in3 <= VN_sign_in(2187) & VN_data_in(2187);
  VN364_in4 <= VN_sign_in(2188) & VN_data_in(2188);
  VN364_in5 <= VN_sign_in(2189) & VN_data_in(2189);
  VN365_in0 <= VN_sign_in(2190) & VN_data_in(2190);
  VN365_in1 <= VN_sign_in(2191) & VN_data_in(2191);
  VN365_in2 <= VN_sign_in(2192) & VN_data_in(2192);
  VN365_in3 <= VN_sign_in(2193) & VN_data_in(2193);
  VN365_in4 <= VN_sign_in(2194) & VN_data_in(2194);
  VN365_in5 <= VN_sign_in(2195) & VN_data_in(2195);
  VN366_in0 <= VN_sign_in(2196) & VN_data_in(2196);
  VN366_in1 <= VN_sign_in(2197) & VN_data_in(2197);
  VN366_in2 <= VN_sign_in(2198) & VN_data_in(2198);
  VN366_in3 <= VN_sign_in(2199) & VN_data_in(2199);
  VN366_in4 <= VN_sign_in(2200) & VN_data_in(2200);
  VN366_in5 <= VN_sign_in(2201) & VN_data_in(2201);
  VN367_in0 <= VN_sign_in(2202) & VN_data_in(2202);
  VN367_in1 <= VN_sign_in(2203) & VN_data_in(2203);
  VN367_in2 <= VN_sign_in(2204) & VN_data_in(2204);
  VN367_in3 <= VN_sign_in(2205) & VN_data_in(2205);
  VN367_in4 <= VN_sign_in(2206) & VN_data_in(2206);
  VN367_in5 <= VN_sign_in(2207) & VN_data_in(2207);
  VN368_in0 <= VN_sign_in(2208) & VN_data_in(2208);
  VN368_in1 <= VN_sign_in(2209) & VN_data_in(2209);
  VN368_in2 <= VN_sign_in(2210) & VN_data_in(2210);
  VN368_in3 <= VN_sign_in(2211) & VN_data_in(2211);
  VN368_in4 <= VN_sign_in(2212) & VN_data_in(2212);
  VN368_in5 <= VN_sign_in(2213) & VN_data_in(2213);
  VN369_in0 <= VN_sign_in(2214) & VN_data_in(2214);
  VN369_in1 <= VN_sign_in(2215) & VN_data_in(2215);
  VN369_in2 <= VN_sign_in(2216) & VN_data_in(2216);
  VN369_in3 <= VN_sign_in(2217) & VN_data_in(2217);
  VN369_in4 <= VN_sign_in(2218) & VN_data_in(2218);
  VN369_in5 <= VN_sign_in(2219) & VN_data_in(2219);
  VN370_in0 <= VN_sign_in(2220) & VN_data_in(2220);
  VN370_in1 <= VN_sign_in(2221) & VN_data_in(2221);
  VN370_in2 <= VN_sign_in(2222) & VN_data_in(2222);
  VN370_in3 <= VN_sign_in(2223) & VN_data_in(2223);
  VN370_in4 <= VN_sign_in(2224) & VN_data_in(2224);
  VN370_in5 <= VN_sign_in(2225) & VN_data_in(2225);
  VN371_in0 <= VN_sign_in(2226) & VN_data_in(2226);
  VN371_in1 <= VN_sign_in(2227) & VN_data_in(2227);
  VN371_in2 <= VN_sign_in(2228) & VN_data_in(2228);
  VN371_in3 <= VN_sign_in(2229) & VN_data_in(2229);
  VN371_in4 <= VN_sign_in(2230) & VN_data_in(2230);
  VN371_in5 <= VN_sign_in(2231) & VN_data_in(2231);
  VN372_in0 <= VN_sign_in(2232) & VN_data_in(2232);
  VN372_in1 <= VN_sign_in(2233) & VN_data_in(2233);
  VN372_in2 <= VN_sign_in(2234) & VN_data_in(2234);
  VN372_in3 <= VN_sign_in(2235) & VN_data_in(2235);
  VN372_in4 <= VN_sign_in(2236) & VN_data_in(2236);
  VN372_in5 <= VN_sign_in(2237) & VN_data_in(2237);
  VN373_in0 <= VN_sign_in(2238) & VN_data_in(2238);
  VN373_in1 <= VN_sign_in(2239) & VN_data_in(2239);
  VN373_in2 <= VN_sign_in(2240) & VN_data_in(2240);
  VN373_in3 <= VN_sign_in(2241) & VN_data_in(2241);
  VN373_in4 <= VN_sign_in(2242) & VN_data_in(2242);
  VN373_in5 <= VN_sign_in(2243) & VN_data_in(2243);
  VN374_in0 <= VN_sign_in(2244) & VN_data_in(2244);
  VN374_in1 <= VN_sign_in(2245) & VN_data_in(2245);
  VN374_in2 <= VN_sign_in(2246) & VN_data_in(2246);
  VN374_in3 <= VN_sign_in(2247) & VN_data_in(2247);
  VN374_in4 <= VN_sign_in(2248) & VN_data_in(2248);
  VN374_in5 <= VN_sign_in(2249) & VN_data_in(2249);
  VN375_in0 <= VN_sign_in(2250) & VN_data_in(2250);
  VN375_in1 <= VN_sign_in(2251) & VN_data_in(2251);
  VN375_in2 <= VN_sign_in(2252) & VN_data_in(2252);
  VN375_in3 <= VN_sign_in(2253) & VN_data_in(2253);
  VN375_in4 <= VN_sign_in(2254) & VN_data_in(2254);
  VN375_in5 <= VN_sign_in(2255) & VN_data_in(2255);
  VN376_in0 <= VN_sign_in(2256) & VN_data_in(2256);
  VN376_in1 <= VN_sign_in(2257) & VN_data_in(2257);
  VN376_in2 <= VN_sign_in(2258) & VN_data_in(2258);
  VN376_in3 <= VN_sign_in(2259) & VN_data_in(2259);
  VN376_in4 <= VN_sign_in(2260) & VN_data_in(2260);
  VN376_in5 <= VN_sign_in(2261) & VN_data_in(2261);
  VN377_in0 <= VN_sign_in(2262) & VN_data_in(2262);
  VN377_in1 <= VN_sign_in(2263) & VN_data_in(2263);
  VN377_in2 <= VN_sign_in(2264) & VN_data_in(2264);
  VN377_in3 <= VN_sign_in(2265) & VN_data_in(2265);
  VN377_in4 <= VN_sign_in(2266) & VN_data_in(2266);
  VN377_in5 <= VN_sign_in(2267) & VN_data_in(2267);
  VN378_in0 <= VN_sign_in(2268) & VN_data_in(2268);
  VN378_in1 <= VN_sign_in(2269) & VN_data_in(2269);
  VN378_in2 <= VN_sign_in(2270) & VN_data_in(2270);
  VN378_in3 <= VN_sign_in(2271) & VN_data_in(2271);
  VN378_in4 <= VN_sign_in(2272) & VN_data_in(2272);
  VN378_in5 <= VN_sign_in(2273) & VN_data_in(2273);
  VN379_in0 <= VN_sign_in(2274) & VN_data_in(2274);
  VN379_in1 <= VN_sign_in(2275) & VN_data_in(2275);
  VN379_in2 <= VN_sign_in(2276) & VN_data_in(2276);
  VN379_in3 <= VN_sign_in(2277) & VN_data_in(2277);
  VN379_in4 <= VN_sign_in(2278) & VN_data_in(2278);
  VN379_in5 <= VN_sign_in(2279) & VN_data_in(2279);
  VN380_in0 <= VN_sign_in(2280) & VN_data_in(2280);
  VN380_in1 <= VN_sign_in(2281) & VN_data_in(2281);
  VN380_in2 <= VN_sign_in(2282) & VN_data_in(2282);
  VN380_in3 <= VN_sign_in(2283) & VN_data_in(2283);
  VN380_in4 <= VN_sign_in(2284) & VN_data_in(2284);
  VN380_in5 <= VN_sign_in(2285) & VN_data_in(2285);
  VN381_in0 <= VN_sign_in(2286) & VN_data_in(2286);
  VN381_in1 <= VN_sign_in(2287) & VN_data_in(2287);
  VN381_in2 <= VN_sign_in(2288) & VN_data_in(2288);
  VN381_in3 <= VN_sign_in(2289) & VN_data_in(2289);
  VN381_in4 <= VN_sign_in(2290) & VN_data_in(2290);
  VN381_in5 <= VN_sign_in(2291) & VN_data_in(2291);
  VN382_in0 <= VN_sign_in(2292) & VN_data_in(2292);
  VN382_in1 <= VN_sign_in(2293) & VN_data_in(2293);
  VN382_in2 <= VN_sign_in(2294) & VN_data_in(2294);
  VN382_in3 <= VN_sign_in(2295) & VN_data_in(2295);
  VN382_in4 <= VN_sign_in(2296) & VN_data_in(2296);
  VN382_in5 <= VN_sign_in(2297) & VN_data_in(2297);
  VN383_in0 <= VN_sign_in(2298) & VN_data_in(2298);
  VN383_in1 <= VN_sign_in(2299) & VN_data_in(2299);
  VN383_in2 <= VN_sign_in(2300) & VN_data_in(2300);
  VN383_in3 <= VN_sign_in(2301) & VN_data_in(2301);
  VN383_in4 <= VN_sign_in(2302) & VN_data_in(2302);
  VN383_in5 <= VN_sign_in(2303) & VN_data_in(2303);
  VN384_in0 <= VN_sign_in(2304) & VN_data_in(2304);
  VN384_in1 <= VN_sign_in(2305) & VN_data_in(2305);
  VN384_in2 <= VN_sign_in(2306) & VN_data_in(2306);
  VN384_in3 <= VN_sign_in(2307) & VN_data_in(2307);
  VN384_in4 <= VN_sign_in(2308) & VN_data_in(2308);
  VN384_in5 <= VN_sign_in(2309) & VN_data_in(2309);
  VN385_in0 <= VN_sign_in(2310) & VN_data_in(2310);
  VN385_in1 <= VN_sign_in(2311) & VN_data_in(2311);
  VN385_in2 <= VN_sign_in(2312) & VN_data_in(2312);
  VN385_in3 <= VN_sign_in(2313) & VN_data_in(2313);
  VN385_in4 <= VN_sign_in(2314) & VN_data_in(2314);
  VN385_in5 <= VN_sign_in(2315) & VN_data_in(2315);
  VN386_in0 <= VN_sign_in(2316) & VN_data_in(2316);
  VN386_in1 <= VN_sign_in(2317) & VN_data_in(2317);
  VN386_in2 <= VN_sign_in(2318) & VN_data_in(2318);
  VN386_in3 <= VN_sign_in(2319) & VN_data_in(2319);
  VN386_in4 <= VN_sign_in(2320) & VN_data_in(2320);
  VN386_in5 <= VN_sign_in(2321) & VN_data_in(2321);
  VN387_in0 <= VN_sign_in(2322) & VN_data_in(2322);
  VN387_in1 <= VN_sign_in(2323) & VN_data_in(2323);
  VN387_in2 <= VN_sign_in(2324) & VN_data_in(2324);
  VN387_in3 <= VN_sign_in(2325) & VN_data_in(2325);
  VN387_in4 <= VN_sign_in(2326) & VN_data_in(2326);
  VN387_in5 <= VN_sign_in(2327) & VN_data_in(2327);
  VN388_in0 <= VN_sign_in(2328) & VN_data_in(2328);
  VN388_in1 <= VN_sign_in(2329) & VN_data_in(2329);
  VN388_in2 <= VN_sign_in(2330) & VN_data_in(2330);
  VN388_in3 <= VN_sign_in(2331) & VN_data_in(2331);
  VN388_in4 <= VN_sign_in(2332) & VN_data_in(2332);
  VN388_in5 <= VN_sign_in(2333) & VN_data_in(2333);
  VN389_in0 <= VN_sign_in(2334) & VN_data_in(2334);
  VN389_in1 <= VN_sign_in(2335) & VN_data_in(2335);
  VN389_in2 <= VN_sign_in(2336) & VN_data_in(2336);
  VN389_in3 <= VN_sign_in(2337) & VN_data_in(2337);
  VN389_in4 <= VN_sign_in(2338) & VN_data_in(2338);
  VN389_in5 <= VN_sign_in(2339) & VN_data_in(2339);
  VN390_in0 <= VN_sign_in(2340) & VN_data_in(2340);
  VN390_in1 <= VN_sign_in(2341) & VN_data_in(2341);
  VN390_in2 <= VN_sign_in(2342) & VN_data_in(2342);
  VN390_in3 <= VN_sign_in(2343) & VN_data_in(2343);
  VN390_in4 <= VN_sign_in(2344) & VN_data_in(2344);
  VN390_in5 <= VN_sign_in(2345) & VN_data_in(2345);
  VN391_in0 <= VN_sign_in(2346) & VN_data_in(2346);
  VN391_in1 <= VN_sign_in(2347) & VN_data_in(2347);
  VN391_in2 <= VN_sign_in(2348) & VN_data_in(2348);
  VN391_in3 <= VN_sign_in(2349) & VN_data_in(2349);
  VN391_in4 <= VN_sign_in(2350) & VN_data_in(2350);
  VN391_in5 <= VN_sign_in(2351) & VN_data_in(2351);
  VN392_in0 <= VN_sign_in(2352) & VN_data_in(2352);
  VN392_in1 <= VN_sign_in(2353) & VN_data_in(2353);
  VN392_in2 <= VN_sign_in(2354) & VN_data_in(2354);
  VN392_in3 <= VN_sign_in(2355) & VN_data_in(2355);
  VN392_in4 <= VN_sign_in(2356) & VN_data_in(2356);
  VN392_in5 <= VN_sign_in(2357) & VN_data_in(2357);
  VN393_in0 <= VN_sign_in(2358) & VN_data_in(2358);
  VN393_in1 <= VN_sign_in(2359) & VN_data_in(2359);
  VN393_in2 <= VN_sign_in(2360) & VN_data_in(2360);
  VN393_in3 <= VN_sign_in(2361) & VN_data_in(2361);
  VN393_in4 <= VN_sign_in(2362) & VN_data_in(2362);
  VN393_in5 <= VN_sign_in(2363) & VN_data_in(2363);
  VN394_in0 <= VN_sign_in(2364) & VN_data_in(2364);
  VN394_in1 <= VN_sign_in(2365) & VN_data_in(2365);
  VN394_in2 <= VN_sign_in(2366) & VN_data_in(2366);
  VN394_in3 <= VN_sign_in(2367) & VN_data_in(2367);
  VN394_in4 <= VN_sign_in(2368) & VN_data_in(2368);
  VN394_in5 <= VN_sign_in(2369) & VN_data_in(2369);
  VN395_in0 <= VN_sign_in(2370) & VN_data_in(2370);
  VN395_in1 <= VN_sign_in(2371) & VN_data_in(2371);
  VN395_in2 <= VN_sign_in(2372) & VN_data_in(2372);
  VN395_in3 <= VN_sign_in(2373) & VN_data_in(2373);
  VN395_in4 <= VN_sign_in(2374) & VN_data_in(2374);
  VN395_in5 <= VN_sign_in(2375) & VN_data_in(2375);
  VN396_in0 <= VN_sign_in(2376) & VN_data_in(2376);
  VN396_in1 <= VN_sign_in(2377) & VN_data_in(2377);
  VN396_in2 <= VN_sign_in(2378) & VN_data_in(2378);
  VN396_in3 <= VN_sign_in(2379) & VN_data_in(2379);
  VN396_in4 <= VN_sign_in(2380) & VN_data_in(2380);
  VN396_in5 <= VN_sign_in(2381) & VN_data_in(2381);
  VN397_in0 <= VN_sign_in(2382) & VN_data_in(2382);
  VN397_in1 <= VN_sign_in(2383) & VN_data_in(2383);
  VN397_in2 <= VN_sign_in(2384) & VN_data_in(2384);
  VN397_in3 <= VN_sign_in(2385) & VN_data_in(2385);
  VN397_in4 <= VN_sign_in(2386) & VN_data_in(2386);
  VN397_in5 <= VN_sign_in(2387) & VN_data_in(2387);
  VN398_in0 <= VN_sign_in(2388) & VN_data_in(2388);
  VN398_in1 <= VN_sign_in(2389) & VN_data_in(2389);
  VN398_in2 <= VN_sign_in(2390) & VN_data_in(2390);
  VN398_in3 <= VN_sign_in(2391) & VN_data_in(2391);
  VN398_in4 <= VN_sign_in(2392) & VN_data_in(2392);
  VN398_in5 <= VN_sign_in(2393) & VN_data_in(2393);
  VN399_in0 <= VN_sign_in(2394) & VN_data_in(2394);
  VN399_in1 <= VN_sign_in(2395) & VN_data_in(2395);
  VN399_in2 <= VN_sign_in(2396) & VN_data_in(2396);
  VN399_in3 <= VN_sign_in(2397) & VN_data_in(2397);
  VN399_in4 <= VN_sign_in(2398) & VN_data_in(2398);
  VN399_in5 <= VN_sign_in(2399) & VN_data_in(2399);
  VN400_in0 <= VN_sign_in(2400) & VN_data_in(2400);
  VN400_in1 <= VN_sign_in(2401) & VN_data_in(2401);
  VN400_in2 <= VN_sign_in(2402) & VN_data_in(2402);
  VN400_in3 <= VN_sign_in(2403) & VN_data_in(2403);
  VN400_in4 <= VN_sign_in(2404) & VN_data_in(2404);
  VN400_in5 <= VN_sign_in(2405) & VN_data_in(2405);
  VN401_in0 <= VN_sign_in(2406) & VN_data_in(2406);
  VN401_in1 <= VN_sign_in(2407) & VN_data_in(2407);
  VN401_in2 <= VN_sign_in(2408) & VN_data_in(2408);
  VN401_in3 <= VN_sign_in(2409) & VN_data_in(2409);
  VN401_in4 <= VN_sign_in(2410) & VN_data_in(2410);
  VN401_in5 <= VN_sign_in(2411) & VN_data_in(2411);
  VN402_in0 <= VN_sign_in(2412) & VN_data_in(2412);
  VN402_in1 <= VN_sign_in(2413) & VN_data_in(2413);
  VN402_in2 <= VN_sign_in(2414) & VN_data_in(2414);
  VN402_in3 <= VN_sign_in(2415) & VN_data_in(2415);
  VN402_in4 <= VN_sign_in(2416) & VN_data_in(2416);
  VN402_in5 <= VN_sign_in(2417) & VN_data_in(2417);
  VN403_in0 <= VN_sign_in(2418) & VN_data_in(2418);
  VN403_in1 <= VN_sign_in(2419) & VN_data_in(2419);
  VN403_in2 <= VN_sign_in(2420) & VN_data_in(2420);
  VN403_in3 <= VN_sign_in(2421) & VN_data_in(2421);
  VN403_in4 <= VN_sign_in(2422) & VN_data_in(2422);
  VN403_in5 <= VN_sign_in(2423) & VN_data_in(2423);
  VN404_in0 <= VN_sign_in(2424) & VN_data_in(2424);
  VN404_in1 <= VN_sign_in(2425) & VN_data_in(2425);
  VN404_in2 <= VN_sign_in(2426) & VN_data_in(2426);
  VN404_in3 <= VN_sign_in(2427) & VN_data_in(2427);
  VN404_in4 <= VN_sign_in(2428) & VN_data_in(2428);
  VN404_in5 <= VN_sign_in(2429) & VN_data_in(2429);
  VN405_in0 <= VN_sign_in(2430) & VN_data_in(2430);
  VN405_in1 <= VN_sign_in(2431) & VN_data_in(2431);
  VN405_in2 <= VN_sign_in(2432) & VN_data_in(2432);
  VN405_in3 <= VN_sign_in(2433) & VN_data_in(2433);
  VN405_in4 <= VN_sign_in(2434) & VN_data_in(2434);
  VN405_in5 <= VN_sign_in(2435) & VN_data_in(2435);
  VN406_in0 <= VN_sign_in(2436) & VN_data_in(2436);
  VN406_in1 <= VN_sign_in(2437) & VN_data_in(2437);
  VN406_in2 <= VN_sign_in(2438) & VN_data_in(2438);
  VN406_in3 <= VN_sign_in(2439) & VN_data_in(2439);
  VN406_in4 <= VN_sign_in(2440) & VN_data_in(2440);
  VN406_in5 <= VN_sign_in(2441) & VN_data_in(2441);
  VN407_in0 <= VN_sign_in(2442) & VN_data_in(2442);
  VN407_in1 <= VN_sign_in(2443) & VN_data_in(2443);
  VN407_in2 <= VN_sign_in(2444) & VN_data_in(2444);
  VN407_in3 <= VN_sign_in(2445) & VN_data_in(2445);
  VN407_in4 <= VN_sign_in(2446) & VN_data_in(2446);
  VN407_in5 <= VN_sign_in(2447) & VN_data_in(2447);
  VN408_in0 <= VN_sign_in(2448) & VN_data_in(2448);
  VN408_in1 <= VN_sign_in(2449) & VN_data_in(2449);
  VN408_in2 <= VN_sign_in(2450) & VN_data_in(2450);
  VN408_in3 <= VN_sign_in(2451) & VN_data_in(2451);
  VN408_in4 <= VN_sign_in(2452) & VN_data_in(2452);
  VN408_in5 <= VN_sign_in(2453) & VN_data_in(2453);
  VN409_in0 <= VN_sign_in(2454) & VN_data_in(2454);
  VN409_in1 <= VN_sign_in(2455) & VN_data_in(2455);
  VN409_in2 <= VN_sign_in(2456) & VN_data_in(2456);
  VN409_in3 <= VN_sign_in(2457) & VN_data_in(2457);
  VN409_in4 <= VN_sign_in(2458) & VN_data_in(2458);
  VN409_in5 <= VN_sign_in(2459) & VN_data_in(2459);
  VN410_in0 <= VN_sign_in(2460) & VN_data_in(2460);
  VN410_in1 <= VN_sign_in(2461) & VN_data_in(2461);
  VN410_in2 <= VN_sign_in(2462) & VN_data_in(2462);
  VN410_in3 <= VN_sign_in(2463) & VN_data_in(2463);
  VN410_in4 <= VN_sign_in(2464) & VN_data_in(2464);
  VN410_in5 <= VN_sign_in(2465) & VN_data_in(2465);
  VN411_in0 <= VN_sign_in(2466) & VN_data_in(2466);
  VN411_in1 <= VN_sign_in(2467) & VN_data_in(2467);
  VN411_in2 <= VN_sign_in(2468) & VN_data_in(2468);
  VN411_in3 <= VN_sign_in(2469) & VN_data_in(2469);
  VN411_in4 <= VN_sign_in(2470) & VN_data_in(2470);
  VN411_in5 <= VN_sign_in(2471) & VN_data_in(2471);
  VN412_in0 <= VN_sign_in(2472) & VN_data_in(2472);
  VN412_in1 <= VN_sign_in(2473) & VN_data_in(2473);
  VN412_in2 <= VN_sign_in(2474) & VN_data_in(2474);
  VN412_in3 <= VN_sign_in(2475) & VN_data_in(2475);
  VN412_in4 <= VN_sign_in(2476) & VN_data_in(2476);
  VN412_in5 <= VN_sign_in(2477) & VN_data_in(2477);
  VN413_in0 <= VN_sign_in(2478) & VN_data_in(2478);
  VN413_in1 <= VN_sign_in(2479) & VN_data_in(2479);
  VN413_in2 <= VN_sign_in(2480) & VN_data_in(2480);
  VN413_in3 <= VN_sign_in(2481) & VN_data_in(2481);
  VN413_in4 <= VN_sign_in(2482) & VN_data_in(2482);
  VN413_in5 <= VN_sign_in(2483) & VN_data_in(2483);
  VN414_in0 <= VN_sign_in(2484) & VN_data_in(2484);
  VN414_in1 <= VN_sign_in(2485) & VN_data_in(2485);
  VN414_in2 <= VN_sign_in(2486) & VN_data_in(2486);
  VN414_in3 <= VN_sign_in(2487) & VN_data_in(2487);
  VN414_in4 <= VN_sign_in(2488) & VN_data_in(2488);
  VN414_in5 <= VN_sign_in(2489) & VN_data_in(2489);
  VN415_in0 <= VN_sign_in(2490) & VN_data_in(2490);
  VN415_in1 <= VN_sign_in(2491) & VN_data_in(2491);
  VN415_in2 <= VN_sign_in(2492) & VN_data_in(2492);
  VN415_in3 <= VN_sign_in(2493) & VN_data_in(2493);
  VN415_in4 <= VN_sign_in(2494) & VN_data_in(2494);
  VN415_in5 <= VN_sign_in(2495) & VN_data_in(2495);
  VN416_in0 <= VN_sign_in(2496) & VN_data_in(2496);
  VN416_in1 <= VN_sign_in(2497) & VN_data_in(2497);
  VN416_in2 <= VN_sign_in(2498) & VN_data_in(2498);
  VN416_in3 <= VN_sign_in(2499) & VN_data_in(2499);
  VN416_in4 <= VN_sign_in(2500) & VN_data_in(2500);
  VN416_in5 <= VN_sign_in(2501) & VN_data_in(2501);
  VN417_in0 <= VN_sign_in(2502) & VN_data_in(2502);
  VN417_in1 <= VN_sign_in(2503) & VN_data_in(2503);
  VN417_in2 <= VN_sign_in(2504) & VN_data_in(2504);
  VN417_in3 <= VN_sign_in(2505) & VN_data_in(2505);
  VN417_in4 <= VN_sign_in(2506) & VN_data_in(2506);
  VN417_in5 <= VN_sign_in(2507) & VN_data_in(2507);
  VN418_in0 <= VN_sign_in(2508) & VN_data_in(2508);
  VN418_in1 <= VN_sign_in(2509) & VN_data_in(2509);
  VN418_in2 <= VN_sign_in(2510) & VN_data_in(2510);
  VN418_in3 <= VN_sign_in(2511) & VN_data_in(2511);
  VN418_in4 <= VN_sign_in(2512) & VN_data_in(2512);
  VN418_in5 <= VN_sign_in(2513) & VN_data_in(2513);
  VN419_in0 <= VN_sign_in(2514) & VN_data_in(2514);
  VN419_in1 <= VN_sign_in(2515) & VN_data_in(2515);
  VN419_in2 <= VN_sign_in(2516) & VN_data_in(2516);
  VN419_in3 <= VN_sign_in(2517) & VN_data_in(2517);
  VN419_in4 <= VN_sign_in(2518) & VN_data_in(2518);
  VN419_in5 <= VN_sign_in(2519) & VN_data_in(2519);
  VN420_in0 <= VN_sign_in(2520) & VN_data_in(2520);
  VN420_in1 <= VN_sign_in(2521) & VN_data_in(2521);
  VN420_in2 <= VN_sign_in(2522) & VN_data_in(2522);
  VN420_in3 <= VN_sign_in(2523) & VN_data_in(2523);
  VN420_in4 <= VN_sign_in(2524) & VN_data_in(2524);
  VN420_in5 <= VN_sign_in(2525) & VN_data_in(2525);
  VN421_in0 <= VN_sign_in(2526) & VN_data_in(2526);
  VN421_in1 <= VN_sign_in(2527) & VN_data_in(2527);
  VN421_in2 <= VN_sign_in(2528) & VN_data_in(2528);
  VN421_in3 <= VN_sign_in(2529) & VN_data_in(2529);
  VN421_in4 <= VN_sign_in(2530) & VN_data_in(2530);
  VN421_in5 <= VN_sign_in(2531) & VN_data_in(2531);
  VN422_in0 <= VN_sign_in(2532) & VN_data_in(2532);
  VN422_in1 <= VN_sign_in(2533) & VN_data_in(2533);
  VN422_in2 <= VN_sign_in(2534) & VN_data_in(2534);
  VN422_in3 <= VN_sign_in(2535) & VN_data_in(2535);
  VN422_in4 <= VN_sign_in(2536) & VN_data_in(2536);
  VN422_in5 <= VN_sign_in(2537) & VN_data_in(2537);
  VN423_in0 <= VN_sign_in(2538) & VN_data_in(2538);
  VN423_in1 <= VN_sign_in(2539) & VN_data_in(2539);
  VN423_in2 <= VN_sign_in(2540) & VN_data_in(2540);
  VN423_in3 <= VN_sign_in(2541) & VN_data_in(2541);
  VN423_in4 <= VN_sign_in(2542) & VN_data_in(2542);
  VN423_in5 <= VN_sign_in(2543) & VN_data_in(2543);
  VN424_in0 <= VN_sign_in(2544) & VN_data_in(2544);
  VN424_in1 <= VN_sign_in(2545) & VN_data_in(2545);
  VN424_in2 <= VN_sign_in(2546) & VN_data_in(2546);
  VN424_in3 <= VN_sign_in(2547) & VN_data_in(2547);
  VN424_in4 <= VN_sign_in(2548) & VN_data_in(2548);
  VN424_in5 <= VN_sign_in(2549) & VN_data_in(2549);
  VN425_in0 <= VN_sign_in(2550) & VN_data_in(2550);
  VN425_in1 <= VN_sign_in(2551) & VN_data_in(2551);
  VN425_in2 <= VN_sign_in(2552) & VN_data_in(2552);
  VN425_in3 <= VN_sign_in(2553) & VN_data_in(2553);
  VN425_in4 <= VN_sign_in(2554) & VN_data_in(2554);
  VN425_in5 <= VN_sign_in(2555) & VN_data_in(2555);
  VN426_in0 <= VN_sign_in(2556) & VN_data_in(2556);
  VN426_in1 <= VN_sign_in(2557) & VN_data_in(2557);
  VN426_in2 <= VN_sign_in(2558) & VN_data_in(2558);
  VN426_in3 <= VN_sign_in(2559) & VN_data_in(2559);
  VN426_in4 <= VN_sign_in(2560) & VN_data_in(2560);
  VN426_in5 <= VN_sign_in(2561) & VN_data_in(2561);
  VN427_in0 <= VN_sign_in(2562) & VN_data_in(2562);
  VN427_in1 <= VN_sign_in(2563) & VN_data_in(2563);
  VN427_in2 <= VN_sign_in(2564) & VN_data_in(2564);
  VN427_in3 <= VN_sign_in(2565) & VN_data_in(2565);
  VN427_in4 <= VN_sign_in(2566) & VN_data_in(2566);
  VN427_in5 <= VN_sign_in(2567) & VN_data_in(2567);
  VN428_in0 <= VN_sign_in(2568) & VN_data_in(2568);
  VN428_in1 <= VN_sign_in(2569) & VN_data_in(2569);
  VN428_in2 <= VN_sign_in(2570) & VN_data_in(2570);
  VN428_in3 <= VN_sign_in(2571) & VN_data_in(2571);
  VN428_in4 <= VN_sign_in(2572) & VN_data_in(2572);
  VN428_in5 <= VN_sign_in(2573) & VN_data_in(2573);
  VN429_in0 <= VN_sign_in(2574) & VN_data_in(2574);
  VN429_in1 <= VN_sign_in(2575) & VN_data_in(2575);
  VN429_in2 <= VN_sign_in(2576) & VN_data_in(2576);
  VN429_in3 <= VN_sign_in(2577) & VN_data_in(2577);
  VN429_in4 <= VN_sign_in(2578) & VN_data_in(2578);
  VN429_in5 <= VN_sign_in(2579) & VN_data_in(2579);
  VN430_in0 <= VN_sign_in(2580) & VN_data_in(2580);
  VN430_in1 <= VN_sign_in(2581) & VN_data_in(2581);
  VN430_in2 <= VN_sign_in(2582) & VN_data_in(2582);
  VN430_in3 <= VN_sign_in(2583) & VN_data_in(2583);
  VN430_in4 <= VN_sign_in(2584) & VN_data_in(2584);
  VN430_in5 <= VN_sign_in(2585) & VN_data_in(2585);
  VN431_in0 <= VN_sign_in(2586) & VN_data_in(2586);
  VN431_in1 <= VN_sign_in(2587) & VN_data_in(2587);
  VN431_in2 <= VN_sign_in(2588) & VN_data_in(2588);
  VN431_in3 <= VN_sign_in(2589) & VN_data_in(2589);
  VN431_in4 <= VN_sign_in(2590) & VN_data_in(2590);
  VN431_in5 <= VN_sign_in(2591) & VN_data_in(2591);
  VN432_in0 <= VN_sign_in(2592) & VN_data_in(2592);
  VN432_in1 <= VN_sign_in(2593) & VN_data_in(2593);
  VN432_in2 <= VN_sign_in(2594) & VN_data_in(2594);
  VN432_in3 <= VN_sign_in(2595) & VN_data_in(2595);
  VN432_in4 <= VN_sign_in(2596) & VN_data_in(2596);
  VN432_in5 <= VN_sign_in(2597) & VN_data_in(2597);
  VN433_in0 <= VN_sign_in(2598) & VN_data_in(2598);
  VN433_in1 <= VN_sign_in(2599) & VN_data_in(2599);
  VN433_in2 <= VN_sign_in(2600) & VN_data_in(2600);
  VN433_in3 <= VN_sign_in(2601) & VN_data_in(2601);
  VN433_in4 <= VN_sign_in(2602) & VN_data_in(2602);
  VN433_in5 <= VN_sign_in(2603) & VN_data_in(2603);
  VN434_in0 <= VN_sign_in(2604) & VN_data_in(2604);
  VN434_in1 <= VN_sign_in(2605) & VN_data_in(2605);
  VN434_in2 <= VN_sign_in(2606) & VN_data_in(2606);
  VN434_in3 <= VN_sign_in(2607) & VN_data_in(2607);
  VN434_in4 <= VN_sign_in(2608) & VN_data_in(2608);
  VN434_in5 <= VN_sign_in(2609) & VN_data_in(2609);
  VN435_in0 <= VN_sign_in(2610) & VN_data_in(2610);
  VN435_in1 <= VN_sign_in(2611) & VN_data_in(2611);
  VN435_in2 <= VN_sign_in(2612) & VN_data_in(2612);
  VN435_in3 <= VN_sign_in(2613) & VN_data_in(2613);
  VN435_in4 <= VN_sign_in(2614) & VN_data_in(2614);
  VN435_in5 <= VN_sign_in(2615) & VN_data_in(2615);
  VN436_in0 <= VN_sign_in(2616) & VN_data_in(2616);
  VN436_in1 <= VN_sign_in(2617) & VN_data_in(2617);
  VN436_in2 <= VN_sign_in(2618) & VN_data_in(2618);
  VN436_in3 <= VN_sign_in(2619) & VN_data_in(2619);
  VN436_in4 <= VN_sign_in(2620) & VN_data_in(2620);
  VN436_in5 <= VN_sign_in(2621) & VN_data_in(2621);
  VN437_in0 <= VN_sign_in(2622) & VN_data_in(2622);
  VN437_in1 <= VN_sign_in(2623) & VN_data_in(2623);
  VN437_in2 <= VN_sign_in(2624) & VN_data_in(2624);
  VN437_in3 <= VN_sign_in(2625) & VN_data_in(2625);
  VN437_in4 <= VN_sign_in(2626) & VN_data_in(2626);
  VN437_in5 <= VN_sign_in(2627) & VN_data_in(2627);
  VN438_in0 <= VN_sign_in(2628) & VN_data_in(2628);
  VN438_in1 <= VN_sign_in(2629) & VN_data_in(2629);
  VN438_in2 <= VN_sign_in(2630) & VN_data_in(2630);
  VN438_in3 <= VN_sign_in(2631) & VN_data_in(2631);
  VN438_in4 <= VN_sign_in(2632) & VN_data_in(2632);
  VN438_in5 <= VN_sign_in(2633) & VN_data_in(2633);
  VN439_in0 <= VN_sign_in(2634) & VN_data_in(2634);
  VN439_in1 <= VN_sign_in(2635) & VN_data_in(2635);
  VN439_in2 <= VN_sign_in(2636) & VN_data_in(2636);
  VN439_in3 <= VN_sign_in(2637) & VN_data_in(2637);
  VN439_in4 <= VN_sign_in(2638) & VN_data_in(2638);
  VN439_in5 <= VN_sign_in(2639) & VN_data_in(2639);
  VN440_in0 <= VN_sign_in(2640) & VN_data_in(2640);
  VN440_in1 <= VN_sign_in(2641) & VN_data_in(2641);
  VN440_in2 <= VN_sign_in(2642) & VN_data_in(2642);
  VN440_in3 <= VN_sign_in(2643) & VN_data_in(2643);
  VN440_in4 <= VN_sign_in(2644) & VN_data_in(2644);
  VN440_in5 <= VN_sign_in(2645) & VN_data_in(2645);
  VN441_in0 <= VN_sign_in(2646) & VN_data_in(2646);
  VN441_in1 <= VN_sign_in(2647) & VN_data_in(2647);
  VN441_in2 <= VN_sign_in(2648) & VN_data_in(2648);
  VN441_in3 <= VN_sign_in(2649) & VN_data_in(2649);
  VN441_in4 <= VN_sign_in(2650) & VN_data_in(2650);
  VN441_in5 <= VN_sign_in(2651) & VN_data_in(2651);
  VN442_in0 <= VN_sign_in(2652) & VN_data_in(2652);
  VN442_in1 <= VN_sign_in(2653) & VN_data_in(2653);
  VN442_in2 <= VN_sign_in(2654) & VN_data_in(2654);
  VN442_in3 <= VN_sign_in(2655) & VN_data_in(2655);
  VN442_in4 <= VN_sign_in(2656) & VN_data_in(2656);
  VN442_in5 <= VN_sign_in(2657) & VN_data_in(2657);
  VN443_in0 <= VN_sign_in(2658) & VN_data_in(2658);
  VN443_in1 <= VN_sign_in(2659) & VN_data_in(2659);
  VN443_in2 <= VN_sign_in(2660) & VN_data_in(2660);
  VN443_in3 <= VN_sign_in(2661) & VN_data_in(2661);
  VN443_in4 <= VN_sign_in(2662) & VN_data_in(2662);
  VN443_in5 <= VN_sign_in(2663) & VN_data_in(2663);
  VN444_in0 <= VN_sign_in(2664) & VN_data_in(2664);
  VN444_in1 <= VN_sign_in(2665) & VN_data_in(2665);
  VN444_in2 <= VN_sign_in(2666) & VN_data_in(2666);
  VN444_in3 <= VN_sign_in(2667) & VN_data_in(2667);
  VN444_in4 <= VN_sign_in(2668) & VN_data_in(2668);
  VN444_in5 <= VN_sign_in(2669) & VN_data_in(2669);
  VN445_in0 <= VN_sign_in(2670) & VN_data_in(2670);
  VN445_in1 <= VN_sign_in(2671) & VN_data_in(2671);
  VN445_in2 <= VN_sign_in(2672) & VN_data_in(2672);
  VN445_in3 <= VN_sign_in(2673) & VN_data_in(2673);
  VN445_in4 <= VN_sign_in(2674) & VN_data_in(2674);
  VN445_in5 <= VN_sign_in(2675) & VN_data_in(2675);
  VN446_in0 <= VN_sign_in(2676) & VN_data_in(2676);
  VN446_in1 <= VN_sign_in(2677) & VN_data_in(2677);
  VN446_in2 <= VN_sign_in(2678) & VN_data_in(2678);
  VN446_in3 <= VN_sign_in(2679) & VN_data_in(2679);
  VN446_in4 <= VN_sign_in(2680) & VN_data_in(2680);
  VN446_in5 <= VN_sign_in(2681) & VN_data_in(2681);
  VN447_in0 <= VN_sign_in(2682) & VN_data_in(2682);
  VN447_in1 <= VN_sign_in(2683) & VN_data_in(2683);
  VN447_in2 <= VN_sign_in(2684) & VN_data_in(2684);
  VN447_in3 <= VN_sign_in(2685) & VN_data_in(2685);
  VN447_in4 <= VN_sign_in(2686) & VN_data_in(2686);
  VN447_in5 <= VN_sign_in(2687) & VN_data_in(2687);
  VN448_in0 <= VN_sign_in(2688) & VN_data_in(2688);
  VN448_in1 <= VN_sign_in(2689) & VN_data_in(2689);
  VN448_in2 <= VN_sign_in(2690) & VN_data_in(2690);
  VN448_in3 <= VN_sign_in(2691) & VN_data_in(2691);
  VN448_in4 <= VN_sign_in(2692) & VN_data_in(2692);
  VN448_in5 <= VN_sign_in(2693) & VN_data_in(2693);
  VN449_in0 <= VN_sign_in(2694) & VN_data_in(2694);
  VN449_in1 <= VN_sign_in(2695) & VN_data_in(2695);
  VN449_in2 <= VN_sign_in(2696) & VN_data_in(2696);
  VN449_in3 <= VN_sign_in(2697) & VN_data_in(2697);
  VN449_in4 <= VN_sign_in(2698) & VN_data_in(2698);
  VN449_in5 <= VN_sign_in(2699) & VN_data_in(2699);
  VN450_in0 <= VN_sign_in(2700) & VN_data_in(2700);
  VN450_in1 <= VN_sign_in(2701) & VN_data_in(2701);
  VN450_in2 <= VN_sign_in(2702) & VN_data_in(2702);
  VN450_in3 <= VN_sign_in(2703) & VN_data_in(2703);
  VN450_in4 <= VN_sign_in(2704) & VN_data_in(2704);
  VN450_in5 <= VN_sign_in(2705) & VN_data_in(2705);
  VN451_in0 <= VN_sign_in(2706) & VN_data_in(2706);
  VN451_in1 <= VN_sign_in(2707) & VN_data_in(2707);
  VN451_in2 <= VN_sign_in(2708) & VN_data_in(2708);
  VN451_in3 <= VN_sign_in(2709) & VN_data_in(2709);
  VN451_in4 <= VN_sign_in(2710) & VN_data_in(2710);
  VN451_in5 <= VN_sign_in(2711) & VN_data_in(2711);
  VN452_in0 <= VN_sign_in(2712) & VN_data_in(2712);
  VN452_in1 <= VN_sign_in(2713) & VN_data_in(2713);
  VN452_in2 <= VN_sign_in(2714) & VN_data_in(2714);
  VN452_in3 <= VN_sign_in(2715) & VN_data_in(2715);
  VN452_in4 <= VN_sign_in(2716) & VN_data_in(2716);
  VN452_in5 <= VN_sign_in(2717) & VN_data_in(2717);
  VN453_in0 <= VN_sign_in(2718) & VN_data_in(2718);
  VN453_in1 <= VN_sign_in(2719) & VN_data_in(2719);
  VN453_in2 <= VN_sign_in(2720) & VN_data_in(2720);
  VN453_in3 <= VN_sign_in(2721) & VN_data_in(2721);
  VN453_in4 <= VN_sign_in(2722) & VN_data_in(2722);
  VN453_in5 <= VN_sign_in(2723) & VN_data_in(2723);
  VN454_in0 <= VN_sign_in(2724) & VN_data_in(2724);
  VN454_in1 <= VN_sign_in(2725) & VN_data_in(2725);
  VN454_in2 <= VN_sign_in(2726) & VN_data_in(2726);
  VN454_in3 <= VN_sign_in(2727) & VN_data_in(2727);
  VN454_in4 <= VN_sign_in(2728) & VN_data_in(2728);
  VN454_in5 <= VN_sign_in(2729) & VN_data_in(2729);
  VN455_in0 <= VN_sign_in(2730) & VN_data_in(2730);
  VN455_in1 <= VN_sign_in(2731) & VN_data_in(2731);
  VN455_in2 <= VN_sign_in(2732) & VN_data_in(2732);
  VN455_in3 <= VN_sign_in(2733) & VN_data_in(2733);
  VN455_in4 <= VN_sign_in(2734) & VN_data_in(2734);
  VN455_in5 <= VN_sign_in(2735) & VN_data_in(2735);
  VN456_in0 <= VN_sign_in(2736) & VN_data_in(2736);
  VN456_in1 <= VN_sign_in(2737) & VN_data_in(2737);
  VN456_in2 <= VN_sign_in(2738) & VN_data_in(2738);
  VN456_in3 <= VN_sign_in(2739) & VN_data_in(2739);
  VN456_in4 <= VN_sign_in(2740) & VN_data_in(2740);
  VN456_in5 <= VN_sign_in(2741) & VN_data_in(2741);
  VN457_in0 <= VN_sign_in(2742) & VN_data_in(2742);
  VN457_in1 <= VN_sign_in(2743) & VN_data_in(2743);
  VN457_in2 <= VN_sign_in(2744) & VN_data_in(2744);
  VN457_in3 <= VN_sign_in(2745) & VN_data_in(2745);
  VN457_in4 <= VN_sign_in(2746) & VN_data_in(2746);
  VN457_in5 <= VN_sign_in(2747) & VN_data_in(2747);
  VN458_in0 <= VN_sign_in(2748) & VN_data_in(2748);
  VN458_in1 <= VN_sign_in(2749) & VN_data_in(2749);
  VN458_in2 <= VN_sign_in(2750) & VN_data_in(2750);
  VN458_in3 <= VN_sign_in(2751) & VN_data_in(2751);
  VN458_in4 <= VN_sign_in(2752) & VN_data_in(2752);
  VN458_in5 <= VN_sign_in(2753) & VN_data_in(2753);
  VN459_in0 <= VN_sign_in(2754) & VN_data_in(2754);
  VN459_in1 <= VN_sign_in(2755) & VN_data_in(2755);
  VN459_in2 <= VN_sign_in(2756) & VN_data_in(2756);
  VN459_in3 <= VN_sign_in(2757) & VN_data_in(2757);
  VN459_in4 <= VN_sign_in(2758) & VN_data_in(2758);
  VN459_in5 <= VN_sign_in(2759) & VN_data_in(2759);
  VN460_in0 <= VN_sign_in(2760) & VN_data_in(2760);
  VN460_in1 <= VN_sign_in(2761) & VN_data_in(2761);
  VN460_in2 <= VN_sign_in(2762) & VN_data_in(2762);
  VN460_in3 <= VN_sign_in(2763) & VN_data_in(2763);
  VN460_in4 <= VN_sign_in(2764) & VN_data_in(2764);
  VN460_in5 <= VN_sign_in(2765) & VN_data_in(2765);
  VN461_in0 <= VN_sign_in(2766) & VN_data_in(2766);
  VN461_in1 <= VN_sign_in(2767) & VN_data_in(2767);
  VN461_in2 <= VN_sign_in(2768) & VN_data_in(2768);
  VN461_in3 <= VN_sign_in(2769) & VN_data_in(2769);
  VN461_in4 <= VN_sign_in(2770) & VN_data_in(2770);
  VN461_in5 <= VN_sign_in(2771) & VN_data_in(2771);
  VN462_in0 <= VN_sign_in(2772) & VN_data_in(2772);
  VN462_in1 <= VN_sign_in(2773) & VN_data_in(2773);
  VN462_in2 <= VN_sign_in(2774) & VN_data_in(2774);
  VN462_in3 <= VN_sign_in(2775) & VN_data_in(2775);
  VN462_in4 <= VN_sign_in(2776) & VN_data_in(2776);
  VN462_in5 <= VN_sign_in(2777) & VN_data_in(2777);
  VN463_in0 <= VN_sign_in(2778) & VN_data_in(2778);
  VN463_in1 <= VN_sign_in(2779) & VN_data_in(2779);
  VN463_in2 <= VN_sign_in(2780) & VN_data_in(2780);
  VN463_in3 <= VN_sign_in(2781) & VN_data_in(2781);
  VN463_in4 <= VN_sign_in(2782) & VN_data_in(2782);
  VN463_in5 <= VN_sign_in(2783) & VN_data_in(2783);
  VN464_in0 <= VN_sign_in(2784) & VN_data_in(2784);
  VN464_in1 <= VN_sign_in(2785) & VN_data_in(2785);
  VN464_in2 <= VN_sign_in(2786) & VN_data_in(2786);
  VN464_in3 <= VN_sign_in(2787) & VN_data_in(2787);
  VN464_in4 <= VN_sign_in(2788) & VN_data_in(2788);
  VN464_in5 <= VN_sign_in(2789) & VN_data_in(2789);
  VN465_in0 <= VN_sign_in(2790) & VN_data_in(2790);
  VN465_in1 <= VN_sign_in(2791) & VN_data_in(2791);
  VN465_in2 <= VN_sign_in(2792) & VN_data_in(2792);
  VN465_in3 <= VN_sign_in(2793) & VN_data_in(2793);
  VN465_in4 <= VN_sign_in(2794) & VN_data_in(2794);
  VN465_in5 <= VN_sign_in(2795) & VN_data_in(2795);
  VN466_in0 <= VN_sign_in(2796) & VN_data_in(2796);
  VN466_in1 <= VN_sign_in(2797) & VN_data_in(2797);
  VN466_in2 <= VN_sign_in(2798) & VN_data_in(2798);
  VN466_in3 <= VN_sign_in(2799) & VN_data_in(2799);
  VN466_in4 <= VN_sign_in(2800) & VN_data_in(2800);
  VN466_in5 <= VN_sign_in(2801) & VN_data_in(2801);
  VN467_in0 <= VN_sign_in(2802) & VN_data_in(2802);
  VN467_in1 <= VN_sign_in(2803) & VN_data_in(2803);
  VN467_in2 <= VN_sign_in(2804) & VN_data_in(2804);
  VN467_in3 <= VN_sign_in(2805) & VN_data_in(2805);
  VN467_in4 <= VN_sign_in(2806) & VN_data_in(2806);
  VN467_in5 <= VN_sign_in(2807) & VN_data_in(2807);
  VN468_in0 <= VN_sign_in(2808) & VN_data_in(2808);
  VN468_in1 <= VN_sign_in(2809) & VN_data_in(2809);
  VN468_in2 <= VN_sign_in(2810) & VN_data_in(2810);
  VN468_in3 <= VN_sign_in(2811) & VN_data_in(2811);
  VN468_in4 <= VN_sign_in(2812) & VN_data_in(2812);
  VN468_in5 <= VN_sign_in(2813) & VN_data_in(2813);
  VN469_in0 <= VN_sign_in(2814) & VN_data_in(2814);
  VN469_in1 <= VN_sign_in(2815) & VN_data_in(2815);
  VN469_in2 <= VN_sign_in(2816) & VN_data_in(2816);
  VN469_in3 <= VN_sign_in(2817) & VN_data_in(2817);
  VN469_in4 <= VN_sign_in(2818) & VN_data_in(2818);
  VN469_in5 <= VN_sign_in(2819) & VN_data_in(2819);
  VN470_in0 <= VN_sign_in(2820) & VN_data_in(2820);
  VN470_in1 <= VN_sign_in(2821) & VN_data_in(2821);
  VN470_in2 <= VN_sign_in(2822) & VN_data_in(2822);
  VN470_in3 <= VN_sign_in(2823) & VN_data_in(2823);
  VN470_in4 <= VN_sign_in(2824) & VN_data_in(2824);
  VN470_in5 <= VN_sign_in(2825) & VN_data_in(2825);
  VN471_in0 <= VN_sign_in(2826) & VN_data_in(2826);
  VN471_in1 <= VN_sign_in(2827) & VN_data_in(2827);
  VN471_in2 <= VN_sign_in(2828) & VN_data_in(2828);
  VN471_in3 <= VN_sign_in(2829) & VN_data_in(2829);
  VN471_in4 <= VN_sign_in(2830) & VN_data_in(2830);
  VN471_in5 <= VN_sign_in(2831) & VN_data_in(2831);
  VN472_in0 <= VN_sign_in(2832) & VN_data_in(2832);
  VN472_in1 <= VN_sign_in(2833) & VN_data_in(2833);
  VN472_in2 <= VN_sign_in(2834) & VN_data_in(2834);
  VN472_in3 <= VN_sign_in(2835) & VN_data_in(2835);
  VN472_in4 <= VN_sign_in(2836) & VN_data_in(2836);
  VN472_in5 <= VN_sign_in(2837) & VN_data_in(2837);
  VN473_in0 <= VN_sign_in(2838) & VN_data_in(2838);
  VN473_in1 <= VN_sign_in(2839) & VN_data_in(2839);
  VN473_in2 <= VN_sign_in(2840) & VN_data_in(2840);
  VN473_in3 <= VN_sign_in(2841) & VN_data_in(2841);
  VN473_in4 <= VN_sign_in(2842) & VN_data_in(2842);
  VN473_in5 <= VN_sign_in(2843) & VN_data_in(2843);
  VN474_in0 <= VN_sign_in(2844) & VN_data_in(2844);
  VN474_in1 <= VN_sign_in(2845) & VN_data_in(2845);
  VN474_in2 <= VN_sign_in(2846) & VN_data_in(2846);
  VN474_in3 <= VN_sign_in(2847) & VN_data_in(2847);
  VN474_in4 <= VN_sign_in(2848) & VN_data_in(2848);
  VN474_in5 <= VN_sign_in(2849) & VN_data_in(2849);
  VN475_in0 <= VN_sign_in(2850) & VN_data_in(2850);
  VN475_in1 <= VN_sign_in(2851) & VN_data_in(2851);
  VN475_in2 <= VN_sign_in(2852) & VN_data_in(2852);
  VN475_in3 <= VN_sign_in(2853) & VN_data_in(2853);
  VN475_in4 <= VN_sign_in(2854) & VN_data_in(2854);
  VN475_in5 <= VN_sign_in(2855) & VN_data_in(2855);
  VN476_in0 <= VN_sign_in(2856) & VN_data_in(2856);
  VN476_in1 <= VN_sign_in(2857) & VN_data_in(2857);
  VN476_in2 <= VN_sign_in(2858) & VN_data_in(2858);
  VN476_in3 <= VN_sign_in(2859) & VN_data_in(2859);
  VN476_in4 <= VN_sign_in(2860) & VN_data_in(2860);
  VN476_in5 <= VN_sign_in(2861) & VN_data_in(2861);
  VN477_in0 <= VN_sign_in(2862) & VN_data_in(2862);
  VN477_in1 <= VN_sign_in(2863) & VN_data_in(2863);
  VN477_in2 <= VN_sign_in(2864) & VN_data_in(2864);
  VN477_in3 <= VN_sign_in(2865) & VN_data_in(2865);
  VN477_in4 <= VN_sign_in(2866) & VN_data_in(2866);
  VN477_in5 <= VN_sign_in(2867) & VN_data_in(2867);
  VN478_in0 <= VN_sign_in(2868) & VN_data_in(2868);
  VN478_in1 <= VN_sign_in(2869) & VN_data_in(2869);
  VN478_in2 <= VN_sign_in(2870) & VN_data_in(2870);
  VN478_in3 <= VN_sign_in(2871) & VN_data_in(2871);
  VN478_in4 <= VN_sign_in(2872) & VN_data_in(2872);
  VN478_in5 <= VN_sign_in(2873) & VN_data_in(2873);
  VN479_in0 <= VN_sign_in(2874) & VN_data_in(2874);
  VN479_in1 <= VN_sign_in(2875) & VN_data_in(2875);
  VN479_in2 <= VN_sign_in(2876) & VN_data_in(2876);
  VN479_in3 <= VN_sign_in(2877) & VN_data_in(2877);
  VN479_in4 <= VN_sign_in(2878) & VN_data_in(2878);
  VN479_in5 <= VN_sign_in(2879) & VN_data_in(2879);
  VN480_in0 <= VN_sign_in(2880) & VN_data_in(2880);
  VN480_in1 <= VN_sign_in(2881) & VN_data_in(2881);
  VN480_in2 <= VN_sign_in(2882) & VN_data_in(2882);
  VN480_in3 <= VN_sign_in(2883) & VN_data_in(2883);
  VN480_in4 <= VN_sign_in(2884) & VN_data_in(2884);
  VN480_in5 <= VN_sign_in(2885) & VN_data_in(2885);
  VN481_in0 <= VN_sign_in(2886) & VN_data_in(2886);
  VN481_in1 <= VN_sign_in(2887) & VN_data_in(2887);
  VN481_in2 <= VN_sign_in(2888) & VN_data_in(2888);
  VN481_in3 <= VN_sign_in(2889) & VN_data_in(2889);
  VN481_in4 <= VN_sign_in(2890) & VN_data_in(2890);
  VN481_in5 <= VN_sign_in(2891) & VN_data_in(2891);
  VN482_in0 <= VN_sign_in(2892) & VN_data_in(2892);
  VN482_in1 <= VN_sign_in(2893) & VN_data_in(2893);
  VN482_in2 <= VN_sign_in(2894) & VN_data_in(2894);
  VN482_in3 <= VN_sign_in(2895) & VN_data_in(2895);
  VN482_in4 <= VN_sign_in(2896) & VN_data_in(2896);
  VN482_in5 <= VN_sign_in(2897) & VN_data_in(2897);
  VN483_in0 <= VN_sign_in(2898) & VN_data_in(2898);
  VN483_in1 <= VN_sign_in(2899) & VN_data_in(2899);
  VN483_in2 <= VN_sign_in(2900) & VN_data_in(2900);
  VN483_in3 <= VN_sign_in(2901) & VN_data_in(2901);
  VN483_in4 <= VN_sign_in(2902) & VN_data_in(2902);
  VN483_in5 <= VN_sign_in(2903) & VN_data_in(2903);
  VN484_in0 <= VN_sign_in(2904) & VN_data_in(2904);
  VN484_in1 <= VN_sign_in(2905) & VN_data_in(2905);
  VN484_in2 <= VN_sign_in(2906) & VN_data_in(2906);
  VN484_in3 <= VN_sign_in(2907) & VN_data_in(2907);
  VN484_in4 <= VN_sign_in(2908) & VN_data_in(2908);
  VN484_in5 <= VN_sign_in(2909) & VN_data_in(2909);
  VN485_in0 <= VN_sign_in(2910) & VN_data_in(2910);
  VN485_in1 <= VN_sign_in(2911) & VN_data_in(2911);
  VN485_in2 <= VN_sign_in(2912) & VN_data_in(2912);
  VN485_in3 <= VN_sign_in(2913) & VN_data_in(2913);
  VN485_in4 <= VN_sign_in(2914) & VN_data_in(2914);
  VN485_in5 <= VN_sign_in(2915) & VN_data_in(2915);
  VN486_in0 <= VN_sign_in(2916) & VN_data_in(2916);
  VN486_in1 <= VN_sign_in(2917) & VN_data_in(2917);
  VN486_in2 <= VN_sign_in(2918) & VN_data_in(2918);
  VN486_in3 <= VN_sign_in(2919) & VN_data_in(2919);
  VN486_in4 <= VN_sign_in(2920) & VN_data_in(2920);
  VN486_in5 <= VN_sign_in(2921) & VN_data_in(2921);
  VN487_in0 <= VN_sign_in(2922) & VN_data_in(2922);
  VN487_in1 <= VN_sign_in(2923) & VN_data_in(2923);
  VN487_in2 <= VN_sign_in(2924) & VN_data_in(2924);
  VN487_in3 <= VN_sign_in(2925) & VN_data_in(2925);
  VN487_in4 <= VN_sign_in(2926) & VN_data_in(2926);
  VN487_in5 <= VN_sign_in(2927) & VN_data_in(2927);
  VN488_in0 <= VN_sign_in(2928) & VN_data_in(2928);
  VN488_in1 <= VN_sign_in(2929) & VN_data_in(2929);
  VN488_in2 <= VN_sign_in(2930) & VN_data_in(2930);
  VN488_in3 <= VN_sign_in(2931) & VN_data_in(2931);
  VN488_in4 <= VN_sign_in(2932) & VN_data_in(2932);
  VN488_in5 <= VN_sign_in(2933) & VN_data_in(2933);
  VN489_in0 <= VN_sign_in(2934) & VN_data_in(2934);
  VN489_in1 <= VN_sign_in(2935) & VN_data_in(2935);
  VN489_in2 <= VN_sign_in(2936) & VN_data_in(2936);
  VN489_in3 <= VN_sign_in(2937) & VN_data_in(2937);
  VN489_in4 <= VN_sign_in(2938) & VN_data_in(2938);
  VN489_in5 <= VN_sign_in(2939) & VN_data_in(2939);
  VN490_in0 <= VN_sign_in(2940) & VN_data_in(2940);
  VN490_in1 <= VN_sign_in(2941) & VN_data_in(2941);
  VN490_in2 <= VN_sign_in(2942) & VN_data_in(2942);
  VN490_in3 <= VN_sign_in(2943) & VN_data_in(2943);
  VN490_in4 <= VN_sign_in(2944) & VN_data_in(2944);
  VN490_in5 <= VN_sign_in(2945) & VN_data_in(2945);
  VN491_in0 <= VN_sign_in(2946) & VN_data_in(2946);
  VN491_in1 <= VN_sign_in(2947) & VN_data_in(2947);
  VN491_in2 <= VN_sign_in(2948) & VN_data_in(2948);
  VN491_in3 <= VN_sign_in(2949) & VN_data_in(2949);
  VN491_in4 <= VN_sign_in(2950) & VN_data_in(2950);
  VN491_in5 <= VN_sign_in(2951) & VN_data_in(2951);
  VN492_in0 <= VN_sign_in(2952) & VN_data_in(2952);
  VN492_in1 <= VN_sign_in(2953) & VN_data_in(2953);
  VN492_in2 <= VN_sign_in(2954) & VN_data_in(2954);
  VN492_in3 <= VN_sign_in(2955) & VN_data_in(2955);
  VN492_in4 <= VN_sign_in(2956) & VN_data_in(2956);
  VN492_in5 <= VN_sign_in(2957) & VN_data_in(2957);
  VN493_in0 <= VN_sign_in(2958) & VN_data_in(2958);
  VN493_in1 <= VN_sign_in(2959) & VN_data_in(2959);
  VN493_in2 <= VN_sign_in(2960) & VN_data_in(2960);
  VN493_in3 <= VN_sign_in(2961) & VN_data_in(2961);
  VN493_in4 <= VN_sign_in(2962) & VN_data_in(2962);
  VN493_in5 <= VN_sign_in(2963) & VN_data_in(2963);
  VN494_in0 <= VN_sign_in(2964) & VN_data_in(2964);
  VN494_in1 <= VN_sign_in(2965) & VN_data_in(2965);
  VN494_in2 <= VN_sign_in(2966) & VN_data_in(2966);
  VN494_in3 <= VN_sign_in(2967) & VN_data_in(2967);
  VN494_in4 <= VN_sign_in(2968) & VN_data_in(2968);
  VN494_in5 <= VN_sign_in(2969) & VN_data_in(2969);
  VN495_in0 <= VN_sign_in(2970) & VN_data_in(2970);
  VN495_in1 <= VN_sign_in(2971) & VN_data_in(2971);
  VN495_in2 <= VN_sign_in(2972) & VN_data_in(2972);
  VN495_in3 <= VN_sign_in(2973) & VN_data_in(2973);
  VN495_in4 <= VN_sign_in(2974) & VN_data_in(2974);
  VN495_in5 <= VN_sign_in(2975) & VN_data_in(2975);
  VN496_in0 <= VN_sign_in(2976) & VN_data_in(2976);
  VN496_in1 <= VN_sign_in(2977) & VN_data_in(2977);
  VN496_in2 <= VN_sign_in(2978) & VN_data_in(2978);
  VN496_in3 <= VN_sign_in(2979) & VN_data_in(2979);
  VN496_in4 <= VN_sign_in(2980) & VN_data_in(2980);
  VN496_in5 <= VN_sign_in(2981) & VN_data_in(2981);
  VN497_in0 <= VN_sign_in(2982) & VN_data_in(2982);
  VN497_in1 <= VN_sign_in(2983) & VN_data_in(2983);
  VN497_in2 <= VN_sign_in(2984) & VN_data_in(2984);
  VN497_in3 <= VN_sign_in(2985) & VN_data_in(2985);
  VN497_in4 <= VN_sign_in(2986) & VN_data_in(2986);
  VN497_in5 <= VN_sign_in(2987) & VN_data_in(2987);
  VN498_in0 <= VN_sign_in(2988) & VN_data_in(2988);
  VN498_in1 <= VN_sign_in(2989) & VN_data_in(2989);
  VN498_in2 <= VN_sign_in(2990) & VN_data_in(2990);
  VN498_in3 <= VN_sign_in(2991) & VN_data_in(2991);
  VN498_in4 <= VN_sign_in(2992) & VN_data_in(2992);
  VN498_in5 <= VN_sign_in(2993) & VN_data_in(2993);
  VN499_in0 <= VN_sign_in(2994) & VN_data_in(2994);
  VN499_in1 <= VN_sign_in(2995) & VN_data_in(2995);
  VN499_in2 <= VN_sign_in(2996) & VN_data_in(2996);
  VN499_in3 <= VN_sign_in(2997) & VN_data_in(2997);
  VN499_in4 <= VN_sign_in(2998) & VN_data_in(2998);
  VN499_in5 <= VN_sign_in(2999) & VN_data_in(2999);
  VN500_in0 <= VN_sign_in(3000) & VN_data_in(3000);
  VN500_in1 <= VN_sign_in(3001) & VN_data_in(3001);
  VN500_in2 <= VN_sign_in(3002) & VN_data_in(3002);
  VN500_in3 <= VN_sign_in(3003) & VN_data_in(3003);
  VN500_in4 <= VN_sign_in(3004) & VN_data_in(3004);
  VN500_in5 <= VN_sign_in(3005) & VN_data_in(3005);
  VN501_in0 <= VN_sign_in(3006) & VN_data_in(3006);
  VN501_in1 <= VN_sign_in(3007) & VN_data_in(3007);
  VN501_in2 <= VN_sign_in(3008) & VN_data_in(3008);
  VN501_in3 <= VN_sign_in(3009) & VN_data_in(3009);
  VN501_in4 <= VN_sign_in(3010) & VN_data_in(3010);
  VN501_in5 <= VN_sign_in(3011) & VN_data_in(3011);
  VN502_in0 <= VN_sign_in(3012) & VN_data_in(3012);
  VN502_in1 <= VN_sign_in(3013) & VN_data_in(3013);
  VN502_in2 <= VN_sign_in(3014) & VN_data_in(3014);
  VN502_in3 <= VN_sign_in(3015) & VN_data_in(3015);
  VN502_in4 <= VN_sign_in(3016) & VN_data_in(3016);
  VN502_in5 <= VN_sign_in(3017) & VN_data_in(3017);
  VN503_in0 <= VN_sign_in(3018) & VN_data_in(3018);
  VN503_in1 <= VN_sign_in(3019) & VN_data_in(3019);
  VN503_in2 <= VN_sign_in(3020) & VN_data_in(3020);
  VN503_in3 <= VN_sign_in(3021) & VN_data_in(3021);
  VN503_in4 <= VN_sign_in(3022) & VN_data_in(3022);
  VN503_in5 <= VN_sign_in(3023) & VN_data_in(3023);
  VN504_in0 <= VN_sign_in(3024) & VN_data_in(3024);
  VN504_in1 <= VN_sign_in(3025) & VN_data_in(3025);
  VN504_in2 <= VN_sign_in(3026) & VN_data_in(3026);
  VN504_in3 <= VN_sign_in(3027) & VN_data_in(3027);
  VN504_in4 <= VN_sign_in(3028) & VN_data_in(3028);
  VN504_in5 <= VN_sign_in(3029) & VN_data_in(3029);
  VN505_in0 <= VN_sign_in(3030) & VN_data_in(3030);
  VN505_in1 <= VN_sign_in(3031) & VN_data_in(3031);
  VN505_in2 <= VN_sign_in(3032) & VN_data_in(3032);
  VN505_in3 <= VN_sign_in(3033) & VN_data_in(3033);
  VN505_in4 <= VN_sign_in(3034) & VN_data_in(3034);
  VN505_in5 <= VN_sign_in(3035) & VN_data_in(3035);
  VN506_in0 <= VN_sign_in(3036) & VN_data_in(3036);
  VN506_in1 <= VN_sign_in(3037) & VN_data_in(3037);
  VN506_in2 <= VN_sign_in(3038) & VN_data_in(3038);
  VN506_in3 <= VN_sign_in(3039) & VN_data_in(3039);
  VN506_in4 <= VN_sign_in(3040) & VN_data_in(3040);
  VN506_in5 <= VN_sign_in(3041) & VN_data_in(3041);
  VN507_in0 <= VN_sign_in(3042) & VN_data_in(3042);
  VN507_in1 <= VN_sign_in(3043) & VN_data_in(3043);
  VN507_in2 <= VN_sign_in(3044) & VN_data_in(3044);
  VN507_in3 <= VN_sign_in(3045) & VN_data_in(3045);
  VN507_in4 <= VN_sign_in(3046) & VN_data_in(3046);
  VN507_in5 <= VN_sign_in(3047) & VN_data_in(3047);
  VN508_in0 <= VN_sign_in(3048) & VN_data_in(3048);
  VN508_in1 <= VN_sign_in(3049) & VN_data_in(3049);
  VN508_in2 <= VN_sign_in(3050) & VN_data_in(3050);
  VN508_in3 <= VN_sign_in(3051) & VN_data_in(3051);
  VN508_in4 <= VN_sign_in(3052) & VN_data_in(3052);
  VN508_in5 <= VN_sign_in(3053) & VN_data_in(3053);
  VN509_in0 <= VN_sign_in(3054) & VN_data_in(3054);
  VN509_in1 <= VN_sign_in(3055) & VN_data_in(3055);
  VN509_in2 <= VN_sign_in(3056) & VN_data_in(3056);
  VN509_in3 <= VN_sign_in(3057) & VN_data_in(3057);
  VN509_in4 <= VN_sign_in(3058) & VN_data_in(3058);
  VN509_in5 <= VN_sign_in(3059) & VN_data_in(3059);
  VN510_in0 <= VN_sign_in(3060) & VN_data_in(3060);
  VN510_in1 <= VN_sign_in(3061) & VN_data_in(3061);
  VN510_in2 <= VN_sign_in(3062) & VN_data_in(3062);
  VN510_in3 <= VN_sign_in(3063) & VN_data_in(3063);
  VN510_in4 <= VN_sign_in(3064) & VN_data_in(3064);
  VN510_in5 <= VN_sign_in(3065) & VN_data_in(3065);
  VN511_in0 <= VN_sign_in(3066) & VN_data_in(3066);
  VN511_in1 <= VN_sign_in(3067) & VN_data_in(3067);
  VN511_in2 <= VN_sign_in(3068) & VN_data_in(3068);
  VN511_in3 <= VN_sign_in(3069) & VN_data_in(3069);
  VN511_in4 <= VN_sign_in(3070) & VN_data_in(3070);
  VN511_in5 <= VN_sign_in(3071) & VN_data_in(3071);
  VN512_in0 <= VN_sign_in(3072) & VN_data_in(3072);
  VN512_in1 <= VN_sign_in(3073) & VN_data_in(3073);
  VN512_in2 <= VN_sign_in(3074) & VN_data_in(3074);
  VN512_in3 <= VN_sign_in(3075) & VN_data_in(3075);
  VN512_in4 <= VN_sign_in(3076) & VN_data_in(3076);
  VN512_in5 <= VN_sign_in(3077) & VN_data_in(3077);
  VN513_in0 <= VN_sign_in(3078) & VN_data_in(3078);
  VN513_in1 <= VN_sign_in(3079) & VN_data_in(3079);
  VN513_in2 <= VN_sign_in(3080) & VN_data_in(3080);
  VN513_in3 <= VN_sign_in(3081) & VN_data_in(3081);
  VN513_in4 <= VN_sign_in(3082) & VN_data_in(3082);
  VN513_in5 <= VN_sign_in(3083) & VN_data_in(3083);
  VN514_in0 <= VN_sign_in(3084) & VN_data_in(3084);
  VN514_in1 <= VN_sign_in(3085) & VN_data_in(3085);
  VN514_in2 <= VN_sign_in(3086) & VN_data_in(3086);
  VN514_in3 <= VN_sign_in(3087) & VN_data_in(3087);
  VN514_in4 <= VN_sign_in(3088) & VN_data_in(3088);
  VN514_in5 <= VN_sign_in(3089) & VN_data_in(3089);
  VN515_in0 <= VN_sign_in(3090) & VN_data_in(3090);
  VN515_in1 <= VN_sign_in(3091) & VN_data_in(3091);
  VN515_in2 <= VN_sign_in(3092) & VN_data_in(3092);
  VN515_in3 <= VN_sign_in(3093) & VN_data_in(3093);
  VN515_in4 <= VN_sign_in(3094) & VN_data_in(3094);
  VN515_in5 <= VN_sign_in(3095) & VN_data_in(3095);
  VN516_in0 <= VN_sign_in(3096) & VN_data_in(3096);
  VN516_in1 <= VN_sign_in(3097) & VN_data_in(3097);
  VN516_in2 <= VN_sign_in(3098) & VN_data_in(3098);
  VN516_in3 <= VN_sign_in(3099) & VN_data_in(3099);
  VN516_in4 <= VN_sign_in(3100) & VN_data_in(3100);
  VN516_in5 <= VN_sign_in(3101) & VN_data_in(3101);
  VN517_in0 <= VN_sign_in(3102) & VN_data_in(3102);
  VN517_in1 <= VN_sign_in(3103) & VN_data_in(3103);
  VN517_in2 <= VN_sign_in(3104) & VN_data_in(3104);
  VN517_in3 <= VN_sign_in(3105) & VN_data_in(3105);
  VN517_in4 <= VN_sign_in(3106) & VN_data_in(3106);
  VN517_in5 <= VN_sign_in(3107) & VN_data_in(3107);
  VN518_in0 <= VN_sign_in(3108) & VN_data_in(3108);
  VN518_in1 <= VN_sign_in(3109) & VN_data_in(3109);
  VN518_in2 <= VN_sign_in(3110) & VN_data_in(3110);
  VN518_in3 <= VN_sign_in(3111) & VN_data_in(3111);
  VN518_in4 <= VN_sign_in(3112) & VN_data_in(3112);
  VN518_in5 <= VN_sign_in(3113) & VN_data_in(3113);
  VN519_in0 <= VN_sign_in(3114) & VN_data_in(3114);
  VN519_in1 <= VN_sign_in(3115) & VN_data_in(3115);
  VN519_in2 <= VN_sign_in(3116) & VN_data_in(3116);
  VN519_in3 <= VN_sign_in(3117) & VN_data_in(3117);
  VN519_in4 <= VN_sign_in(3118) & VN_data_in(3118);
  VN519_in5 <= VN_sign_in(3119) & VN_data_in(3119);
  VN520_in0 <= VN_sign_in(3120) & VN_data_in(3120);
  VN520_in1 <= VN_sign_in(3121) & VN_data_in(3121);
  VN520_in2 <= VN_sign_in(3122) & VN_data_in(3122);
  VN520_in3 <= VN_sign_in(3123) & VN_data_in(3123);
  VN520_in4 <= VN_sign_in(3124) & VN_data_in(3124);
  VN520_in5 <= VN_sign_in(3125) & VN_data_in(3125);
  VN521_in0 <= VN_sign_in(3126) & VN_data_in(3126);
  VN521_in1 <= VN_sign_in(3127) & VN_data_in(3127);
  VN521_in2 <= VN_sign_in(3128) & VN_data_in(3128);
  VN521_in3 <= VN_sign_in(3129) & VN_data_in(3129);
  VN521_in4 <= VN_sign_in(3130) & VN_data_in(3130);
  VN521_in5 <= VN_sign_in(3131) & VN_data_in(3131);
  VN522_in0 <= VN_sign_in(3132) & VN_data_in(3132);
  VN522_in1 <= VN_sign_in(3133) & VN_data_in(3133);
  VN522_in2 <= VN_sign_in(3134) & VN_data_in(3134);
  VN522_in3 <= VN_sign_in(3135) & VN_data_in(3135);
  VN522_in4 <= VN_sign_in(3136) & VN_data_in(3136);
  VN522_in5 <= VN_sign_in(3137) & VN_data_in(3137);
  VN523_in0 <= VN_sign_in(3138) & VN_data_in(3138);
  VN523_in1 <= VN_sign_in(3139) & VN_data_in(3139);
  VN523_in2 <= VN_sign_in(3140) & VN_data_in(3140);
  VN523_in3 <= VN_sign_in(3141) & VN_data_in(3141);
  VN523_in4 <= VN_sign_in(3142) & VN_data_in(3142);
  VN523_in5 <= VN_sign_in(3143) & VN_data_in(3143);
  VN524_in0 <= VN_sign_in(3144) & VN_data_in(3144);
  VN524_in1 <= VN_sign_in(3145) & VN_data_in(3145);
  VN524_in2 <= VN_sign_in(3146) & VN_data_in(3146);
  VN524_in3 <= VN_sign_in(3147) & VN_data_in(3147);
  VN524_in4 <= VN_sign_in(3148) & VN_data_in(3148);
  VN524_in5 <= VN_sign_in(3149) & VN_data_in(3149);
  VN525_in0 <= VN_sign_in(3150) & VN_data_in(3150);
  VN525_in1 <= VN_sign_in(3151) & VN_data_in(3151);
  VN525_in2 <= VN_sign_in(3152) & VN_data_in(3152);
  VN525_in3 <= VN_sign_in(3153) & VN_data_in(3153);
  VN525_in4 <= VN_sign_in(3154) & VN_data_in(3154);
  VN525_in5 <= VN_sign_in(3155) & VN_data_in(3155);
  VN526_in0 <= VN_sign_in(3156) & VN_data_in(3156);
  VN526_in1 <= VN_sign_in(3157) & VN_data_in(3157);
  VN526_in2 <= VN_sign_in(3158) & VN_data_in(3158);
  VN526_in3 <= VN_sign_in(3159) & VN_data_in(3159);
  VN526_in4 <= VN_sign_in(3160) & VN_data_in(3160);
  VN526_in5 <= VN_sign_in(3161) & VN_data_in(3161);
  VN527_in0 <= VN_sign_in(3162) & VN_data_in(3162);
  VN527_in1 <= VN_sign_in(3163) & VN_data_in(3163);
  VN527_in2 <= VN_sign_in(3164) & VN_data_in(3164);
  VN527_in3 <= VN_sign_in(3165) & VN_data_in(3165);
  VN527_in4 <= VN_sign_in(3166) & VN_data_in(3166);
  VN527_in5 <= VN_sign_in(3167) & VN_data_in(3167);
  VN528_in0 <= VN_sign_in(3168) & VN_data_in(3168);
  VN528_in1 <= VN_sign_in(3169) & VN_data_in(3169);
  VN528_in2 <= VN_sign_in(3170) & VN_data_in(3170);
  VN528_in3 <= VN_sign_in(3171) & VN_data_in(3171);
  VN528_in4 <= VN_sign_in(3172) & VN_data_in(3172);
  VN528_in5 <= VN_sign_in(3173) & VN_data_in(3173);
  VN529_in0 <= VN_sign_in(3174) & VN_data_in(3174);
  VN529_in1 <= VN_sign_in(3175) & VN_data_in(3175);
  VN529_in2 <= VN_sign_in(3176) & VN_data_in(3176);
  VN529_in3 <= VN_sign_in(3177) & VN_data_in(3177);
  VN529_in4 <= VN_sign_in(3178) & VN_data_in(3178);
  VN529_in5 <= VN_sign_in(3179) & VN_data_in(3179);
  VN530_in0 <= VN_sign_in(3180) & VN_data_in(3180);
  VN530_in1 <= VN_sign_in(3181) & VN_data_in(3181);
  VN530_in2 <= VN_sign_in(3182) & VN_data_in(3182);
  VN530_in3 <= VN_sign_in(3183) & VN_data_in(3183);
  VN530_in4 <= VN_sign_in(3184) & VN_data_in(3184);
  VN530_in5 <= VN_sign_in(3185) & VN_data_in(3185);
  VN531_in0 <= VN_sign_in(3186) & VN_data_in(3186);
  VN531_in1 <= VN_sign_in(3187) & VN_data_in(3187);
  VN531_in2 <= VN_sign_in(3188) & VN_data_in(3188);
  VN531_in3 <= VN_sign_in(3189) & VN_data_in(3189);
  VN531_in4 <= VN_sign_in(3190) & VN_data_in(3190);
  VN531_in5 <= VN_sign_in(3191) & VN_data_in(3191);
  VN532_in0 <= VN_sign_in(3192) & VN_data_in(3192);
  VN532_in1 <= VN_sign_in(3193) & VN_data_in(3193);
  VN532_in2 <= VN_sign_in(3194) & VN_data_in(3194);
  VN532_in3 <= VN_sign_in(3195) & VN_data_in(3195);
  VN532_in4 <= VN_sign_in(3196) & VN_data_in(3196);
  VN532_in5 <= VN_sign_in(3197) & VN_data_in(3197);
  VN533_in0 <= VN_sign_in(3198) & VN_data_in(3198);
  VN533_in1 <= VN_sign_in(3199) & VN_data_in(3199);
  VN533_in2 <= VN_sign_in(3200) & VN_data_in(3200);
  VN533_in3 <= VN_sign_in(3201) & VN_data_in(3201);
  VN533_in4 <= VN_sign_in(3202) & VN_data_in(3202);
  VN533_in5 <= VN_sign_in(3203) & VN_data_in(3203);
  VN534_in0 <= VN_sign_in(3204) & VN_data_in(3204);
  VN534_in1 <= VN_sign_in(3205) & VN_data_in(3205);
  VN534_in2 <= VN_sign_in(3206) & VN_data_in(3206);
  VN534_in3 <= VN_sign_in(3207) & VN_data_in(3207);
  VN534_in4 <= VN_sign_in(3208) & VN_data_in(3208);
  VN534_in5 <= VN_sign_in(3209) & VN_data_in(3209);
  VN535_in0 <= VN_sign_in(3210) & VN_data_in(3210);
  VN535_in1 <= VN_sign_in(3211) & VN_data_in(3211);
  VN535_in2 <= VN_sign_in(3212) & VN_data_in(3212);
  VN535_in3 <= VN_sign_in(3213) & VN_data_in(3213);
  VN535_in4 <= VN_sign_in(3214) & VN_data_in(3214);
  VN535_in5 <= VN_sign_in(3215) & VN_data_in(3215);
  VN536_in0 <= VN_sign_in(3216) & VN_data_in(3216);
  VN536_in1 <= VN_sign_in(3217) & VN_data_in(3217);
  VN536_in2 <= VN_sign_in(3218) & VN_data_in(3218);
  VN536_in3 <= VN_sign_in(3219) & VN_data_in(3219);
  VN536_in4 <= VN_sign_in(3220) & VN_data_in(3220);
  VN536_in5 <= VN_sign_in(3221) & VN_data_in(3221);
  VN537_in0 <= VN_sign_in(3222) & VN_data_in(3222);
  VN537_in1 <= VN_sign_in(3223) & VN_data_in(3223);
  VN537_in2 <= VN_sign_in(3224) & VN_data_in(3224);
  VN537_in3 <= VN_sign_in(3225) & VN_data_in(3225);
  VN537_in4 <= VN_sign_in(3226) & VN_data_in(3226);
  VN537_in5 <= VN_sign_in(3227) & VN_data_in(3227);
  VN538_in0 <= VN_sign_in(3228) & VN_data_in(3228);
  VN538_in1 <= VN_sign_in(3229) & VN_data_in(3229);
  VN538_in2 <= VN_sign_in(3230) & VN_data_in(3230);
  VN538_in3 <= VN_sign_in(3231) & VN_data_in(3231);
  VN538_in4 <= VN_sign_in(3232) & VN_data_in(3232);
  VN538_in5 <= VN_sign_in(3233) & VN_data_in(3233);
  VN539_in0 <= VN_sign_in(3234) & VN_data_in(3234);
  VN539_in1 <= VN_sign_in(3235) & VN_data_in(3235);
  VN539_in2 <= VN_sign_in(3236) & VN_data_in(3236);
  VN539_in3 <= VN_sign_in(3237) & VN_data_in(3237);
  VN539_in4 <= VN_sign_in(3238) & VN_data_in(3238);
  VN539_in5 <= VN_sign_in(3239) & VN_data_in(3239);
  VN540_in0 <= VN_sign_in(3240) & VN_data_in(3240);
  VN540_in1 <= VN_sign_in(3241) & VN_data_in(3241);
  VN540_in2 <= VN_sign_in(3242) & VN_data_in(3242);
  VN540_in3 <= VN_sign_in(3243) & VN_data_in(3243);
  VN540_in4 <= VN_sign_in(3244) & VN_data_in(3244);
  VN540_in5 <= VN_sign_in(3245) & VN_data_in(3245);
  VN541_in0 <= VN_sign_in(3246) & VN_data_in(3246);
  VN541_in1 <= VN_sign_in(3247) & VN_data_in(3247);
  VN541_in2 <= VN_sign_in(3248) & VN_data_in(3248);
  VN541_in3 <= VN_sign_in(3249) & VN_data_in(3249);
  VN541_in4 <= VN_sign_in(3250) & VN_data_in(3250);
  VN541_in5 <= VN_sign_in(3251) & VN_data_in(3251);
  VN542_in0 <= VN_sign_in(3252) & VN_data_in(3252);
  VN542_in1 <= VN_sign_in(3253) & VN_data_in(3253);
  VN542_in2 <= VN_sign_in(3254) & VN_data_in(3254);
  VN542_in3 <= VN_sign_in(3255) & VN_data_in(3255);
  VN542_in4 <= VN_sign_in(3256) & VN_data_in(3256);
  VN542_in5 <= VN_sign_in(3257) & VN_data_in(3257);
  VN543_in0 <= VN_sign_in(3258) & VN_data_in(3258);
  VN543_in1 <= VN_sign_in(3259) & VN_data_in(3259);
  VN543_in2 <= VN_sign_in(3260) & VN_data_in(3260);
  VN543_in3 <= VN_sign_in(3261) & VN_data_in(3261);
  VN543_in4 <= VN_sign_in(3262) & VN_data_in(3262);
  VN543_in5 <= VN_sign_in(3263) & VN_data_in(3263);
  VN544_in0 <= VN_sign_in(3264) & VN_data_in(3264);
  VN544_in1 <= VN_sign_in(3265) & VN_data_in(3265);
  VN544_in2 <= VN_sign_in(3266) & VN_data_in(3266);
  VN544_in3 <= VN_sign_in(3267) & VN_data_in(3267);
  VN544_in4 <= VN_sign_in(3268) & VN_data_in(3268);
  VN544_in5 <= VN_sign_in(3269) & VN_data_in(3269);
  VN545_in0 <= VN_sign_in(3270) & VN_data_in(3270);
  VN545_in1 <= VN_sign_in(3271) & VN_data_in(3271);
  VN545_in2 <= VN_sign_in(3272) & VN_data_in(3272);
  VN545_in3 <= VN_sign_in(3273) & VN_data_in(3273);
  VN545_in4 <= VN_sign_in(3274) & VN_data_in(3274);
  VN545_in5 <= VN_sign_in(3275) & VN_data_in(3275);
  VN546_in0 <= VN_sign_in(3276) & VN_data_in(3276);
  VN546_in1 <= VN_sign_in(3277) & VN_data_in(3277);
  VN546_in2 <= VN_sign_in(3278) & VN_data_in(3278);
  VN546_in3 <= VN_sign_in(3279) & VN_data_in(3279);
  VN546_in4 <= VN_sign_in(3280) & VN_data_in(3280);
  VN546_in5 <= VN_sign_in(3281) & VN_data_in(3281);
  VN547_in0 <= VN_sign_in(3282) & VN_data_in(3282);
  VN547_in1 <= VN_sign_in(3283) & VN_data_in(3283);
  VN547_in2 <= VN_sign_in(3284) & VN_data_in(3284);
  VN547_in3 <= VN_sign_in(3285) & VN_data_in(3285);
  VN547_in4 <= VN_sign_in(3286) & VN_data_in(3286);
  VN547_in5 <= VN_sign_in(3287) & VN_data_in(3287);
  VN548_in0 <= VN_sign_in(3288) & VN_data_in(3288);
  VN548_in1 <= VN_sign_in(3289) & VN_data_in(3289);
  VN548_in2 <= VN_sign_in(3290) & VN_data_in(3290);
  VN548_in3 <= VN_sign_in(3291) & VN_data_in(3291);
  VN548_in4 <= VN_sign_in(3292) & VN_data_in(3292);
  VN548_in5 <= VN_sign_in(3293) & VN_data_in(3293);
  VN549_in0 <= VN_sign_in(3294) & VN_data_in(3294);
  VN549_in1 <= VN_sign_in(3295) & VN_data_in(3295);
  VN549_in2 <= VN_sign_in(3296) & VN_data_in(3296);
  VN549_in3 <= VN_sign_in(3297) & VN_data_in(3297);
  VN549_in4 <= VN_sign_in(3298) & VN_data_in(3298);
  VN549_in5 <= VN_sign_in(3299) & VN_data_in(3299);
  VN550_in0 <= VN_sign_in(3300) & VN_data_in(3300);
  VN550_in1 <= VN_sign_in(3301) & VN_data_in(3301);
  VN550_in2 <= VN_sign_in(3302) & VN_data_in(3302);
  VN550_in3 <= VN_sign_in(3303) & VN_data_in(3303);
  VN550_in4 <= VN_sign_in(3304) & VN_data_in(3304);
  VN550_in5 <= VN_sign_in(3305) & VN_data_in(3305);
  VN551_in0 <= VN_sign_in(3306) & VN_data_in(3306);
  VN551_in1 <= VN_sign_in(3307) & VN_data_in(3307);
  VN551_in2 <= VN_sign_in(3308) & VN_data_in(3308);
  VN551_in3 <= VN_sign_in(3309) & VN_data_in(3309);
  VN551_in4 <= VN_sign_in(3310) & VN_data_in(3310);
  VN551_in5 <= VN_sign_in(3311) & VN_data_in(3311);
  VN552_in0 <= VN_sign_in(3312) & VN_data_in(3312);
  VN552_in1 <= VN_sign_in(3313) & VN_data_in(3313);
  VN552_in2 <= VN_sign_in(3314) & VN_data_in(3314);
  VN552_in3 <= VN_sign_in(3315) & VN_data_in(3315);
  VN552_in4 <= VN_sign_in(3316) & VN_data_in(3316);
  VN552_in5 <= VN_sign_in(3317) & VN_data_in(3317);
  VN553_in0 <= VN_sign_in(3318) & VN_data_in(3318);
  VN553_in1 <= VN_sign_in(3319) & VN_data_in(3319);
  VN553_in2 <= VN_sign_in(3320) & VN_data_in(3320);
  VN553_in3 <= VN_sign_in(3321) & VN_data_in(3321);
  VN553_in4 <= VN_sign_in(3322) & VN_data_in(3322);
  VN553_in5 <= VN_sign_in(3323) & VN_data_in(3323);
  VN554_in0 <= VN_sign_in(3324) & VN_data_in(3324);
  VN554_in1 <= VN_sign_in(3325) & VN_data_in(3325);
  VN554_in2 <= VN_sign_in(3326) & VN_data_in(3326);
  VN554_in3 <= VN_sign_in(3327) & VN_data_in(3327);
  VN554_in4 <= VN_sign_in(3328) & VN_data_in(3328);
  VN554_in5 <= VN_sign_in(3329) & VN_data_in(3329);
  VN555_in0 <= VN_sign_in(3330) & VN_data_in(3330);
  VN555_in1 <= VN_sign_in(3331) & VN_data_in(3331);
  VN555_in2 <= VN_sign_in(3332) & VN_data_in(3332);
  VN555_in3 <= VN_sign_in(3333) & VN_data_in(3333);
  VN555_in4 <= VN_sign_in(3334) & VN_data_in(3334);
  VN555_in5 <= VN_sign_in(3335) & VN_data_in(3335);
  VN556_in0 <= VN_sign_in(3336) & VN_data_in(3336);
  VN556_in1 <= VN_sign_in(3337) & VN_data_in(3337);
  VN556_in2 <= VN_sign_in(3338) & VN_data_in(3338);
  VN556_in3 <= VN_sign_in(3339) & VN_data_in(3339);
  VN556_in4 <= VN_sign_in(3340) & VN_data_in(3340);
  VN556_in5 <= VN_sign_in(3341) & VN_data_in(3341);
  VN557_in0 <= VN_sign_in(3342) & VN_data_in(3342);
  VN557_in1 <= VN_sign_in(3343) & VN_data_in(3343);
  VN557_in2 <= VN_sign_in(3344) & VN_data_in(3344);
  VN557_in3 <= VN_sign_in(3345) & VN_data_in(3345);
  VN557_in4 <= VN_sign_in(3346) & VN_data_in(3346);
  VN557_in5 <= VN_sign_in(3347) & VN_data_in(3347);
  VN558_in0 <= VN_sign_in(3348) & VN_data_in(3348);
  VN558_in1 <= VN_sign_in(3349) & VN_data_in(3349);
  VN558_in2 <= VN_sign_in(3350) & VN_data_in(3350);
  VN558_in3 <= VN_sign_in(3351) & VN_data_in(3351);
  VN558_in4 <= VN_sign_in(3352) & VN_data_in(3352);
  VN558_in5 <= VN_sign_in(3353) & VN_data_in(3353);
  VN559_in0 <= VN_sign_in(3354) & VN_data_in(3354);
  VN559_in1 <= VN_sign_in(3355) & VN_data_in(3355);
  VN559_in2 <= VN_sign_in(3356) & VN_data_in(3356);
  VN559_in3 <= VN_sign_in(3357) & VN_data_in(3357);
  VN559_in4 <= VN_sign_in(3358) & VN_data_in(3358);
  VN559_in5 <= VN_sign_in(3359) & VN_data_in(3359);
  VN560_in0 <= VN_sign_in(3360) & VN_data_in(3360);
  VN560_in1 <= VN_sign_in(3361) & VN_data_in(3361);
  VN560_in2 <= VN_sign_in(3362) & VN_data_in(3362);
  VN560_in3 <= VN_sign_in(3363) & VN_data_in(3363);
  VN560_in4 <= VN_sign_in(3364) & VN_data_in(3364);
  VN560_in5 <= VN_sign_in(3365) & VN_data_in(3365);
  VN561_in0 <= VN_sign_in(3366) & VN_data_in(3366);
  VN561_in1 <= VN_sign_in(3367) & VN_data_in(3367);
  VN561_in2 <= VN_sign_in(3368) & VN_data_in(3368);
  VN561_in3 <= VN_sign_in(3369) & VN_data_in(3369);
  VN561_in4 <= VN_sign_in(3370) & VN_data_in(3370);
  VN561_in5 <= VN_sign_in(3371) & VN_data_in(3371);
  VN562_in0 <= VN_sign_in(3372) & VN_data_in(3372);
  VN562_in1 <= VN_sign_in(3373) & VN_data_in(3373);
  VN562_in2 <= VN_sign_in(3374) & VN_data_in(3374);
  VN562_in3 <= VN_sign_in(3375) & VN_data_in(3375);
  VN562_in4 <= VN_sign_in(3376) & VN_data_in(3376);
  VN562_in5 <= VN_sign_in(3377) & VN_data_in(3377);
  VN563_in0 <= VN_sign_in(3378) & VN_data_in(3378);
  VN563_in1 <= VN_sign_in(3379) & VN_data_in(3379);
  VN563_in2 <= VN_sign_in(3380) & VN_data_in(3380);
  VN563_in3 <= VN_sign_in(3381) & VN_data_in(3381);
  VN563_in4 <= VN_sign_in(3382) & VN_data_in(3382);
  VN563_in5 <= VN_sign_in(3383) & VN_data_in(3383);
  VN564_in0 <= VN_sign_in(3384) & VN_data_in(3384);
  VN564_in1 <= VN_sign_in(3385) & VN_data_in(3385);
  VN564_in2 <= VN_sign_in(3386) & VN_data_in(3386);
  VN564_in3 <= VN_sign_in(3387) & VN_data_in(3387);
  VN564_in4 <= VN_sign_in(3388) & VN_data_in(3388);
  VN564_in5 <= VN_sign_in(3389) & VN_data_in(3389);
  VN565_in0 <= VN_sign_in(3390) & VN_data_in(3390);
  VN565_in1 <= VN_sign_in(3391) & VN_data_in(3391);
  VN565_in2 <= VN_sign_in(3392) & VN_data_in(3392);
  VN565_in3 <= VN_sign_in(3393) & VN_data_in(3393);
  VN565_in4 <= VN_sign_in(3394) & VN_data_in(3394);
  VN565_in5 <= VN_sign_in(3395) & VN_data_in(3395);
  VN566_in0 <= VN_sign_in(3396) & VN_data_in(3396);
  VN566_in1 <= VN_sign_in(3397) & VN_data_in(3397);
  VN566_in2 <= VN_sign_in(3398) & VN_data_in(3398);
  VN566_in3 <= VN_sign_in(3399) & VN_data_in(3399);
  VN566_in4 <= VN_sign_in(3400) & VN_data_in(3400);
  VN566_in5 <= VN_sign_in(3401) & VN_data_in(3401);
  VN567_in0 <= VN_sign_in(3402) & VN_data_in(3402);
  VN567_in1 <= VN_sign_in(3403) & VN_data_in(3403);
  VN567_in2 <= VN_sign_in(3404) & VN_data_in(3404);
  VN567_in3 <= VN_sign_in(3405) & VN_data_in(3405);
  VN567_in4 <= VN_sign_in(3406) & VN_data_in(3406);
  VN567_in5 <= VN_sign_in(3407) & VN_data_in(3407);
  VN568_in0 <= VN_sign_in(3408) & VN_data_in(3408);
  VN568_in1 <= VN_sign_in(3409) & VN_data_in(3409);
  VN568_in2 <= VN_sign_in(3410) & VN_data_in(3410);
  VN568_in3 <= VN_sign_in(3411) & VN_data_in(3411);
  VN568_in4 <= VN_sign_in(3412) & VN_data_in(3412);
  VN568_in5 <= VN_sign_in(3413) & VN_data_in(3413);
  VN569_in0 <= VN_sign_in(3414) & VN_data_in(3414);
  VN569_in1 <= VN_sign_in(3415) & VN_data_in(3415);
  VN569_in2 <= VN_sign_in(3416) & VN_data_in(3416);
  VN569_in3 <= VN_sign_in(3417) & VN_data_in(3417);
  VN569_in4 <= VN_sign_in(3418) & VN_data_in(3418);
  VN569_in5 <= VN_sign_in(3419) & VN_data_in(3419);
  VN570_in0 <= VN_sign_in(3420) & VN_data_in(3420);
  VN570_in1 <= VN_sign_in(3421) & VN_data_in(3421);
  VN570_in2 <= VN_sign_in(3422) & VN_data_in(3422);
  VN570_in3 <= VN_sign_in(3423) & VN_data_in(3423);
  VN570_in4 <= VN_sign_in(3424) & VN_data_in(3424);
  VN570_in5 <= VN_sign_in(3425) & VN_data_in(3425);
  VN571_in0 <= VN_sign_in(3426) & VN_data_in(3426);
  VN571_in1 <= VN_sign_in(3427) & VN_data_in(3427);
  VN571_in2 <= VN_sign_in(3428) & VN_data_in(3428);
  VN571_in3 <= VN_sign_in(3429) & VN_data_in(3429);
  VN571_in4 <= VN_sign_in(3430) & VN_data_in(3430);
  VN571_in5 <= VN_sign_in(3431) & VN_data_in(3431);
  VN572_in0 <= VN_sign_in(3432) & VN_data_in(3432);
  VN572_in1 <= VN_sign_in(3433) & VN_data_in(3433);
  VN572_in2 <= VN_sign_in(3434) & VN_data_in(3434);
  VN572_in3 <= VN_sign_in(3435) & VN_data_in(3435);
  VN572_in4 <= VN_sign_in(3436) & VN_data_in(3436);
  VN572_in5 <= VN_sign_in(3437) & VN_data_in(3437);
  VN573_in0 <= VN_sign_in(3438) & VN_data_in(3438);
  VN573_in1 <= VN_sign_in(3439) & VN_data_in(3439);
  VN573_in2 <= VN_sign_in(3440) & VN_data_in(3440);
  VN573_in3 <= VN_sign_in(3441) & VN_data_in(3441);
  VN573_in4 <= VN_sign_in(3442) & VN_data_in(3442);
  VN573_in5 <= VN_sign_in(3443) & VN_data_in(3443);
  VN574_in0 <= VN_sign_in(3444) & VN_data_in(3444);
  VN574_in1 <= VN_sign_in(3445) & VN_data_in(3445);
  VN574_in2 <= VN_sign_in(3446) & VN_data_in(3446);
  VN574_in3 <= VN_sign_in(3447) & VN_data_in(3447);
  VN574_in4 <= VN_sign_in(3448) & VN_data_in(3448);
  VN574_in5 <= VN_sign_in(3449) & VN_data_in(3449);
  VN575_in0 <= VN_sign_in(3450) & VN_data_in(3450);
  VN575_in1 <= VN_sign_in(3451) & VN_data_in(3451);
  VN575_in2 <= VN_sign_in(3452) & VN_data_in(3452);
  VN575_in3 <= VN_sign_in(3453) & VN_data_in(3453);
  VN575_in4 <= VN_sign_in(3454) & VN_data_in(3454);
  VN575_in5 <= VN_sign_in(3455) & VN_data_in(3455);
  VN576_in0 <= VN_sign_in(3456) & VN_data_in(3456);
  VN576_in1 <= VN_sign_in(3457) & VN_data_in(3457);
  VN576_in2 <= VN_sign_in(3458) & VN_data_in(3458);
  VN576_in3 <= VN_sign_in(3459) & VN_data_in(3459);
  VN576_in4 <= VN_sign_in(3460) & VN_data_in(3460);
  VN576_in5 <= VN_sign_in(3461) & VN_data_in(3461);
  VN577_in0 <= VN_sign_in(3462) & VN_data_in(3462);
  VN577_in1 <= VN_sign_in(3463) & VN_data_in(3463);
  VN577_in2 <= VN_sign_in(3464) & VN_data_in(3464);
  VN577_in3 <= VN_sign_in(3465) & VN_data_in(3465);
  VN577_in4 <= VN_sign_in(3466) & VN_data_in(3466);
  VN577_in5 <= VN_sign_in(3467) & VN_data_in(3467);
  VN578_in0 <= VN_sign_in(3468) & VN_data_in(3468);
  VN578_in1 <= VN_sign_in(3469) & VN_data_in(3469);
  VN578_in2 <= VN_sign_in(3470) & VN_data_in(3470);
  VN578_in3 <= VN_sign_in(3471) & VN_data_in(3471);
  VN578_in4 <= VN_sign_in(3472) & VN_data_in(3472);
  VN578_in5 <= VN_sign_in(3473) & VN_data_in(3473);
  VN579_in0 <= VN_sign_in(3474) & VN_data_in(3474);
  VN579_in1 <= VN_sign_in(3475) & VN_data_in(3475);
  VN579_in2 <= VN_sign_in(3476) & VN_data_in(3476);
  VN579_in3 <= VN_sign_in(3477) & VN_data_in(3477);
  VN579_in4 <= VN_sign_in(3478) & VN_data_in(3478);
  VN579_in5 <= VN_sign_in(3479) & VN_data_in(3479);
  VN580_in0 <= VN_sign_in(3480) & VN_data_in(3480);
  VN580_in1 <= VN_sign_in(3481) & VN_data_in(3481);
  VN580_in2 <= VN_sign_in(3482) & VN_data_in(3482);
  VN580_in3 <= VN_sign_in(3483) & VN_data_in(3483);
  VN580_in4 <= VN_sign_in(3484) & VN_data_in(3484);
  VN580_in5 <= VN_sign_in(3485) & VN_data_in(3485);
  VN581_in0 <= VN_sign_in(3486) & VN_data_in(3486);
  VN581_in1 <= VN_sign_in(3487) & VN_data_in(3487);
  VN581_in2 <= VN_sign_in(3488) & VN_data_in(3488);
  VN581_in3 <= VN_sign_in(3489) & VN_data_in(3489);
  VN581_in4 <= VN_sign_in(3490) & VN_data_in(3490);
  VN581_in5 <= VN_sign_in(3491) & VN_data_in(3491);
  VN582_in0 <= VN_sign_in(3492) & VN_data_in(3492);
  VN582_in1 <= VN_sign_in(3493) & VN_data_in(3493);
  VN582_in2 <= VN_sign_in(3494) & VN_data_in(3494);
  VN582_in3 <= VN_sign_in(3495) & VN_data_in(3495);
  VN582_in4 <= VN_sign_in(3496) & VN_data_in(3496);
  VN582_in5 <= VN_sign_in(3497) & VN_data_in(3497);
  VN583_in0 <= VN_sign_in(3498) & VN_data_in(3498);
  VN583_in1 <= VN_sign_in(3499) & VN_data_in(3499);
  VN583_in2 <= VN_sign_in(3500) & VN_data_in(3500);
  VN583_in3 <= VN_sign_in(3501) & VN_data_in(3501);
  VN583_in4 <= VN_sign_in(3502) & VN_data_in(3502);
  VN583_in5 <= VN_sign_in(3503) & VN_data_in(3503);
  VN584_in0 <= VN_sign_in(3504) & VN_data_in(3504);
  VN584_in1 <= VN_sign_in(3505) & VN_data_in(3505);
  VN584_in2 <= VN_sign_in(3506) & VN_data_in(3506);
  VN584_in3 <= VN_sign_in(3507) & VN_data_in(3507);
  VN584_in4 <= VN_sign_in(3508) & VN_data_in(3508);
  VN584_in5 <= VN_sign_in(3509) & VN_data_in(3509);
  VN585_in0 <= VN_sign_in(3510) & VN_data_in(3510);
  VN585_in1 <= VN_sign_in(3511) & VN_data_in(3511);
  VN585_in2 <= VN_sign_in(3512) & VN_data_in(3512);
  VN585_in3 <= VN_sign_in(3513) & VN_data_in(3513);
  VN585_in4 <= VN_sign_in(3514) & VN_data_in(3514);
  VN585_in5 <= VN_sign_in(3515) & VN_data_in(3515);
  VN586_in0 <= VN_sign_in(3516) & VN_data_in(3516);
  VN586_in1 <= VN_sign_in(3517) & VN_data_in(3517);
  VN586_in2 <= VN_sign_in(3518) & VN_data_in(3518);
  VN586_in3 <= VN_sign_in(3519) & VN_data_in(3519);
  VN586_in4 <= VN_sign_in(3520) & VN_data_in(3520);
  VN586_in5 <= VN_sign_in(3521) & VN_data_in(3521);
  VN587_in0 <= VN_sign_in(3522) & VN_data_in(3522);
  VN587_in1 <= VN_sign_in(3523) & VN_data_in(3523);
  VN587_in2 <= VN_sign_in(3524) & VN_data_in(3524);
  VN587_in3 <= VN_sign_in(3525) & VN_data_in(3525);
  VN587_in4 <= VN_sign_in(3526) & VN_data_in(3526);
  VN587_in5 <= VN_sign_in(3527) & VN_data_in(3527);
  VN588_in0 <= VN_sign_in(3528) & VN_data_in(3528);
  VN588_in1 <= VN_sign_in(3529) & VN_data_in(3529);
  VN588_in2 <= VN_sign_in(3530) & VN_data_in(3530);
  VN588_in3 <= VN_sign_in(3531) & VN_data_in(3531);
  VN588_in4 <= VN_sign_in(3532) & VN_data_in(3532);
  VN588_in5 <= VN_sign_in(3533) & VN_data_in(3533);
  VN589_in0 <= VN_sign_in(3534) & VN_data_in(3534);
  VN589_in1 <= VN_sign_in(3535) & VN_data_in(3535);
  VN589_in2 <= VN_sign_in(3536) & VN_data_in(3536);
  VN589_in3 <= VN_sign_in(3537) & VN_data_in(3537);
  VN589_in4 <= VN_sign_in(3538) & VN_data_in(3538);
  VN589_in5 <= VN_sign_in(3539) & VN_data_in(3539);
  VN590_in0 <= VN_sign_in(3540) & VN_data_in(3540);
  VN590_in1 <= VN_sign_in(3541) & VN_data_in(3541);
  VN590_in2 <= VN_sign_in(3542) & VN_data_in(3542);
  VN590_in3 <= VN_sign_in(3543) & VN_data_in(3543);
  VN590_in4 <= VN_sign_in(3544) & VN_data_in(3544);
  VN590_in5 <= VN_sign_in(3545) & VN_data_in(3545);
  VN591_in0 <= VN_sign_in(3546) & VN_data_in(3546);
  VN591_in1 <= VN_sign_in(3547) & VN_data_in(3547);
  VN591_in2 <= VN_sign_in(3548) & VN_data_in(3548);
  VN591_in3 <= VN_sign_in(3549) & VN_data_in(3549);
  VN591_in4 <= VN_sign_in(3550) & VN_data_in(3550);
  VN591_in5 <= VN_sign_in(3551) & VN_data_in(3551);
  VN592_in0 <= VN_sign_in(3552) & VN_data_in(3552);
  VN592_in1 <= VN_sign_in(3553) & VN_data_in(3553);
  VN592_in2 <= VN_sign_in(3554) & VN_data_in(3554);
  VN592_in3 <= VN_sign_in(3555) & VN_data_in(3555);
  VN592_in4 <= VN_sign_in(3556) & VN_data_in(3556);
  VN592_in5 <= VN_sign_in(3557) & VN_data_in(3557);
  VN593_in0 <= VN_sign_in(3558) & VN_data_in(3558);
  VN593_in1 <= VN_sign_in(3559) & VN_data_in(3559);
  VN593_in2 <= VN_sign_in(3560) & VN_data_in(3560);
  VN593_in3 <= VN_sign_in(3561) & VN_data_in(3561);
  VN593_in4 <= VN_sign_in(3562) & VN_data_in(3562);
  VN593_in5 <= VN_sign_in(3563) & VN_data_in(3563);
  VN594_in0 <= VN_sign_in(3564) & VN_data_in(3564);
  VN594_in1 <= VN_sign_in(3565) & VN_data_in(3565);
  VN594_in2 <= VN_sign_in(3566) & VN_data_in(3566);
  VN594_in3 <= VN_sign_in(3567) & VN_data_in(3567);
  VN594_in4 <= VN_sign_in(3568) & VN_data_in(3568);
  VN594_in5 <= VN_sign_in(3569) & VN_data_in(3569);
  VN595_in0 <= VN_sign_in(3570) & VN_data_in(3570);
  VN595_in1 <= VN_sign_in(3571) & VN_data_in(3571);
  VN595_in2 <= VN_sign_in(3572) & VN_data_in(3572);
  VN595_in3 <= VN_sign_in(3573) & VN_data_in(3573);
  VN595_in4 <= VN_sign_in(3574) & VN_data_in(3574);
  VN595_in5 <= VN_sign_in(3575) & VN_data_in(3575);
  VN596_in0 <= VN_sign_in(3576) & VN_data_in(3576);
  VN596_in1 <= VN_sign_in(3577) & VN_data_in(3577);
  VN596_in2 <= VN_sign_in(3578) & VN_data_in(3578);
  VN596_in3 <= VN_sign_in(3579) & VN_data_in(3579);
  VN596_in4 <= VN_sign_in(3580) & VN_data_in(3580);
  VN596_in5 <= VN_sign_in(3581) & VN_data_in(3581);
  VN597_in0 <= VN_sign_in(3582) & VN_data_in(3582);
  VN597_in1 <= VN_sign_in(3583) & VN_data_in(3583);
  VN597_in2 <= VN_sign_in(3584) & VN_data_in(3584);
  VN597_in3 <= VN_sign_in(3585) & VN_data_in(3585);
  VN597_in4 <= VN_sign_in(3586) & VN_data_in(3586);
  VN597_in5 <= VN_sign_in(3587) & VN_data_in(3587);
  VN598_in0 <= VN_sign_in(3588) & VN_data_in(3588);
  VN598_in1 <= VN_sign_in(3589) & VN_data_in(3589);
  VN598_in2 <= VN_sign_in(3590) & VN_data_in(3590);
  VN598_in3 <= VN_sign_in(3591) & VN_data_in(3591);
  VN598_in4 <= VN_sign_in(3592) & VN_data_in(3592);
  VN598_in5 <= VN_sign_in(3593) & VN_data_in(3593);
  VN599_in0 <= VN_sign_in(3594) & VN_data_in(3594);
  VN599_in1 <= VN_sign_in(3595) & VN_data_in(3595);
  VN599_in2 <= VN_sign_in(3596) & VN_data_in(3596);
  VN599_in3 <= VN_sign_in(3597) & VN_data_in(3597);
  VN599_in4 <= VN_sign_in(3598) & VN_data_in(3598);
  VN599_in5 <= VN_sign_in(3599) & VN_data_in(3599);
  VN600_in0 <= VN_sign_in(3600) & VN_data_in(3600);
  VN600_in1 <= VN_sign_in(3601) & VN_data_in(3601);
  VN600_in2 <= VN_sign_in(3602) & VN_data_in(3602);
  VN600_in3 <= VN_sign_in(3603) & VN_data_in(3603);
  VN600_in4 <= VN_sign_in(3604) & VN_data_in(3604);
  VN600_in5 <= VN_sign_in(3605) & VN_data_in(3605);
  VN601_in0 <= VN_sign_in(3606) & VN_data_in(3606);
  VN601_in1 <= VN_sign_in(3607) & VN_data_in(3607);
  VN601_in2 <= VN_sign_in(3608) & VN_data_in(3608);
  VN601_in3 <= VN_sign_in(3609) & VN_data_in(3609);
  VN601_in4 <= VN_sign_in(3610) & VN_data_in(3610);
  VN601_in5 <= VN_sign_in(3611) & VN_data_in(3611);
  VN602_in0 <= VN_sign_in(3612) & VN_data_in(3612);
  VN602_in1 <= VN_sign_in(3613) & VN_data_in(3613);
  VN602_in2 <= VN_sign_in(3614) & VN_data_in(3614);
  VN602_in3 <= VN_sign_in(3615) & VN_data_in(3615);
  VN602_in4 <= VN_sign_in(3616) & VN_data_in(3616);
  VN602_in5 <= VN_sign_in(3617) & VN_data_in(3617);
  VN603_in0 <= VN_sign_in(3618) & VN_data_in(3618);
  VN603_in1 <= VN_sign_in(3619) & VN_data_in(3619);
  VN603_in2 <= VN_sign_in(3620) & VN_data_in(3620);
  VN603_in3 <= VN_sign_in(3621) & VN_data_in(3621);
  VN603_in4 <= VN_sign_in(3622) & VN_data_in(3622);
  VN603_in5 <= VN_sign_in(3623) & VN_data_in(3623);
  VN604_in0 <= VN_sign_in(3624) & VN_data_in(3624);
  VN604_in1 <= VN_sign_in(3625) & VN_data_in(3625);
  VN604_in2 <= VN_sign_in(3626) & VN_data_in(3626);
  VN604_in3 <= VN_sign_in(3627) & VN_data_in(3627);
  VN604_in4 <= VN_sign_in(3628) & VN_data_in(3628);
  VN604_in5 <= VN_sign_in(3629) & VN_data_in(3629);
  VN605_in0 <= VN_sign_in(3630) & VN_data_in(3630);
  VN605_in1 <= VN_sign_in(3631) & VN_data_in(3631);
  VN605_in2 <= VN_sign_in(3632) & VN_data_in(3632);
  VN605_in3 <= VN_sign_in(3633) & VN_data_in(3633);
  VN605_in4 <= VN_sign_in(3634) & VN_data_in(3634);
  VN605_in5 <= VN_sign_in(3635) & VN_data_in(3635);
  VN606_in0 <= VN_sign_in(3636) & VN_data_in(3636);
  VN606_in1 <= VN_sign_in(3637) & VN_data_in(3637);
  VN606_in2 <= VN_sign_in(3638) & VN_data_in(3638);
  VN606_in3 <= VN_sign_in(3639) & VN_data_in(3639);
  VN606_in4 <= VN_sign_in(3640) & VN_data_in(3640);
  VN606_in5 <= VN_sign_in(3641) & VN_data_in(3641);
  VN607_in0 <= VN_sign_in(3642) & VN_data_in(3642);
  VN607_in1 <= VN_sign_in(3643) & VN_data_in(3643);
  VN607_in2 <= VN_sign_in(3644) & VN_data_in(3644);
  VN607_in3 <= VN_sign_in(3645) & VN_data_in(3645);
  VN607_in4 <= VN_sign_in(3646) & VN_data_in(3646);
  VN607_in5 <= VN_sign_in(3647) & VN_data_in(3647);
  VN608_in0 <= VN_sign_in(3648) & VN_data_in(3648);
  VN608_in1 <= VN_sign_in(3649) & VN_data_in(3649);
  VN608_in2 <= VN_sign_in(3650) & VN_data_in(3650);
  VN608_in3 <= VN_sign_in(3651) & VN_data_in(3651);
  VN608_in4 <= VN_sign_in(3652) & VN_data_in(3652);
  VN608_in5 <= VN_sign_in(3653) & VN_data_in(3653);
  VN609_in0 <= VN_sign_in(3654) & VN_data_in(3654);
  VN609_in1 <= VN_sign_in(3655) & VN_data_in(3655);
  VN609_in2 <= VN_sign_in(3656) & VN_data_in(3656);
  VN609_in3 <= VN_sign_in(3657) & VN_data_in(3657);
  VN609_in4 <= VN_sign_in(3658) & VN_data_in(3658);
  VN609_in5 <= VN_sign_in(3659) & VN_data_in(3659);
  VN610_in0 <= VN_sign_in(3660) & VN_data_in(3660);
  VN610_in1 <= VN_sign_in(3661) & VN_data_in(3661);
  VN610_in2 <= VN_sign_in(3662) & VN_data_in(3662);
  VN610_in3 <= VN_sign_in(3663) & VN_data_in(3663);
  VN610_in4 <= VN_sign_in(3664) & VN_data_in(3664);
  VN610_in5 <= VN_sign_in(3665) & VN_data_in(3665);
  VN611_in0 <= VN_sign_in(3666) & VN_data_in(3666);
  VN611_in1 <= VN_sign_in(3667) & VN_data_in(3667);
  VN611_in2 <= VN_sign_in(3668) & VN_data_in(3668);
  VN611_in3 <= VN_sign_in(3669) & VN_data_in(3669);
  VN611_in4 <= VN_sign_in(3670) & VN_data_in(3670);
  VN611_in5 <= VN_sign_in(3671) & VN_data_in(3671);
  VN612_in0 <= VN_sign_in(3672) & VN_data_in(3672);
  VN612_in1 <= VN_sign_in(3673) & VN_data_in(3673);
  VN612_in2 <= VN_sign_in(3674) & VN_data_in(3674);
  VN612_in3 <= VN_sign_in(3675) & VN_data_in(3675);
  VN612_in4 <= VN_sign_in(3676) & VN_data_in(3676);
  VN612_in5 <= VN_sign_in(3677) & VN_data_in(3677);
  VN613_in0 <= VN_sign_in(3678) & VN_data_in(3678);
  VN613_in1 <= VN_sign_in(3679) & VN_data_in(3679);
  VN613_in2 <= VN_sign_in(3680) & VN_data_in(3680);
  VN613_in3 <= VN_sign_in(3681) & VN_data_in(3681);
  VN613_in4 <= VN_sign_in(3682) & VN_data_in(3682);
  VN613_in5 <= VN_sign_in(3683) & VN_data_in(3683);
  VN614_in0 <= VN_sign_in(3684) & VN_data_in(3684);
  VN614_in1 <= VN_sign_in(3685) & VN_data_in(3685);
  VN614_in2 <= VN_sign_in(3686) & VN_data_in(3686);
  VN614_in3 <= VN_sign_in(3687) & VN_data_in(3687);
  VN614_in4 <= VN_sign_in(3688) & VN_data_in(3688);
  VN614_in5 <= VN_sign_in(3689) & VN_data_in(3689);
  VN615_in0 <= VN_sign_in(3690) & VN_data_in(3690);
  VN615_in1 <= VN_sign_in(3691) & VN_data_in(3691);
  VN615_in2 <= VN_sign_in(3692) & VN_data_in(3692);
  VN615_in3 <= VN_sign_in(3693) & VN_data_in(3693);
  VN615_in4 <= VN_sign_in(3694) & VN_data_in(3694);
  VN615_in5 <= VN_sign_in(3695) & VN_data_in(3695);
  VN616_in0 <= VN_sign_in(3696) & VN_data_in(3696);
  VN616_in1 <= VN_sign_in(3697) & VN_data_in(3697);
  VN616_in2 <= VN_sign_in(3698) & VN_data_in(3698);
  VN616_in3 <= VN_sign_in(3699) & VN_data_in(3699);
  VN616_in4 <= VN_sign_in(3700) & VN_data_in(3700);
  VN616_in5 <= VN_sign_in(3701) & VN_data_in(3701);
  VN617_in0 <= VN_sign_in(3702) & VN_data_in(3702);
  VN617_in1 <= VN_sign_in(3703) & VN_data_in(3703);
  VN617_in2 <= VN_sign_in(3704) & VN_data_in(3704);
  VN617_in3 <= VN_sign_in(3705) & VN_data_in(3705);
  VN617_in4 <= VN_sign_in(3706) & VN_data_in(3706);
  VN617_in5 <= VN_sign_in(3707) & VN_data_in(3707);
  VN618_in0 <= VN_sign_in(3708) & VN_data_in(3708);
  VN618_in1 <= VN_sign_in(3709) & VN_data_in(3709);
  VN618_in2 <= VN_sign_in(3710) & VN_data_in(3710);
  VN618_in3 <= VN_sign_in(3711) & VN_data_in(3711);
  VN618_in4 <= VN_sign_in(3712) & VN_data_in(3712);
  VN618_in5 <= VN_sign_in(3713) & VN_data_in(3713);
  VN619_in0 <= VN_sign_in(3714) & VN_data_in(3714);
  VN619_in1 <= VN_sign_in(3715) & VN_data_in(3715);
  VN619_in2 <= VN_sign_in(3716) & VN_data_in(3716);
  VN619_in3 <= VN_sign_in(3717) & VN_data_in(3717);
  VN619_in4 <= VN_sign_in(3718) & VN_data_in(3718);
  VN619_in5 <= VN_sign_in(3719) & VN_data_in(3719);
  VN620_in0 <= VN_sign_in(3720) & VN_data_in(3720);
  VN620_in1 <= VN_sign_in(3721) & VN_data_in(3721);
  VN620_in2 <= VN_sign_in(3722) & VN_data_in(3722);
  VN620_in3 <= VN_sign_in(3723) & VN_data_in(3723);
  VN620_in4 <= VN_sign_in(3724) & VN_data_in(3724);
  VN620_in5 <= VN_sign_in(3725) & VN_data_in(3725);
  VN621_in0 <= VN_sign_in(3726) & VN_data_in(3726);
  VN621_in1 <= VN_sign_in(3727) & VN_data_in(3727);
  VN621_in2 <= VN_sign_in(3728) & VN_data_in(3728);
  VN621_in3 <= VN_sign_in(3729) & VN_data_in(3729);
  VN621_in4 <= VN_sign_in(3730) & VN_data_in(3730);
  VN621_in5 <= VN_sign_in(3731) & VN_data_in(3731);
  VN622_in0 <= VN_sign_in(3732) & VN_data_in(3732);
  VN622_in1 <= VN_sign_in(3733) & VN_data_in(3733);
  VN622_in2 <= VN_sign_in(3734) & VN_data_in(3734);
  VN622_in3 <= VN_sign_in(3735) & VN_data_in(3735);
  VN622_in4 <= VN_sign_in(3736) & VN_data_in(3736);
  VN622_in5 <= VN_sign_in(3737) & VN_data_in(3737);
  VN623_in0 <= VN_sign_in(3738) & VN_data_in(3738);
  VN623_in1 <= VN_sign_in(3739) & VN_data_in(3739);
  VN623_in2 <= VN_sign_in(3740) & VN_data_in(3740);
  VN623_in3 <= VN_sign_in(3741) & VN_data_in(3741);
  VN623_in4 <= VN_sign_in(3742) & VN_data_in(3742);
  VN623_in5 <= VN_sign_in(3743) & VN_data_in(3743);
  VN624_in0 <= VN_sign_in(3744) & VN_data_in(3744);
  VN624_in1 <= VN_sign_in(3745) & VN_data_in(3745);
  VN624_in2 <= VN_sign_in(3746) & VN_data_in(3746);
  VN624_in3 <= VN_sign_in(3747) & VN_data_in(3747);
  VN624_in4 <= VN_sign_in(3748) & VN_data_in(3748);
  VN624_in5 <= VN_sign_in(3749) & VN_data_in(3749);
  VN625_in0 <= VN_sign_in(3750) & VN_data_in(3750);
  VN625_in1 <= VN_sign_in(3751) & VN_data_in(3751);
  VN625_in2 <= VN_sign_in(3752) & VN_data_in(3752);
  VN625_in3 <= VN_sign_in(3753) & VN_data_in(3753);
  VN625_in4 <= VN_sign_in(3754) & VN_data_in(3754);
  VN625_in5 <= VN_sign_in(3755) & VN_data_in(3755);
  VN626_in0 <= VN_sign_in(3756) & VN_data_in(3756);
  VN626_in1 <= VN_sign_in(3757) & VN_data_in(3757);
  VN626_in2 <= VN_sign_in(3758) & VN_data_in(3758);
  VN626_in3 <= VN_sign_in(3759) & VN_data_in(3759);
  VN626_in4 <= VN_sign_in(3760) & VN_data_in(3760);
  VN626_in5 <= VN_sign_in(3761) & VN_data_in(3761);
  VN627_in0 <= VN_sign_in(3762) & VN_data_in(3762);
  VN627_in1 <= VN_sign_in(3763) & VN_data_in(3763);
  VN627_in2 <= VN_sign_in(3764) & VN_data_in(3764);
  VN627_in3 <= VN_sign_in(3765) & VN_data_in(3765);
  VN627_in4 <= VN_sign_in(3766) & VN_data_in(3766);
  VN627_in5 <= VN_sign_in(3767) & VN_data_in(3767);
  VN628_in0 <= VN_sign_in(3768) & VN_data_in(3768);
  VN628_in1 <= VN_sign_in(3769) & VN_data_in(3769);
  VN628_in2 <= VN_sign_in(3770) & VN_data_in(3770);
  VN628_in3 <= VN_sign_in(3771) & VN_data_in(3771);
  VN628_in4 <= VN_sign_in(3772) & VN_data_in(3772);
  VN628_in5 <= VN_sign_in(3773) & VN_data_in(3773);
  VN629_in0 <= VN_sign_in(3774) & VN_data_in(3774);
  VN629_in1 <= VN_sign_in(3775) & VN_data_in(3775);
  VN629_in2 <= VN_sign_in(3776) & VN_data_in(3776);
  VN629_in3 <= VN_sign_in(3777) & VN_data_in(3777);
  VN629_in4 <= VN_sign_in(3778) & VN_data_in(3778);
  VN629_in5 <= VN_sign_in(3779) & VN_data_in(3779);
  VN630_in0 <= VN_sign_in(3780) & VN_data_in(3780);
  VN630_in1 <= VN_sign_in(3781) & VN_data_in(3781);
  VN630_in2 <= VN_sign_in(3782) & VN_data_in(3782);
  VN630_in3 <= VN_sign_in(3783) & VN_data_in(3783);
  VN630_in4 <= VN_sign_in(3784) & VN_data_in(3784);
  VN630_in5 <= VN_sign_in(3785) & VN_data_in(3785);
  VN631_in0 <= VN_sign_in(3786) & VN_data_in(3786);
  VN631_in1 <= VN_sign_in(3787) & VN_data_in(3787);
  VN631_in2 <= VN_sign_in(3788) & VN_data_in(3788);
  VN631_in3 <= VN_sign_in(3789) & VN_data_in(3789);
  VN631_in4 <= VN_sign_in(3790) & VN_data_in(3790);
  VN631_in5 <= VN_sign_in(3791) & VN_data_in(3791);
  VN632_in0 <= VN_sign_in(3792) & VN_data_in(3792);
  VN632_in1 <= VN_sign_in(3793) & VN_data_in(3793);
  VN632_in2 <= VN_sign_in(3794) & VN_data_in(3794);
  VN632_in3 <= VN_sign_in(3795) & VN_data_in(3795);
  VN632_in4 <= VN_sign_in(3796) & VN_data_in(3796);
  VN632_in5 <= VN_sign_in(3797) & VN_data_in(3797);
  VN633_in0 <= VN_sign_in(3798) & VN_data_in(3798);
  VN633_in1 <= VN_sign_in(3799) & VN_data_in(3799);
  VN633_in2 <= VN_sign_in(3800) & VN_data_in(3800);
  VN633_in3 <= VN_sign_in(3801) & VN_data_in(3801);
  VN633_in4 <= VN_sign_in(3802) & VN_data_in(3802);
  VN633_in5 <= VN_sign_in(3803) & VN_data_in(3803);
  VN634_in0 <= VN_sign_in(3804) & VN_data_in(3804);
  VN634_in1 <= VN_sign_in(3805) & VN_data_in(3805);
  VN634_in2 <= VN_sign_in(3806) & VN_data_in(3806);
  VN634_in3 <= VN_sign_in(3807) & VN_data_in(3807);
  VN634_in4 <= VN_sign_in(3808) & VN_data_in(3808);
  VN634_in5 <= VN_sign_in(3809) & VN_data_in(3809);
  VN635_in0 <= VN_sign_in(3810) & VN_data_in(3810);
  VN635_in1 <= VN_sign_in(3811) & VN_data_in(3811);
  VN635_in2 <= VN_sign_in(3812) & VN_data_in(3812);
  VN635_in3 <= VN_sign_in(3813) & VN_data_in(3813);
  VN635_in4 <= VN_sign_in(3814) & VN_data_in(3814);
  VN635_in5 <= VN_sign_in(3815) & VN_data_in(3815);
  VN636_in0 <= VN_sign_in(3816) & VN_data_in(3816);
  VN636_in1 <= VN_sign_in(3817) & VN_data_in(3817);
  VN636_in2 <= VN_sign_in(3818) & VN_data_in(3818);
  VN636_in3 <= VN_sign_in(3819) & VN_data_in(3819);
  VN636_in4 <= VN_sign_in(3820) & VN_data_in(3820);
  VN636_in5 <= VN_sign_in(3821) & VN_data_in(3821);
  VN637_in0 <= VN_sign_in(3822) & VN_data_in(3822);
  VN637_in1 <= VN_sign_in(3823) & VN_data_in(3823);
  VN637_in2 <= VN_sign_in(3824) & VN_data_in(3824);
  VN637_in3 <= VN_sign_in(3825) & VN_data_in(3825);
  VN637_in4 <= VN_sign_in(3826) & VN_data_in(3826);
  VN637_in5 <= VN_sign_in(3827) & VN_data_in(3827);
  VN638_in0 <= VN_sign_in(3828) & VN_data_in(3828);
  VN638_in1 <= VN_sign_in(3829) & VN_data_in(3829);
  VN638_in2 <= VN_sign_in(3830) & VN_data_in(3830);
  VN638_in3 <= VN_sign_in(3831) & VN_data_in(3831);
  VN638_in4 <= VN_sign_in(3832) & VN_data_in(3832);
  VN638_in5 <= VN_sign_in(3833) & VN_data_in(3833);
  VN639_in0 <= VN_sign_in(3834) & VN_data_in(3834);
  VN639_in1 <= VN_sign_in(3835) & VN_data_in(3835);
  VN639_in2 <= VN_sign_in(3836) & VN_data_in(3836);
  VN639_in3 <= VN_sign_in(3837) & VN_data_in(3837);
  VN639_in4 <= VN_sign_in(3838) & VN_data_in(3838);
  VN639_in5 <= VN_sign_in(3839) & VN_data_in(3839);
  VN640_in0 <= VN_sign_in(3840) & VN_data_in(3840);
  VN640_in1 <= VN_sign_in(3841) & VN_data_in(3841);
  VN640_in2 <= VN_sign_in(3842) & VN_data_in(3842);
  VN640_in3 <= VN_sign_in(3843) & VN_data_in(3843);
  VN640_in4 <= VN_sign_in(3844) & VN_data_in(3844);
  VN640_in5 <= VN_sign_in(3845) & VN_data_in(3845);
  VN641_in0 <= VN_sign_in(3846) & VN_data_in(3846);
  VN641_in1 <= VN_sign_in(3847) & VN_data_in(3847);
  VN641_in2 <= VN_sign_in(3848) & VN_data_in(3848);
  VN641_in3 <= VN_sign_in(3849) & VN_data_in(3849);
  VN641_in4 <= VN_sign_in(3850) & VN_data_in(3850);
  VN641_in5 <= VN_sign_in(3851) & VN_data_in(3851);
  VN642_in0 <= VN_sign_in(3852) & VN_data_in(3852);
  VN642_in1 <= VN_sign_in(3853) & VN_data_in(3853);
  VN642_in2 <= VN_sign_in(3854) & VN_data_in(3854);
  VN642_in3 <= VN_sign_in(3855) & VN_data_in(3855);
  VN642_in4 <= VN_sign_in(3856) & VN_data_in(3856);
  VN642_in5 <= VN_sign_in(3857) & VN_data_in(3857);
  VN643_in0 <= VN_sign_in(3858) & VN_data_in(3858);
  VN643_in1 <= VN_sign_in(3859) & VN_data_in(3859);
  VN643_in2 <= VN_sign_in(3860) & VN_data_in(3860);
  VN643_in3 <= VN_sign_in(3861) & VN_data_in(3861);
  VN643_in4 <= VN_sign_in(3862) & VN_data_in(3862);
  VN643_in5 <= VN_sign_in(3863) & VN_data_in(3863);
  VN644_in0 <= VN_sign_in(3864) & VN_data_in(3864);
  VN644_in1 <= VN_sign_in(3865) & VN_data_in(3865);
  VN644_in2 <= VN_sign_in(3866) & VN_data_in(3866);
  VN644_in3 <= VN_sign_in(3867) & VN_data_in(3867);
  VN644_in4 <= VN_sign_in(3868) & VN_data_in(3868);
  VN644_in5 <= VN_sign_in(3869) & VN_data_in(3869);
  VN645_in0 <= VN_sign_in(3870) & VN_data_in(3870);
  VN645_in1 <= VN_sign_in(3871) & VN_data_in(3871);
  VN645_in2 <= VN_sign_in(3872) & VN_data_in(3872);
  VN645_in3 <= VN_sign_in(3873) & VN_data_in(3873);
  VN645_in4 <= VN_sign_in(3874) & VN_data_in(3874);
  VN645_in5 <= VN_sign_in(3875) & VN_data_in(3875);
  VN646_in0 <= VN_sign_in(3876) & VN_data_in(3876);
  VN646_in1 <= VN_sign_in(3877) & VN_data_in(3877);
  VN646_in2 <= VN_sign_in(3878) & VN_data_in(3878);
  VN646_in3 <= VN_sign_in(3879) & VN_data_in(3879);
  VN646_in4 <= VN_sign_in(3880) & VN_data_in(3880);
  VN646_in5 <= VN_sign_in(3881) & VN_data_in(3881);
  VN647_in0 <= VN_sign_in(3882) & VN_data_in(3882);
  VN647_in1 <= VN_sign_in(3883) & VN_data_in(3883);
  VN647_in2 <= VN_sign_in(3884) & VN_data_in(3884);
  VN647_in3 <= VN_sign_in(3885) & VN_data_in(3885);
  VN647_in4 <= VN_sign_in(3886) & VN_data_in(3886);
  VN647_in5 <= VN_sign_in(3887) & VN_data_in(3887);
  VN648_in0 <= VN_sign_in(3888) & VN_data_in(3888);
  VN648_in1 <= VN_sign_in(3889) & VN_data_in(3889);
  VN648_in2 <= VN_sign_in(3890) & VN_data_in(3890);
  VN648_in3 <= VN_sign_in(3891) & VN_data_in(3891);
  VN648_in4 <= VN_sign_in(3892) & VN_data_in(3892);
  VN648_in5 <= VN_sign_in(3893) & VN_data_in(3893);
  VN649_in0 <= VN_sign_in(3894) & VN_data_in(3894);
  VN649_in1 <= VN_sign_in(3895) & VN_data_in(3895);
  VN649_in2 <= VN_sign_in(3896) & VN_data_in(3896);
  VN649_in3 <= VN_sign_in(3897) & VN_data_in(3897);
  VN649_in4 <= VN_sign_in(3898) & VN_data_in(3898);
  VN649_in5 <= VN_sign_in(3899) & VN_data_in(3899);
  VN650_in0 <= VN_sign_in(3900) & VN_data_in(3900);
  VN650_in1 <= VN_sign_in(3901) & VN_data_in(3901);
  VN650_in2 <= VN_sign_in(3902) & VN_data_in(3902);
  VN650_in3 <= VN_sign_in(3903) & VN_data_in(3903);
  VN650_in4 <= VN_sign_in(3904) & VN_data_in(3904);
  VN650_in5 <= VN_sign_in(3905) & VN_data_in(3905);
  VN651_in0 <= VN_sign_in(3906) & VN_data_in(3906);
  VN651_in1 <= VN_sign_in(3907) & VN_data_in(3907);
  VN651_in2 <= VN_sign_in(3908) & VN_data_in(3908);
  VN651_in3 <= VN_sign_in(3909) & VN_data_in(3909);
  VN651_in4 <= VN_sign_in(3910) & VN_data_in(3910);
  VN651_in5 <= VN_sign_in(3911) & VN_data_in(3911);
  VN652_in0 <= VN_sign_in(3912) & VN_data_in(3912);
  VN652_in1 <= VN_sign_in(3913) & VN_data_in(3913);
  VN652_in2 <= VN_sign_in(3914) & VN_data_in(3914);
  VN652_in3 <= VN_sign_in(3915) & VN_data_in(3915);
  VN652_in4 <= VN_sign_in(3916) & VN_data_in(3916);
  VN652_in5 <= VN_sign_in(3917) & VN_data_in(3917);
  VN653_in0 <= VN_sign_in(3918) & VN_data_in(3918);
  VN653_in1 <= VN_sign_in(3919) & VN_data_in(3919);
  VN653_in2 <= VN_sign_in(3920) & VN_data_in(3920);
  VN653_in3 <= VN_sign_in(3921) & VN_data_in(3921);
  VN653_in4 <= VN_sign_in(3922) & VN_data_in(3922);
  VN653_in5 <= VN_sign_in(3923) & VN_data_in(3923);
  VN654_in0 <= VN_sign_in(3924) & VN_data_in(3924);
  VN654_in1 <= VN_sign_in(3925) & VN_data_in(3925);
  VN654_in2 <= VN_sign_in(3926) & VN_data_in(3926);
  VN654_in3 <= VN_sign_in(3927) & VN_data_in(3927);
  VN654_in4 <= VN_sign_in(3928) & VN_data_in(3928);
  VN654_in5 <= VN_sign_in(3929) & VN_data_in(3929);
  VN655_in0 <= VN_sign_in(3930) & VN_data_in(3930);
  VN655_in1 <= VN_sign_in(3931) & VN_data_in(3931);
  VN655_in2 <= VN_sign_in(3932) & VN_data_in(3932);
  VN655_in3 <= VN_sign_in(3933) & VN_data_in(3933);
  VN655_in4 <= VN_sign_in(3934) & VN_data_in(3934);
  VN655_in5 <= VN_sign_in(3935) & VN_data_in(3935);
  VN656_in0 <= VN_sign_in(3936) & VN_data_in(3936);
  VN656_in1 <= VN_sign_in(3937) & VN_data_in(3937);
  VN656_in2 <= VN_sign_in(3938) & VN_data_in(3938);
  VN656_in3 <= VN_sign_in(3939) & VN_data_in(3939);
  VN656_in4 <= VN_sign_in(3940) & VN_data_in(3940);
  VN656_in5 <= VN_sign_in(3941) & VN_data_in(3941);
  VN657_in0 <= VN_sign_in(3942) & VN_data_in(3942);
  VN657_in1 <= VN_sign_in(3943) & VN_data_in(3943);
  VN657_in2 <= VN_sign_in(3944) & VN_data_in(3944);
  VN657_in3 <= VN_sign_in(3945) & VN_data_in(3945);
  VN657_in4 <= VN_sign_in(3946) & VN_data_in(3946);
  VN657_in5 <= VN_sign_in(3947) & VN_data_in(3947);
  VN658_in0 <= VN_sign_in(3948) & VN_data_in(3948);
  VN658_in1 <= VN_sign_in(3949) & VN_data_in(3949);
  VN658_in2 <= VN_sign_in(3950) & VN_data_in(3950);
  VN658_in3 <= VN_sign_in(3951) & VN_data_in(3951);
  VN658_in4 <= VN_sign_in(3952) & VN_data_in(3952);
  VN658_in5 <= VN_sign_in(3953) & VN_data_in(3953);
  VN659_in0 <= VN_sign_in(3954) & VN_data_in(3954);
  VN659_in1 <= VN_sign_in(3955) & VN_data_in(3955);
  VN659_in2 <= VN_sign_in(3956) & VN_data_in(3956);
  VN659_in3 <= VN_sign_in(3957) & VN_data_in(3957);
  VN659_in4 <= VN_sign_in(3958) & VN_data_in(3958);
  VN659_in5 <= VN_sign_in(3959) & VN_data_in(3959);
  VN660_in0 <= VN_sign_in(3960) & VN_data_in(3960);
  VN660_in1 <= VN_sign_in(3961) & VN_data_in(3961);
  VN660_in2 <= VN_sign_in(3962) & VN_data_in(3962);
  VN660_in3 <= VN_sign_in(3963) & VN_data_in(3963);
  VN660_in4 <= VN_sign_in(3964) & VN_data_in(3964);
  VN660_in5 <= VN_sign_in(3965) & VN_data_in(3965);
  VN661_in0 <= VN_sign_in(3966) & VN_data_in(3966);
  VN661_in1 <= VN_sign_in(3967) & VN_data_in(3967);
  VN661_in2 <= VN_sign_in(3968) & VN_data_in(3968);
  VN661_in3 <= VN_sign_in(3969) & VN_data_in(3969);
  VN661_in4 <= VN_sign_in(3970) & VN_data_in(3970);
  VN661_in5 <= VN_sign_in(3971) & VN_data_in(3971);
  VN662_in0 <= VN_sign_in(3972) & VN_data_in(3972);
  VN662_in1 <= VN_sign_in(3973) & VN_data_in(3973);
  VN662_in2 <= VN_sign_in(3974) & VN_data_in(3974);
  VN662_in3 <= VN_sign_in(3975) & VN_data_in(3975);
  VN662_in4 <= VN_sign_in(3976) & VN_data_in(3976);
  VN662_in5 <= VN_sign_in(3977) & VN_data_in(3977);
  VN663_in0 <= VN_sign_in(3978) & VN_data_in(3978);
  VN663_in1 <= VN_sign_in(3979) & VN_data_in(3979);
  VN663_in2 <= VN_sign_in(3980) & VN_data_in(3980);
  VN663_in3 <= VN_sign_in(3981) & VN_data_in(3981);
  VN663_in4 <= VN_sign_in(3982) & VN_data_in(3982);
  VN663_in5 <= VN_sign_in(3983) & VN_data_in(3983);
  VN664_in0 <= VN_sign_in(3984) & VN_data_in(3984);
  VN664_in1 <= VN_sign_in(3985) & VN_data_in(3985);
  VN664_in2 <= VN_sign_in(3986) & VN_data_in(3986);
  VN664_in3 <= VN_sign_in(3987) & VN_data_in(3987);
  VN664_in4 <= VN_sign_in(3988) & VN_data_in(3988);
  VN664_in5 <= VN_sign_in(3989) & VN_data_in(3989);
  VN665_in0 <= VN_sign_in(3990) & VN_data_in(3990);
  VN665_in1 <= VN_sign_in(3991) & VN_data_in(3991);
  VN665_in2 <= VN_sign_in(3992) & VN_data_in(3992);
  VN665_in3 <= VN_sign_in(3993) & VN_data_in(3993);
  VN665_in4 <= VN_sign_in(3994) & VN_data_in(3994);
  VN665_in5 <= VN_sign_in(3995) & VN_data_in(3995);
  VN666_in0 <= VN_sign_in(3996) & VN_data_in(3996);
  VN666_in1 <= VN_sign_in(3997) & VN_data_in(3997);
  VN666_in2 <= VN_sign_in(3998) & VN_data_in(3998);
  VN666_in3 <= VN_sign_in(3999) & VN_data_in(3999);
  VN666_in4 <= VN_sign_in(4000) & VN_data_in(4000);
  VN666_in5 <= VN_sign_in(4001) & VN_data_in(4001);
  VN667_in0 <= VN_sign_in(4002) & VN_data_in(4002);
  VN667_in1 <= VN_sign_in(4003) & VN_data_in(4003);
  VN667_in2 <= VN_sign_in(4004) & VN_data_in(4004);
  VN667_in3 <= VN_sign_in(4005) & VN_data_in(4005);
  VN667_in4 <= VN_sign_in(4006) & VN_data_in(4006);
  VN667_in5 <= VN_sign_in(4007) & VN_data_in(4007);
  VN668_in0 <= VN_sign_in(4008) & VN_data_in(4008);
  VN668_in1 <= VN_sign_in(4009) & VN_data_in(4009);
  VN668_in2 <= VN_sign_in(4010) & VN_data_in(4010);
  VN668_in3 <= VN_sign_in(4011) & VN_data_in(4011);
  VN668_in4 <= VN_sign_in(4012) & VN_data_in(4012);
  VN668_in5 <= VN_sign_in(4013) & VN_data_in(4013);
  VN669_in0 <= VN_sign_in(4014) & VN_data_in(4014);
  VN669_in1 <= VN_sign_in(4015) & VN_data_in(4015);
  VN669_in2 <= VN_sign_in(4016) & VN_data_in(4016);
  VN669_in3 <= VN_sign_in(4017) & VN_data_in(4017);
  VN669_in4 <= VN_sign_in(4018) & VN_data_in(4018);
  VN669_in5 <= VN_sign_in(4019) & VN_data_in(4019);
  VN670_in0 <= VN_sign_in(4020) & VN_data_in(4020);
  VN670_in1 <= VN_sign_in(4021) & VN_data_in(4021);
  VN670_in2 <= VN_sign_in(4022) & VN_data_in(4022);
  VN670_in3 <= VN_sign_in(4023) & VN_data_in(4023);
  VN670_in4 <= VN_sign_in(4024) & VN_data_in(4024);
  VN670_in5 <= VN_sign_in(4025) & VN_data_in(4025);
  VN671_in0 <= VN_sign_in(4026) & VN_data_in(4026);
  VN671_in1 <= VN_sign_in(4027) & VN_data_in(4027);
  VN671_in2 <= VN_sign_in(4028) & VN_data_in(4028);
  VN671_in3 <= VN_sign_in(4029) & VN_data_in(4029);
  VN671_in4 <= VN_sign_in(4030) & VN_data_in(4030);
  VN671_in5 <= VN_sign_in(4031) & VN_data_in(4031);
  VN672_in0 <= VN_sign_in(4032) & VN_data_in(4032);
  VN672_in1 <= VN_sign_in(4033) & VN_data_in(4033);
  VN672_in2 <= VN_sign_in(4034) & VN_data_in(4034);
  VN672_in3 <= VN_sign_in(4035) & VN_data_in(4035);
  VN672_in4 <= VN_sign_in(4036) & VN_data_in(4036);
  VN672_in5 <= VN_sign_in(4037) & VN_data_in(4037);
  VN673_in0 <= VN_sign_in(4038) & VN_data_in(4038);
  VN673_in1 <= VN_sign_in(4039) & VN_data_in(4039);
  VN673_in2 <= VN_sign_in(4040) & VN_data_in(4040);
  VN673_in3 <= VN_sign_in(4041) & VN_data_in(4041);
  VN673_in4 <= VN_sign_in(4042) & VN_data_in(4042);
  VN673_in5 <= VN_sign_in(4043) & VN_data_in(4043);
  VN674_in0 <= VN_sign_in(4044) & VN_data_in(4044);
  VN674_in1 <= VN_sign_in(4045) & VN_data_in(4045);
  VN674_in2 <= VN_sign_in(4046) & VN_data_in(4046);
  VN674_in3 <= VN_sign_in(4047) & VN_data_in(4047);
  VN674_in4 <= VN_sign_in(4048) & VN_data_in(4048);
  VN674_in5 <= VN_sign_in(4049) & VN_data_in(4049);
  VN675_in0 <= VN_sign_in(4050) & VN_data_in(4050);
  VN675_in1 <= VN_sign_in(4051) & VN_data_in(4051);
  VN675_in2 <= VN_sign_in(4052) & VN_data_in(4052);
  VN675_in3 <= VN_sign_in(4053) & VN_data_in(4053);
  VN675_in4 <= VN_sign_in(4054) & VN_data_in(4054);
  VN675_in5 <= VN_sign_in(4055) & VN_data_in(4055);
  VN676_in0 <= VN_sign_in(4056) & VN_data_in(4056);
  VN676_in1 <= VN_sign_in(4057) & VN_data_in(4057);
  VN676_in2 <= VN_sign_in(4058) & VN_data_in(4058);
  VN676_in3 <= VN_sign_in(4059) & VN_data_in(4059);
  VN676_in4 <= VN_sign_in(4060) & VN_data_in(4060);
  VN676_in5 <= VN_sign_in(4061) & VN_data_in(4061);
  VN677_in0 <= VN_sign_in(4062) & VN_data_in(4062);
  VN677_in1 <= VN_sign_in(4063) & VN_data_in(4063);
  VN677_in2 <= VN_sign_in(4064) & VN_data_in(4064);
  VN677_in3 <= VN_sign_in(4065) & VN_data_in(4065);
  VN677_in4 <= VN_sign_in(4066) & VN_data_in(4066);
  VN677_in5 <= VN_sign_in(4067) & VN_data_in(4067);
  VN678_in0 <= VN_sign_in(4068) & VN_data_in(4068);
  VN678_in1 <= VN_sign_in(4069) & VN_data_in(4069);
  VN678_in2 <= VN_sign_in(4070) & VN_data_in(4070);
  VN678_in3 <= VN_sign_in(4071) & VN_data_in(4071);
  VN678_in4 <= VN_sign_in(4072) & VN_data_in(4072);
  VN678_in5 <= VN_sign_in(4073) & VN_data_in(4073);
  VN679_in0 <= VN_sign_in(4074) & VN_data_in(4074);
  VN679_in1 <= VN_sign_in(4075) & VN_data_in(4075);
  VN679_in2 <= VN_sign_in(4076) & VN_data_in(4076);
  VN679_in3 <= VN_sign_in(4077) & VN_data_in(4077);
  VN679_in4 <= VN_sign_in(4078) & VN_data_in(4078);
  VN679_in5 <= VN_sign_in(4079) & VN_data_in(4079);
  VN680_in0 <= VN_sign_in(4080) & VN_data_in(4080);
  VN680_in1 <= VN_sign_in(4081) & VN_data_in(4081);
  VN680_in2 <= VN_sign_in(4082) & VN_data_in(4082);
  VN680_in3 <= VN_sign_in(4083) & VN_data_in(4083);
  VN680_in4 <= VN_sign_in(4084) & VN_data_in(4084);
  VN680_in5 <= VN_sign_in(4085) & VN_data_in(4085);
  VN681_in0 <= VN_sign_in(4086) & VN_data_in(4086);
  VN681_in1 <= VN_sign_in(4087) & VN_data_in(4087);
  VN681_in2 <= VN_sign_in(4088) & VN_data_in(4088);
  VN681_in3 <= VN_sign_in(4089) & VN_data_in(4089);
  VN681_in4 <= VN_sign_in(4090) & VN_data_in(4090);
  VN681_in5 <= VN_sign_in(4091) & VN_data_in(4091);
  VN682_in0 <= VN_sign_in(4092) & VN_data_in(4092);
  VN682_in1 <= VN_sign_in(4093) & VN_data_in(4093);
  VN682_in2 <= VN_sign_in(4094) & VN_data_in(4094);
  VN682_in3 <= VN_sign_in(4095) & VN_data_in(4095);
  VN682_in4 <= VN_sign_in(4096) & VN_data_in(4096);
  VN682_in5 <= VN_sign_in(4097) & VN_data_in(4097);
  VN683_in0 <= VN_sign_in(4098) & VN_data_in(4098);
  VN683_in1 <= VN_sign_in(4099) & VN_data_in(4099);
  VN683_in2 <= VN_sign_in(4100) & VN_data_in(4100);
  VN683_in3 <= VN_sign_in(4101) & VN_data_in(4101);
  VN683_in4 <= VN_sign_in(4102) & VN_data_in(4102);
  VN683_in5 <= VN_sign_in(4103) & VN_data_in(4103);
  VN684_in0 <= VN_sign_in(4104) & VN_data_in(4104);
  VN684_in1 <= VN_sign_in(4105) & VN_data_in(4105);
  VN684_in2 <= VN_sign_in(4106) & VN_data_in(4106);
  VN684_in3 <= VN_sign_in(4107) & VN_data_in(4107);
  VN684_in4 <= VN_sign_in(4108) & VN_data_in(4108);
  VN684_in5 <= VN_sign_in(4109) & VN_data_in(4109);
  VN685_in0 <= VN_sign_in(4110) & VN_data_in(4110);
  VN685_in1 <= VN_sign_in(4111) & VN_data_in(4111);
  VN685_in2 <= VN_sign_in(4112) & VN_data_in(4112);
  VN685_in3 <= VN_sign_in(4113) & VN_data_in(4113);
  VN685_in4 <= VN_sign_in(4114) & VN_data_in(4114);
  VN685_in5 <= VN_sign_in(4115) & VN_data_in(4115);
  VN686_in0 <= VN_sign_in(4116) & VN_data_in(4116);
  VN686_in1 <= VN_sign_in(4117) & VN_data_in(4117);
  VN686_in2 <= VN_sign_in(4118) & VN_data_in(4118);
  VN686_in3 <= VN_sign_in(4119) & VN_data_in(4119);
  VN686_in4 <= VN_sign_in(4120) & VN_data_in(4120);
  VN686_in5 <= VN_sign_in(4121) & VN_data_in(4121);
  VN687_in0 <= VN_sign_in(4122) & VN_data_in(4122);
  VN687_in1 <= VN_sign_in(4123) & VN_data_in(4123);
  VN687_in2 <= VN_sign_in(4124) & VN_data_in(4124);
  VN687_in3 <= VN_sign_in(4125) & VN_data_in(4125);
  VN687_in4 <= VN_sign_in(4126) & VN_data_in(4126);
  VN687_in5 <= VN_sign_in(4127) & VN_data_in(4127);
  VN688_in0 <= VN_sign_in(4128) & VN_data_in(4128);
  VN688_in1 <= VN_sign_in(4129) & VN_data_in(4129);
  VN688_in2 <= VN_sign_in(4130) & VN_data_in(4130);
  VN688_in3 <= VN_sign_in(4131) & VN_data_in(4131);
  VN688_in4 <= VN_sign_in(4132) & VN_data_in(4132);
  VN688_in5 <= VN_sign_in(4133) & VN_data_in(4133);
  VN689_in0 <= VN_sign_in(4134) & VN_data_in(4134);
  VN689_in1 <= VN_sign_in(4135) & VN_data_in(4135);
  VN689_in2 <= VN_sign_in(4136) & VN_data_in(4136);
  VN689_in3 <= VN_sign_in(4137) & VN_data_in(4137);
  VN689_in4 <= VN_sign_in(4138) & VN_data_in(4138);
  VN689_in5 <= VN_sign_in(4139) & VN_data_in(4139);
  VN690_in0 <= VN_sign_in(4140) & VN_data_in(4140);
  VN690_in1 <= VN_sign_in(4141) & VN_data_in(4141);
  VN690_in2 <= VN_sign_in(4142) & VN_data_in(4142);
  VN690_in3 <= VN_sign_in(4143) & VN_data_in(4143);
  VN690_in4 <= VN_sign_in(4144) & VN_data_in(4144);
  VN690_in5 <= VN_sign_in(4145) & VN_data_in(4145);
  VN691_in0 <= VN_sign_in(4146) & VN_data_in(4146);
  VN691_in1 <= VN_sign_in(4147) & VN_data_in(4147);
  VN691_in2 <= VN_sign_in(4148) & VN_data_in(4148);
  VN691_in3 <= VN_sign_in(4149) & VN_data_in(4149);
  VN691_in4 <= VN_sign_in(4150) & VN_data_in(4150);
  VN691_in5 <= VN_sign_in(4151) & VN_data_in(4151);
  VN692_in0 <= VN_sign_in(4152) & VN_data_in(4152);
  VN692_in1 <= VN_sign_in(4153) & VN_data_in(4153);
  VN692_in2 <= VN_sign_in(4154) & VN_data_in(4154);
  VN692_in3 <= VN_sign_in(4155) & VN_data_in(4155);
  VN692_in4 <= VN_sign_in(4156) & VN_data_in(4156);
  VN692_in5 <= VN_sign_in(4157) & VN_data_in(4157);
  VN693_in0 <= VN_sign_in(4158) & VN_data_in(4158);
  VN693_in1 <= VN_sign_in(4159) & VN_data_in(4159);
  VN693_in2 <= VN_sign_in(4160) & VN_data_in(4160);
  VN693_in3 <= VN_sign_in(4161) & VN_data_in(4161);
  VN693_in4 <= VN_sign_in(4162) & VN_data_in(4162);
  VN693_in5 <= VN_sign_in(4163) & VN_data_in(4163);
  VN694_in0 <= VN_sign_in(4164) & VN_data_in(4164);
  VN694_in1 <= VN_sign_in(4165) & VN_data_in(4165);
  VN694_in2 <= VN_sign_in(4166) & VN_data_in(4166);
  VN694_in3 <= VN_sign_in(4167) & VN_data_in(4167);
  VN694_in4 <= VN_sign_in(4168) & VN_data_in(4168);
  VN694_in5 <= VN_sign_in(4169) & VN_data_in(4169);
  VN695_in0 <= VN_sign_in(4170) & VN_data_in(4170);
  VN695_in1 <= VN_sign_in(4171) & VN_data_in(4171);
  VN695_in2 <= VN_sign_in(4172) & VN_data_in(4172);
  VN695_in3 <= VN_sign_in(4173) & VN_data_in(4173);
  VN695_in4 <= VN_sign_in(4174) & VN_data_in(4174);
  VN695_in5 <= VN_sign_in(4175) & VN_data_in(4175);
  VN696_in0 <= VN_sign_in(4176) & VN_data_in(4176);
  VN696_in1 <= VN_sign_in(4177) & VN_data_in(4177);
  VN696_in2 <= VN_sign_in(4178) & VN_data_in(4178);
  VN696_in3 <= VN_sign_in(4179) & VN_data_in(4179);
  VN696_in4 <= VN_sign_in(4180) & VN_data_in(4180);
  VN696_in5 <= VN_sign_in(4181) & VN_data_in(4181);
  VN697_in0 <= VN_sign_in(4182) & VN_data_in(4182);
  VN697_in1 <= VN_sign_in(4183) & VN_data_in(4183);
  VN697_in2 <= VN_sign_in(4184) & VN_data_in(4184);
  VN697_in3 <= VN_sign_in(4185) & VN_data_in(4185);
  VN697_in4 <= VN_sign_in(4186) & VN_data_in(4186);
  VN697_in5 <= VN_sign_in(4187) & VN_data_in(4187);
  VN698_in0 <= VN_sign_in(4188) & VN_data_in(4188);
  VN698_in1 <= VN_sign_in(4189) & VN_data_in(4189);
  VN698_in2 <= VN_sign_in(4190) & VN_data_in(4190);
  VN698_in3 <= VN_sign_in(4191) & VN_data_in(4191);
  VN698_in4 <= VN_sign_in(4192) & VN_data_in(4192);
  VN698_in5 <= VN_sign_in(4193) & VN_data_in(4193);
  VN699_in0 <= VN_sign_in(4194) & VN_data_in(4194);
  VN699_in1 <= VN_sign_in(4195) & VN_data_in(4195);
  VN699_in2 <= VN_sign_in(4196) & VN_data_in(4196);
  VN699_in3 <= VN_sign_in(4197) & VN_data_in(4197);
  VN699_in4 <= VN_sign_in(4198) & VN_data_in(4198);
  VN699_in5 <= VN_sign_in(4199) & VN_data_in(4199);
  VN700_in0 <= VN_sign_in(4200) & VN_data_in(4200);
  VN700_in1 <= VN_sign_in(4201) & VN_data_in(4201);
  VN700_in2 <= VN_sign_in(4202) & VN_data_in(4202);
  VN700_in3 <= VN_sign_in(4203) & VN_data_in(4203);
  VN700_in4 <= VN_sign_in(4204) & VN_data_in(4204);
  VN700_in5 <= VN_sign_in(4205) & VN_data_in(4205);
  VN701_in0 <= VN_sign_in(4206) & VN_data_in(4206);
  VN701_in1 <= VN_sign_in(4207) & VN_data_in(4207);
  VN701_in2 <= VN_sign_in(4208) & VN_data_in(4208);
  VN701_in3 <= VN_sign_in(4209) & VN_data_in(4209);
  VN701_in4 <= VN_sign_in(4210) & VN_data_in(4210);
  VN701_in5 <= VN_sign_in(4211) & VN_data_in(4211);
  VN702_in0 <= VN_sign_in(4212) & VN_data_in(4212);
  VN702_in1 <= VN_sign_in(4213) & VN_data_in(4213);
  VN702_in2 <= VN_sign_in(4214) & VN_data_in(4214);
  VN702_in3 <= VN_sign_in(4215) & VN_data_in(4215);
  VN702_in4 <= VN_sign_in(4216) & VN_data_in(4216);
  VN702_in5 <= VN_sign_in(4217) & VN_data_in(4217);
  VN703_in0 <= VN_sign_in(4218) & VN_data_in(4218);
  VN703_in1 <= VN_sign_in(4219) & VN_data_in(4219);
  VN703_in2 <= VN_sign_in(4220) & VN_data_in(4220);
  VN703_in3 <= VN_sign_in(4221) & VN_data_in(4221);
  VN703_in4 <= VN_sign_in(4222) & VN_data_in(4222);
  VN703_in5 <= VN_sign_in(4223) & VN_data_in(4223);
  VN704_in0 <= VN_sign_in(4224) & VN_data_in(4224);
  VN704_in1 <= VN_sign_in(4225) & VN_data_in(4225);
  VN704_in2 <= VN_sign_in(4226) & VN_data_in(4226);
  VN704_in3 <= VN_sign_in(4227) & VN_data_in(4227);
  VN704_in4 <= VN_sign_in(4228) & VN_data_in(4228);
  VN704_in5 <= VN_sign_in(4229) & VN_data_in(4229);
  VN705_in0 <= VN_sign_in(4230) & VN_data_in(4230);
  VN705_in1 <= VN_sign_in(4231) & VN_data_in(4231);
  VN705_in2 <= VN_sign_in(4232) & VN_data_in(4232);
  VN705_in3 <= VN_sign_in(4233) & VN_data_in(4233);
  VN705_in4 <= VN_sign_in(4234) & VN_data_in(4234);
  VN705_in5 <= VN_sign_in(4235) & VN_data_in(4235);
  VN706_in0 <= VN_sign_in(4236) & VN_data_in(4236);
  VN706_in1 <= VN_sign_in(4237) & VN_data_in(4237);
  VN706_in2 <= VN_sign_in(4238) & VN_data_in(4238);
  VN706_in3 <= VN_sign_in(4239) & VN_data_in(4239);
  VN706_in4 <= VN_sign_in(4240) & VN_data_in(4240);
  VN706_in5 <= VN_sign_in(4241) & VN_data_in(4241);
  VN707_in0 <= VN_sign_in(4242) & VN_data_in(4242);
  VN707_in1 <= VN_sign_in(4243) & VN_data_in(4243);
  VN707_in2 <= VN_sign_in(4244) & VN_data_in(4244);
  VN707_in3 <= VN_sign_in(4245) & VN_data_in(4245);
  VN707_in4 <= VN_sign_in(4246) & VN_data_in(4246);
  VN707_in5 <= VN_sign_in(4247) & VN_data_in(4247);
  VN708_in0 <= VN_sign_in(4248) & VN_data_in(4248);
  VN708_in1 <= VN_sign_in(4249) & VN_data_in(4249);
  VN708_in2 <= VN_sign_in(4250) & VN_data_in(4250);
  VN708_in3 <= VN_sign_in(4251) & VN_data_in(4251);
  VN708_in4 <= VN_sign_in(4252) & VN_data_in(4252);
  VN708_in5 <= VN_sign_in(4253) & VN_data_in(4253);
  VN709_in0 <= VN_sign_in(4254) & VN_data_in(4254);
  VN709_in1 <= VN_sign_in(4255) & VN_data_in(4255);
  VN709_in2 <= VN_sign_in(4256) & VN_data_in(4256);
  VN709_in3 <= VN_sign_in(4257) & VN_data_in(4257);
  VN709_in4 <= VN_sign_in(4258) & VN_data_in(4258);
  VN709_in5 <= VN_sign_in(4259) & VN_data_in(4259);
  VN710_in0 <= VN_sign_in(4260) & VN_data_in(4260);
  VN710_in1 <= VN_sign_in(4261) & VN_data_in(4261);
  VN710_in2 <= VN_sign_in(4262) & VN_data_in(4262);
  VN710_in3 <= VN_sign_in(4263) & VN_data_in(4263);
  VN710_in4 <= VN_sign_in(4264) & VN_data_in(4264);
  VN710_in5 <= VN_sign_in(4265) & VN_data_in(4265);
  VN711_in0 <= VN_sign_in(4266) & VN_data_in(4266);
  VN711_in1 <= VN_sign_in(4267) & VN_data_in(4267);
  VN711_in2 <= VN_sign_in(4268) & VN_data_in(4268);
  VN711_in3 <= VN_sign_in(4269) & VN_data_in(4269);
  VN711_in4 <= VN_sign_in(4270) & VN_data_in(4270);
  VN711_in5 <= VN_sign_in(4271) & VN_data_in(4271);
  VN712_in0 <= VN_sign_in(4272) & VN_data_in(4272);
  VN712_in1 <= VN_sign_in(4273) & VN_data_in(4273);
  VN712_in2 <= VN_sign_in(4274) & VN_data_in(4274);
  VN712_in3 <= VN_sign_in(4275) & VN_data_in(4275);
  VN712_in4 <= VN_sign_in(4276) & VN_data_in(4276);
  VN712_in5 <= VN_sign_in(4277) & VN_data_in(4277);
  VN713_in0 <= VN_sign_in(4278) & VN_data_in(4278);
  VN713_in1 <= VN_sign_in(4279) & VN_data_in(4279);
  VN713_in2 <= VN_sign_in(4280) & VN_data_in(4280);
  VN713_in3 <= VN_sign_in(4281) & VN_data_in(4281);
  VN713_in4 <= VN_sign_in(4282) & VN_data_in(4282);
  VN713_in5 <= VN_sign_in(4283) & VN_data_in(4283);
  VN714_in0 <= VN_sign_in(4284) & VN_data_in(4284);
  VN714_in1 <= VN_sign_in(4285) & VN_data_in(4285);
  VN714_in2 <= VN_sign_in(4286) & VN_data_in(4286);
  VN714_in3 <= VN_sign_in(4287) & VN_data_in(4287);
  VN714_in4 <= VN_sign_in(4288) & VN_data_in(4288);
  VN714_in5 <= VN_sign_in(4289) & VN_data_in(4289);
  VN715_in0 <= VN_sign_in(4290) & VN_data_in(4290);
  VN715_in1 <= VN_sign_in(4291) & VN_data_in(4291);
  VN715_in2 <= VN_sign_in(4292) & VN_data_in(4292);
  VN715_in3 <= VN_sign_in(4293) & VN_data_in(4293);
  VN715_in4 <= VN_sign_in(4294) & VN_data_in(4294);
  VN715_in5 <= VN_sign_in(4295) & VN_data_in(4295);
  VN716_in0 <= VN_sign_in(4296) & VN_data_in(4296);
  VN716_in1 <= VN_sign_in(4297) & VN_data_in(4297);
  VN716_in2 <= VN_sign_in(4298) & VN_data_in(4298);
  VN716_in3 <= VN_sign_in(4299) & VN_data_in(4299);
  VN716_in4 <= VN_sign_in(4300) & VN_data_in(4300);
  VN716_in5 <= VN_sign_in(4301) & VN_data_in(4301);
  VN717_in0 <= VN_sign_in(4302) & VN_data_in(4302);
  VN717_in1 <= VN_sign_in(4303) & VN_data_in(4303);
  VN717_in2 <= VN_sign_in(4304) & VN_data_in(4304);
  VN717_in3 <= VN_sign_in(4305) & VN_data_in(4305);
  VN717_in4 <= VN_sign_in(4306) & VN_data_in(4306);
  VN717_in5 <= VN_sign_in(4307) & VN_data_in(4307);
  VN718_in0 <= VN_sign_in(4308) & VN_data_in(4308);
  VN718_in1 <= VN_sign_in(4309) & VN_data_in(4309);
  VN718_in2 <= VN_sign_in(4310) & VN_data_in(4310);
  VN718_in3 <= VN_sign_in(4311) & VN_data_in(4311);
  VN718_in4 <= VN_sign_in(4312) & VN_data_in(4312);
  VN718_in5 <= VN_sign_in(4313) & VN_data_in(4313);
  VN719_in0 <= VN_sign_in(4314) & VN_data_in(4314);
  VN719_in1 <= VN_sign_in(4315) & VN_data_in(4315);
  VN719_in2 <= VN_sign_in(4316) & VN_data_in(4316);
  VN719_in3 <= VN_sign_in(4317) & VN_data_in(4317);
  VN719_in4 <= VN_sign_in(4318) & VN_data_in(4318);
  VN719_in5 <= VN_sign_in(4319) & VN_data_in(4319);
  VN720_in0 <= VN_sign_in(4320) & VN_data_in(4320);
  VN720_in1 <= VN_sign_in(4321) & VN_data_in(4321);
  VN720_in2 <= VN_sign_in(4322) & VN_data_in(4322);
  VN720_in3 <= VN_sign_in(4323) & VN_data_in(4323);
  VN720_in4 <= VN_sign_in(4324) & VN_data_in(4324);
  VN720_in5 <= VN_sign_in(4325) & VN_data_in(4325);
  VN721_in0 <= VN_sign_in(4326) & VN_data_in(4326);
  VN721_in1 <= VN_sign_in(4327) & VN_data_in(4327);
  VN721_in2 <= VN_sign_in(4328) & VN_data_in(4328);
  VN721_in3 <= VN_sign_in(4329) & VN_data_in(4329);
  VN721_in4 <= VN_sign_in(4330) & VN_data_in(4330);
  VN721_in5 <= VN_sign_in(4331) & VN_data_in(4331);
  VN722_in0 <= VN_sign_in(4332) & VN_data_in(4332);
  VN722_in1 <= VN_sign_in(4333) & VN_data_in(4333);
  VN722_in2 <= VN_sign_in(4334) & VN_data_in(4334);
  VN722_in3 <= VN_sign_in(4335) & VN_data_in(4335);
  VN722_in4 <= VN_sign_in(4336) & VN_data_in(4336);
  VN722_in5 <= VN_sign_in(4337) & VN_data_in(4337);
  VN723_in0 <= VN_sign_in(4338) & VN_data_in(4338);
  VN723_in1 <= VN_sign_in(4339) & VN_data_in(4339);
  VN723_in2 <= VN_sign_in(4340) & VN_data_in(4340);
  VN723_in3 <= VN_sign_in(4341) & VN_data_in(4341);
  VN723_in4 <= VN_sign_in(4342) & VN_data_in(4342);
  VN723_in5 <= VN_sign_in(4343) & VN_data_in(4343);
  VN724_in0 <= VN_sign_in(4344) & VN_data_in(4344);
  VN724_in1 <= VN_sign_in(4345) & VN_data_in(4345);
  VN724_in2 <= VN_sign_in(4346) & VN_data_in(4346);
  VN724_in3 <= VN_sign_in(4347) & VN_data_in(4347);
  VN724_in4 <= VN_sign_in(4348) & VN_data_in(4348);
  VN724_in5 <= VN_sign_in(4349) & VN_data_in(4349);
  VN725_in0 <= VN_sign_in(4350) & VN_data_in(4350);
  VN725_in1 <= VN_sign_in(4351) & VN_data_in(4351);
  VN725_in2 <= VN_sign_in(4352) & VN_data_in(4352);
  VN725_in3 <= VN_sign_in(4353) & VN_data_in(4353);
  VN725_in4 <= VN_sign_in(4354) & VN_data_in(4354);
  VN725_in5 <= VN_sign_in(4355) & VN_data_in(4355);
  VN726_in0 <= VN_sign_in(4356) & VN_data_in(4356);
  VN726_in1 <= VN_sign_in(4357) & VN_data_in(4357);
  VN726_in2 <= VN_sign_in(4358) & VN_data_in(4358);
  VN726_in3 <= VN_sign_in(4359) & VN_data_in(4359);
  VN726_in4 <= VN_sign_in(4360) & VN_data_in(4360);
  VN726_in5 <= VN_sign_in(4361) & VN_data_in(4361);
  VN727_in0 <= VN_sign_in(4362) & VN_data_in(4362);
  VN727_in1 <= VN_sign_in(4363) & VN_data_in(4363);
  VN727_in2 <= VN_sign_in(4364) & VN_data_in(4364);
  VN727_in3 <= VN_sign_in(4365) & VN_data_in(4365);
  VN727_in4 <= VN_sign_in(4366) & VN_data_in(4366);
  VN727_in5 <= VN_sign_in(4367) & VN_data_in(4367);
  VN728_in0 <= VN_sign_in(4368) & VN_data_in(4368);
  VN728_in1 <= VN_sign_in(4369) & VN_data_in(4369);
  VN728_in2 <= VN_sign_in(4370) & VN_data_in(4370);
  VN728_in3 <= VN_sign_in(4371) & VN_data_in(4371);
  VN728_in4 <= VN_sign_in(4372) & VN_data_in(4372);
  VN728_in5 <= VN_sign_in(4373) & VN_data_in(4373);
  VN729_in0 <= VN_sign_in(4374) & VN_data_in(4374);
  VN729_in1 <= VN_sign_in(4375) & VN_data_in(4375);
  VN729_in2 <= VN_sign_in(4376) & VN_data_in(4376);
  VN729_in3 <= VN_sign_in(4377) & VN_data_in(4377);
  VN729_in4 <= VN_sign_in(4378) & VN_data_in(4378);
  VN729_in5 <= VN_sign_in(4379) & VN_data_in(4379);
  VN730_in0 <= VN_sign_in(4380) & VN_data_in(4380);
  VN730_in1 <= VN_sign_in(4381) & VN_data_in(4381);
  VN730_in2 <= VN_sign_in(4382) & VN_data_in(4382);
  VN730_in3 <= VN_sign_in(4383) & VN_data_in(4383);
  VN730_in4 <= VN_sign_in(4384) & VN_data_in(4384);
  VN730_in5 <= VN_sign_in(4385) & VN_data_in(4385);
  VN731_in0 <= VN_sign_in(4386) & VN_data_in(4386);
  VN731_in1 <= VN_sign_in(4387) & VN_data_in(4387);
  VN731_in2 <= VN_sign_in(4388) & VN_data_in(4388);
  VN731_in3 <= VN_sign_in(4389) & VN_data_in(4389);
  VN731_in4 <= VN_sign_in(4390) & VN_data_in(4390);
  VN731_in5 <= VN_sign_in(4391) & VN_data_in(4391);
  VN732_in0 <= VN_sign_in(4392) & VN_data_in(4392);
  VN732_in1 <= VN_sign_in(4393) & VN_data_in(4393);
  VN732_in2 <= VN_sign_in(4394) & VN_data_in(4394);
  VN732_in3 <= VN_sign_in(4395) & VN_data_in(4395);
  VN732_in4 <= VN_sign_in(4396) & VN_data_in(4396);
  VN732_in5 <= VN_sign_in(4397) & VN_data_in(4397);
  VN733_in0 <= VN_sign_in(4398) & VN_data_in(4398);
  VN733_in1 <= VN_sign_in(4399) & VN_data_in(4399);
  VN733_in2 <= VN_sign_in(4400) & VN_data_in(4400);
  VN733_in3 <= VN_sign_in(4401) & VN_data_in(4401);
  VN733_in4 <= VN_sign_in(4402) & VN_data_in(4402);
  VN733_in5 <= VN_sign_in(4403) & VN_data_in(4403);
  VN734_in0 <= VN_sign_in(4404) & VN_data_in(4404);
  VN734_in1 <= VN_sign_in(4405) & VN_data_in(4405);
  VN734_in2 <= VN_sign_in(4406) & VN_data_in(4406);
  VN734_in3 <= VN_sign_in(4407) & VN_data_in(4407);
  VN734_in4 <= VN_sign_in(4408) & VN_data_in(4408);
  VN734_in5 <= VN_sign_in(4409) & VN_data_in(4409);
  VN735_in0 <= VN_sign_in(4410) & VN_data_in(4410);
  VN735_in1 <= VN_sign_in(4411) & VN_data_in(4411);
  VN735_in2 <= VN_sign_in(4412) & VN_data_in(4412);
  VN735_in3 <= VN_sign_in(4413) & VN_data_in(4413);
  VN735_in4 <= VN_sign_in(4414) & VN_data_in(4414);
  VN735_in5 <= VN_sign_in(4415) & VN_data_in(4415);
  VN736_in0 <= VN_sign_in(4416) & VN_data_in(4416);
  VN736_in1 <= VN_sign_in(4417) & VN_data_in(4417);
  VN736_in2 <= VN_sign_in(4418) & VN_data_in(4418);
  VN736_in3 <= VN_sign_in(4419) & VN_data_in(4419);
  VN736_in4 <= VN_sign_in(4420) & VN_data_in(4420);
  VN736_in5 <= VN_sign_in(4421) & VN_data_in(4421);
  VN737_in0 <= VN_sign_in(4422) & VN_data_in(4422);
  VN737_in1 <= VN_sign_in(4423) & VN_data_in(4423);
  VN737_in2 <= VN_sign_in(4424) & VN_data_in(4424);
  VN737_in3 <= VN_sign_in(4425) & VN_data_in(4425);
  VN737_in4 <= VN_sign_in(4426) & VN_data_in(4426);
  VN737_in5 <= VN_sign_in(4427) & VN_data_in(4427);
  VN738_in0 <= VN_sign_in(4428) & VN_data_in(4428);
  VN738_in1 <= VN_sign_in(4429) & VN_data_in(4429);
  VN738_in2 <= VN_sign_in(4430) & VN_data_in(4430);
  VN738_in3 <= VN_sign_in(4431) & VN_data_in(4431);
  VN738_in4 <= VN_sign_in(4432) & VN_data_in(4432);
  VN738_in5 <= VN_sign_in(4433) & VN_data_in(4433);
  VN739_in0 <= VN_sign_in(4434) & VN_data_in(4434);
  VN739_in1 <= VN_sign_in(4435) & VN_data_in(4435);
  VN739_in2 <= VN_sign_in(4436) & VN_data_in(4436);
  VN739_in3 <= VN_sign_in(4437) & VN_data_in(4437);
  VN739_in4 <= VN_sign_in(4438) & VN_data_in(4438);
  VN739_in5 <= VN_sign_in(4439) & VN_data_in(4439);
  VN740_in0 <= VN_sign_in(4440) & VN_data_in(4440);
  VN740_in1 <= VN_sign_in(4441) & VN_data_in(4441);
  VN740_in2 <= VN_sign_in(4442) & VN_data_in(4442);
  VN740_in3 <= VN_sign_in(4443) & VN_data_in(4443);
  VN740_in4 <= VN_sign_in(4444) & VN_data_in(4444);
  VN740_in5 <= VN_sign_in(4445) & VN_data_in(4445);
  VN741_in0 <= VN_sign_in(4446) & VN_data_in(4446);
  VN741_in1 <= VN_sign_in(4447) & VN_data_in(4447);
  VN741_in2 <= VN_sign_in(4448) & VN_data_in(4448);
  VN741_in3 <= VN_sign_in(4449) & VN_data_in(4449);
  VN741_in4 <= VN_sign_in(4450) & VN_data_in(4450);
  VN741_in5 <= VN_sign_in(4451) & VN_data_in(4451);
  VN742_in0 <= VN_sign_in(4452) & VN_data_in(4452);
  VN742_in1 <= VN_sign_in(4453) & VN_data_in(4453);
  VN742_in2 <= VN_sign_in(4454) & VN_data_in(4454);
  VN742_in3 <= VN_sign_in(4455) & VN_data_in(4455);
  VN742_in4 <= VN_sign_in(4456) & VN_data_in(4456);
  VN742_in5 <= VN_sign_in(4457) & VN_data_in(4457);
  VN743_in0 <= VN_sign_in(4458) & VN_data_in(4458);
  VN743_in1 <= VN_sign_in(4459) & VN_data_in(4459);
  VN743_in2 <= VN_sign_in(4460) & VN_data_in(4460);
  VN743_in3 <= VN_sign_in(4461) & VN_data_in(4461);
  VN743_in4 <= VN_sign_in(4462) & VN_data_in(4462);
  VN743_in5 <= VN_sign_in(4463) & VN_data_in(4463);
  VN744_in0 <= VN_sign_in(4464) & VN_data_in(4464);
  VN744_in1 <= VN_sign_in(4465) & VN_data_in(4465);
  VN744_in2 <= VN_sign_in(4466) & VN_data_in(4466);
  VN744_in3 <= VN_sign_in(4467) & VN_data_in(4467);
  VN744_in4 <= VN_sign_in(4468) & VN_data_in(4468);
  VN744_in5 <= VN_sign_in(4469) & VN_data_in(4469);
  VN745_in0 <= VN_sign_in(4470) & VN_data_in(4470);
  VN745_in1 <= VN_sign_in(4471) & VN_data_in(4471);
  VN745_in2 <= VN_sign_in(4472) & VN_data_in(4472);
  VN745_in3 <= VN_sign_in(4473) & VN_data_in(4473);
  VN745_in4 <= VN_sign_in(4474) & VN_data_in(4474);
  VN745_in5 <= VN_sign_in(4475) & VN_data_in(4475);
  VN746_in0 <= VN_sign_in(4476) & VN_data_in(4476);
  VN746_in1 <= VN_sign_in(4477) & VN_data_in(4477);
  VN746_in2 <= VN_sign_in(4478) & VN_data_in(4478);
  VN746_in3 <= VN_sign_in(4479) & VN_data_in(4479);
  VN746_in4 <= VN_sign_in(4480) & VN_data_in(4480);
  VN746_in5 <= VN_sign_in(4481) & VN_data_in(4481);
  VN747_in0 <= VN_sign_in(4482) & VN_data_in(4482);
  VN747_in1 <= VN_sign_in(4483) & VN_data_in(4483);
  VN747_in2 <= VN_sign_in(4484) & VN_data_in(4484);
  VN747_in3 <= VN_sign_in(4485) & VN_data_in(4485);
  VN747_in4 <= VN_sign_in(4486) & VN_data_in(4486);
  VN747_in5 <= VN_sign_in(4487) & VN_data_in(4487);
  VN748_in0 <= VN_sign_in(4488) & VN_data_in(4488);
  VN748_in1 <= VN_sign_in(4489) & VN_data_in(4489);
  VN748_in2 <= VN_sign_in(4490) & VN_data_in(4490);
  VN748_in3 <= VN_sign_in(4491) & VN_data_in(4491);
  VN748_in4 <= VN_sign_in(4492) & VN_data_in(4492);
  VN748_in5 <= VN_sign_in(4493) & VN_data_in(4493);
  VN749_in0 <= VN_sign_in(4494) & VN_data_in(4494);
  VN749_in1 <= VN_sign_in(4495) & VN_data_in(4495);
  VN749_in2 <= VN_sign_in(4496) & VN_data_in(4496);
  VN749_in3 <= VN_sign_in(4497) & VN_data_in(4497);
  VN749_in4 <= VN_sign_in(4498) & VN_data_in(4498);
  VN749_in5 <= VN_sign_in(4499) & VN_data_in(4499);
  VN750_in0 <= VN_sign_in(4500) & VN_data_in(4500);
  VN750_in1 <= VN_sign_in(4501) & VN_data_in(4501);
  VN750_in2 <= VN_sign_in(4502) & VN_data_in(4502);
  VN750_in3 <= VN_sign_in(4503) & VN_data_in(4503);
  VN750_in4 <= VN_sign_in(4504) & VN_data_in(4504);
  VN750_in5 <= VN_sign_in(4505) & VN_data_in(4505);
  VN751_in0 <= VN_sign_in(4506) & VN_data_in(4506);
  VN751_in1 <= VN_sign_in(4507) & VN_data_in(4507);
  VN751_in2 <= VN_sign_in(4508) & VN_data_in(4508);
  VN751_in3 <= VN_sign_in(4509) & VN_data_in(4509);
  VN751_in4 <= VN_sign_in(4510) & VN_data_in(4510);
  VN751_in5 <= VN_sign_in(4511) & VN_data_in(4511);
  VN752_in0 <= VN_sign_in(4512) & VN_data_in(4512);
  VN752_in1 <= VN_sign_in(4513) & VN_data_in(4513);
  VN752_in2 <= VN_sign_in(4514) & VN_data_in(4514);
  VN752_in3 <= VN_sign_in(4515) & VN_data_in(4515);
  VN752_in4 <= VN_sign_in(4516) & VN_data_in(4516);
  VN752_in5 <= VN_sign_in(4517) & VN_data_in(4517);
  VN753_in0 <= VN_sign_in(4518) & VN_data_in(4518);
  VN753_in1 <= VN_sign_in(4519) & VN_data_in(4519);
  VN753_in2 <= VN_sign_in(4520) & VN_data_in(4520);
  VN753_in3 <= VN_sign_in(4521) & VN_data_in(4521);
  VN753_in4 <= VN_sign_in(4522) & VN_data_in(4522);
  VN753_in5 <= VN_sign_in(4523) & VN_data_in(4523);
  VN754_in0 <= VN_sign_in(4524) & VN_data_in(4524);
  VN754_in1 <= VN_sign_in(4525) & VN_data_in(4525);
  VN754_in2 <= VN_sign_in(4526) & VN_data_in(4526);
  VN754_in3 <= VN_sign_in(4527) & VN_data_in(4527);
  VN754_in4 <= VN_sign_in(4528) & VN_data_in(4528);
  VN754_in5 <= VN_sign_in(4529) & VN_data_in(4529);
  VN755_in0 <= VN_sign_in(4530) & VN_data_in(4530);
  VN755_in1 <= VN_sign_in(4531) & VN_data_in(4531);
  VN755_in2 <= VN_sign_in(4532) & VN_data_in(4532);
  VN755_in3 <= VN_sign_in(4533) & VN_data_in(4533);
  VN755_in4 <= VN_sign_in(4534) & VN_data_in(4534);
  VN755_in5 <= VN_sign_in(4535) & VN_data_in(4535);
  VN756_in0 <= VN_sign_in(4536) & VN_data_in(4536);
  VN756_in1 <= VN_sign_in(4537) & VN_data_in(4537);
  VN756_in2 <= VN_sign_in(4538) & VN_data_in(4538);
  VN756_in3 <= VN_sign_in(4539) & VN_data_in(4539);
  VN756_in4 <= VN_sign_in(4540) & VN_data_in(4540);
  VN756_in5 <= VN_sign_in(4541) & VN_data_in(4541);
  VN757_in0 <= VN_sign_in(4542) & VN_data_in(4542);
  VN757_in1 <= VN_sign_in(4543) & VN_data_in(4543);
  VN757_in2 <= VN_sign_in(4544) & VN_data_in(4544);
  VN757_in3 <= VN_sign_in(4545) & VN_data_in(4545);
  VN757_in4 <= VN_sign_in(4546) & VN_data_in(4546);
  VN757_in5 <= VN_sign_in(4547) & VN_data_in(4547);
  VN758_in0 <= VN_sign_in(4548) & VN_data_in(4548);
  VN758_in1 <= VN_sign_in(4549) & VN_data_in(4549);
  VN758_in2 <= VN_sign_in(4550) & VN_data_in(4550);
  VN758_in3 <= VN_sign_in(4551) & VN_data_in(4551);
  VN758_in4 <= VN_sign_in(4552) & VN_data_in(4552);
  VN758_in5 <= VN_sign_in(4553) & VN_data_in(4553);
  VN759_in0 <= VN_sign_in(4554) & VN_data_in(4554);
  VN759_in1 <= VN_sign_in(4555) & VN_data_in(4555);
  VN759_in2 <= VN_sign_in(4556) & VN_data_in(4556);
  VN759_in3 <= VN_sign_in(4557) & VN_data_in(4557);
  VN759_in4 <= VN_sign_in(4558) & VN_data_in(4558);
  VN759_in5 <= VN_sign_in(4559) & VN_data_in(4559);
  VN760_in0 <= VN_sign_in(4560) & VN_data_in(4560);
  VN760_in1 <= VN_sign_in(4561) & VN_data_in(4561);
  VN760_in2 <= VN_sign_in(4562) & VN_data_in(4562);
  VN760_in3 <= VN_sign_in(4563) & VN_data_in(4563);
  VN760_in4 <= VN_sign_in(4564) & VN_data_in(4564);
  VN760_in5 <= VN_sign_in(4565) & VN_data_in(4565);
  VN761_in0 <= VN_sign_in(4566) & VN_data_in(4566);
  VN761_in1 <= VN_sign_in(4567) & VN_data_in(4567);
  VN761_in2 <= VN_sign_in(4568) & VN_data_in(4568);
  VN761_in3 <= VN_sign_in(4569) & VN_data_in(4569);
  VN761_in4 <= VN_sign_in(4570) & VN_data_in(4570);
  VN761_in5 <= VN_sign_in(4571) & VN_data_in(4571);
  VN762_in0 <= VN_sign_in(4572) & VN_data_in(4572);
  VN762_in1 <= VN_sign_in(4573) & VN_data_in(4573);
  VN762_in2 <= VN_sign_in(4574) & VN_data_in(4574);
  VN762_in3 <= VN_sign_in(4575) & VN_data_in(4575);
  VN762_in4 <= VN_sign_in(4576) & VN_data_in(4576);
  VN762_in5 <= VN_sign_in(4577) & VN_data_in(4577);
  VN763_in0 <= VN_sign_in(4578) & VN_data_in(4578);
  VN763_in1 <= VN_sign_in(4579) & VN_data_in(4579);
  VN763_in2 <= VN_sign_in(4580) & VN_data_in(4580);
  VN763_in3 <= VN_sign_in(4581) & VN_data_in(4581);
  VN763_in4 <= VN_sign_in(4582) & VN_data_in(4582);
  VN763_in5 <= VN_sign_in(4583) & VN_data_in(4583);
  VN764_in0 <= VN_sign_in(4584) & VN_data_in(4584);
  VN764_in1 <= VN_sign_in(4585) & VN_data_in(4585);
  VN764_in2 <= VN_sign_in(4586) & VN_data_in(4586);
  VN764_in3 <= VN_sign_in(4587) & VN_data_in(4587);
  VN764_in4 <= VN_sign_in(4588) & VN_data_in(4588);
  VN764_in5 <= VN_sign_in(4589) & VN_data_in(4589);
  VN765_in0 <= VN_sign_in(4590) & VN_data_in(4590);
  VN765_in1 <= VN_sign_in(4591) & VN_data_in(4591);
  VN765_in2 <= VN_sign_in(4592) & VN_data_in(4592);
  VN765_in3 <= VN_sign_in(4593) & VN_data_in(4593);
  VN765_in4 <= VN_sign_in(4594) & VN_data_in(4594);
  VN765_in5 <= VN_sign_in(4595) & VN_data_in(4595);
  VN766_in0 <= VN_sign_in(4596) & VN_data_in(4596);
  VN766_in1 <= VN_sign_in(4597) & VN_data_in(4597);
  VN766_in2 <= VN_sign_in(4598) & VN_data_in(4598);
  VN766_in3 <= VN_sign_in(4599) & VN_data_in(4599);
  VN766_in4 <= VN_sign_in(4600) & VN_data_in(4600);
  VN766_in5 <= VN_sign_in(4601) & VN_data_in(4601);
  VN767_in0 <= VN_sign_in(4602) & VN_data_in(4602);
  VN767_in1 <= VN_sign_in(4603) & VN_data_in(4603);
  VN767_in2 <= VN_sign_in(4604) & VN_data_in(4604);
  VN767_in3 <= VN_sign_in(4605) & VN_data_in(4605);
  VN767_in4 <= VN_sign_in(4606) & VN_data_in(4606);
  VN767_in5 <= VN_sign_in(4607) & VN_data_in(4607);
  VN768_in0 <= VN_sign_in(4608) & VN_data_in(4608);
  VN768_in1 <= VN_sign_in(4609) & VN_data_in(4609);
  VN768_in2 <= VN_sign_in(4610) & VN_data_in(4610);
  VN768_in3 <= VN_sign_in(4611) & VN_data_in(4611);
  VN768_in4 <= VN_sign_in(4612) & VN_data_in(4612);
  VN768_in5 <= VN_sign_in(4613) & VN_data_in(4613);
  VN769_in0 <= VN_sign_in(4614) & VN_data_in(4614);
  VN769_in1 <= VN_sign_in(4615) & VN_data_in(4615);
  VN769_in2 <= VN_sign_in(4616) & VN_data_in(4616);
  VN769_in3 <= VN_sign_in(4617) & VN_data_in(4617);
  VN769_in4 <= VN_sign_in(4618) & VN_data_in(4618);
  VN769_in5 <= VN_sign_in(4619) & VN_data_in(4619);
  VN770_in0 <= VN_sign_in(4620) & VN_data_in(4620);
  VN770_in1 <= VN_sign_in(4621) & VN_data_in(4621);
  VN770_in2 <= VN_sign_in(4622) & VN_data_in(4622);
  VN770_in3 <= VN_sign_in(4623) & VN_data_in(4623);
  VN770_in4 <= VN_sign_in(4624) & VN_data_in(4624);
  VN770_in5 <= VN_sign_in(4625) & VN_data_in(4625);
  VN771_in0 <= VN_sign_in(4626) & VN_data_in(4626);
  VN771_in1 <= VN_sign_in(4627) & VN_data_in(4627);
  VN771_in2 <= VN_sign_in(4628) & VN_data_in(4628);
  VN771_in3 <= VN_sign_in(4629) & VN_data_in(4629);
  VN771_in4 <= VN_sign_in(4630) & VN_data_in(4630);
  VN771_in5 <= VN_sign_in(4631) & VN_data_in(4631);
  VN772_in0 <= VN_sign_in(4632) & VN_data_in(4632);
  VN772_in1 <= VN_sign_in(4633) & VN_data_in(4633);
  VN772_in2 <= VN_sign_in(4634) & VN_data_in(4634);
  VN772_in3 <= VN_sign_in(4635) & VN_data_in(4635);
  VN772_in4 <= VN_sign_in(4636) & VN_data_in(4636);
  VN772_in5 <= VN_sign_in(4637) & VN_data_in(4637);
  VN773_in0 <= VN_sign_in(4638) & VN_data_in(4638);
  VN773_in1 <= VN_sign_in(4639) & VN_data_in(4639);
  VN773_in2 <= VN_sign_in(4640) & VN_data_in(4640);
  VN773_in3 <= VN_sign_in(4641) & VN_data_in(4641);
  VN773_in4 <= VN_sign_in(4642) & VN_data_in(4642);
  VN773_in5 <= VN_sign_in(4643) & VN_data_in(4643);
  VN774_in0 <= VN_sign_in(4644) & VN_data_in(4644);
  VN774_in1 <= VN_sign_in(4645) & VN_data_in(4645);
  VN774_in2 <= VN_sign_in(4646) & VN_data_in(4646);
  VN774_in3 <= VN_sign_in(4647) & VN_data_in(4647);
  VN774_in4 <= VN_sign_in(4648) & VN_data_in(4648);
  VN774_in5 <= VN_sign_in(4649) & VN_data_in(4649);
  VN775_in0 <= VN_sign_in(4650) & VN_data_in(4650);
  VN775_in1 <= VN_sign_in(4651) & VN_data_in(4651);
  VN775_in2 <= VN_sign_in(4652) & VN_data_in(4652);
  VN775_in3 <= VN_sign_in(4653) & VN_data_in(4653);
  VN775_in4 <= VN_sign_in(4654) & VN_data_in(4654);
  VN775_in5 <= VN_sign_in(4655) & VN_data_in(4655);
  VN776_in0 <= VN_sign_in(4656) & VN_data_in(4656);
  VN776_in1 <= VN_sign_in(4657) & VN_data_in(4657);
  VN776_in2 <= VN_sign_in(4658) & VN_data_in(4658);
  VN776_in3 <= VN_sign_in(4659) & VN_data_in(4659);
  VN776_in4 <= VN_sign_in(4660) & VN_data_in(4660);
  VN776_in5 <= VN_sign_in(4661) & VN_data_in(4661);
  VN777_in0 <= VN_sign_in(4662) & VN_data_in(4662);
  VN777_in1 <= VN_sign_in(4663) & VN_data_in(4663);
  VN777_in2 <= VN_sign_in(4664) & VN_data_in(4664);
  VN777_in3 <= VN_sign_in(4665) & VN_data_in(4665);
  VN777_in4 <= VN_sign_in(4666) & VN_data_in(4666);
  VN777_in5 <= VN_sign_in(4667) & VN_data_in(4667);
  VN778_in0 <= VN_sign_in(4668) & VN_data_in(4668);
  VN778_in1 <= VN_sign_in(4669) & VN_data_in(4669);
  VN778_in2 <= VN_sign_in(4670) & VN_data_in(4670);
  VN778_in3 <= VN_sign_in(4671) & VN_data_in(4671);
  VN778_in4 <= VN_sign_in(4672) & VN_data_in(4672);
  VN778_in5 <= VN_sign_in(4673) & VN_data_in(4673);
  VN779_in0 <= VN_sign_in(4674) & VN_data_in(4674);
  VN779_in1 <= VN_sign_in(4675) & VN_data_in(4675);
  VN779_in2 <= VN_sign_in(4676) & VN_data_in(4676);
  VN779_in3 <= VN_sign_in(4677) & VN_data_in(4677);
  VN779_in4 <= VN_sign_in(4678) & VN_data_in(4678);
  VN779_in5 <= VN_sign_in(4679) & VN_data_in(4679);
  VN780_in0 <= VN_sign_in(4680) & VN_data_in(4680);
  VN780_in1 <= VN_sign_in(4681) & VN_data_in(4681);
  VN780_in2 <= VN_sign_in(4682) & VN_data_in(4682);
  VN780_in3 <= VN_sign_in(4683) & VN_data_in(4683);
  VN780_in4 <= VN_sign_in(4684) & VN_data_in(4684);
  VN780_in5 <= VN_sign_in(4685) & VN_data_in(4685);
  VN781_in0 <= VN_sign_in(4686) & VN_data_in(4686);
  VN781_in1 <= VN_sign_in(4687) & VN_data_in(4687);
  VN781_in2 <= VN_sign_in(4688) & VN_data_in(4688);
  VN781_in3 <= VN_sign_in(4689) & VN_data_in(4689);
  VN781_in4 <= VN_sign_in(4690) & VN_data_in(4690);
  VN781_in5 <= VN_sign_in(4691) & VN_data_in(4691);
  VN782_in0 <= VN_sign_in(4692) & VN_data_in(4692);
  VN782_in1 <= VN_sign_in(4693) & VN_data_in(4693);
  VN782_in2 <= VN_sign_in(4694) & VN_data_in(4694);
  VN782_in3 <= VN_sign_in(4695) & VN_data_in(4695);
  VN782_in4 <= VN_sign_in(4696) & VN_data_in(4696);
  VN782_in5 <= VN_sign_in(4697) & VN_data_in(4697);
  VN783_in0 <= VN_sign_in(4698) & VN_data_in(4698);
  VN783_in1 <= VN_sign_in(4699) & VN_data_in(4699);
  VN783_in2 <= VN_sign_in(4700) & VN_data_in(4700);
  VN783_in3 <= VN_sign_in(4701) & VN_data_in(4701);
  VN783_in4 <= VN_sign_in(4702) & VN_data_in(4702);
  VN783_in5 <= VN_sign_in(4703) & VN_data_in(4703);
  VN784_in0 <= VN_sign_in(4704) & VN_data_in(4704);
  VN784_in1 <= VN_sign_in(4705) & VN_data_in(4705);
  VN784_in2 <= VN_sign_in(4706) & VN_data_in(4706);
  VN784_in3 <= VN_sign_in(4707) & VN_data_in(4707);
  VN784_in4 <= VN_sign_in(4708) & VN_data_in(4708);
  VN784_in5 <= VN_sign_in(4709) & VN_data_in(4709);
  VN785_in0 <= VN_sign_in(4710) & VN_data_in(4710);
  VN785_in1 <= VN_sign_in(4711) & VN_data_in(4711);
  VN785_in2 <= VN_sign_in(4712) & VN_data_in(4712);
  VN785_in3 <= VN_sign_in(4713) & VN_data_in(4713);
  VN785_in4 <= VN_sign_in(4714) & VN_data_in(4714);
  VN785_in5 <= VN_sign_in(4715) & VN_data_in(4715);
  VN786_in0 <= VN_sign_in(4716) & VN_data_in(4716);
  VN786_in1 <= VN_sign_in(4717) & VN_data_in(4717);
  VN786_in2 <= VN_sign_in(4718) & VN_data_in(4718);
  VN786_in3 <= VN_sign_in(4719) & VN_data_in(4719);
  VN786_in4 <= VN_sign_in(4720) & VN_data_in(4720);
  VN786_in5 <= VN_sign_in(4721) & VN_data_in(4721);
  VN787_in0 <= VN_sign_in(4722) & VN_data_in(4722);
  VN787_in1 <= VN_sign_in(4723) & VN_data_in(4723);
  VN787_in2 <= VN_sign_in(4724) & VN_data_in(4724);
  VN787_in3 <= VN_sign_in(4725) & VN_data_in(4725);
  VN787_in4 <= VN_sign_in(4726) & VN_data_in(4726);
  VN787_in5 <= VN_sign_in(4727) & VN_data_in(4727);
  VN788_in0 <= VN_sign_in(4728) & VN_data_in(4728);
  VN788_in1 <= VN_sign_in(4729) & VN_data_in(4729);
  VN788_in2 <= VN_sign_in(4730) & VN_data_in(4730);
  VN788_in3 <= VN_sign_in(4731) & VN_data_in(4731);
  VN788_in4 <= VN_sign_in(4732) & VN_data_in(4732);
  VN788_in5 <= VN_sign_in(4733) & VN_data_in(4733);
  VN789_in0 <= VN_sign_in(4734) & VN_data_in(4734);
  VN789_in1 <= VN_sign_in(4735) & VN_data_in(4735);
  VN789_in2 <= VN_sign_in(4736) & VN_data_in(4736);
  VN789_in3 <= VN_sign_in(4737) & VN_data_in(4737);
  VN789_in4 <= VN_sign_in(4738) & VN_data_in(4738);
  VN789_in5 <= VN_sign_in(4739) & VN_data_in(4739);
  VN790_in0 <= VN_sign_in(4740) & VN_data_in(4740);
  VN790_in1 <= VN_sign_in(4741) & VN_data_in(4741);
  VN790_in2 <= VN_sign_in(4742) & VN_data_in(4742);
  VN790_in3 <= VN_sign_in(4743) & VN_data_in(4743);
  VN790_in4 <= VN_sign_in(4744) & VN_data_in(4744);
  VN790_in5 <= VN_sign_in(4745) & VN_data_in(4745);
  VN791_in0 <= VN_sign_in(4746) & VN_data_in(4746);
  VN791_in1 <= VN_sign_in(4747) & VN_data_in(4747);
  VN791_in2 <= VN_sign_in(4748) & VN_data_in(4748);
  VN791_in3 <= VN_sign_in(4749) & VN_data_in(4749);
  VN791_in4 <= VN_sign_in(4750) & VN_data_in(4750);
  VN791_in5 <= VN_sign_in(4751) & VN_data_in(4751);
  VN792_in0 <= VN_sign_in(4752) & VN_data_in(4752);
  VN792_in1 <= VN_sign_in(4753) & VN_data_in(4753);
  VN792_in2 <= VN_sign_in(4754) & VN_data_in(4754);
  VN792_in3 <= VN_sign_in(4755) & VN_data_in(4755);
  VN792_in4 <= VN_sign_in(4756) & VN_data_in(4756);
  VN792_in5 <= VN_sign_in(4757) & VN_data_in(4757);
  VN793_in0 <= VN_sign_in(4758) & VN_data_in(4758);
  VN793_in1 <= VN_sign_in(4759) & VN_data_in(4759);
  VN793_in2 <= VN_sign_in(4760) & VN_data_in(4760);
  VN793_in3 <= VN_sign_in(4761) & VN_data_in(4761);
  VN793_in4 <= VN_sign_in(4762) & VN_data_in(4762);
  VN793_in5 <= VN_sign_in(4763) & VN_data_in(4763);
  VN794_in0 <= VN_sign_in(4764) & VN_data_in(4764);
  VN794_in1 <= VN_sign_in(4765) & VN_data_in(4765);
  VN794_in2 <= VN_sign_in(4766) & VN_data_in(4766);
  VN794_in3 <= VN_sign_in(4767) & VN_data_in(4767);
  VN794_in4 <= VN_sign_in(4768) & VN_data_in(4768);
  VN794_in5 <= VN_sign_in(4769) & VN_data_in(4769);
  VN795_in0 <= VN_sign_in(4770) & VN_data_in(4770);
  VN795_in1 <= VN_sign_in(4771) & VN_data_in(4771);
  VN795_in2 <= VN_sign_in(4772) & VN_data_in(4772);
  VN795_in3 <= VN_sign_in(4773) & VN_data_in(4773);
  VN795_in4 <= VN_sign_in(4774) & VN_data_in(4774);
  VN795_in5 <= VN_sign_in(4775) & VN_data_in(4775);
  VN796_in0 <= VN_sign_in(4776) & VN_data_in(4776);
  VN796_in1 <= VN_sign_in(4777) & VN_data_in(4777);
  VN796_in2 <= VN_sign_in(4778) & VN_data_in(4778);
  VN796_in3 <= VN_sign_in(4779) & VN_data_in(4779);
  VN796_in4 <= VN_sign_in(4780) & VN_data_in(4780);
  VN796_in5 <= VN_sign_in(4781) & VN_data_in(4781);
  VN797_in0 <= VN_sign_in(4782) & VN_data_in(4782);
  VN797_in1 <= VN_sign_in(4783) & VN_data_in(4783);
  VN797_in2 <= VN_sign_in(4784) & VN_data_in(4784);
  VN797_in3 <= VN_sign_in(4785) & VN_data_in(4785);
  VN797_in4 <= VN_sign_in(4786) & VN_data_in(4786);
  VN797_in5 <= VN_sign_in(4787) & VN_data_in(4787);
  VN798_in0 <= VN_sign_in(4788) & VN_data_in(4788);
  VN798_in1 <= VN_sign_in(4789) & VN_data_in(4789);
  VN798_in2 <= VN_sign_in(4790) & VN_data_in(4790);
  VN798_in3 <= VN_sign_in(4791) & VN_data_in(4791);
  VN798_in4 <= VN_sign_in(4792) & VN_data_in(4792);
  VN798_in5 <= VN_sign_in(4793) & VN_data_in(4793);
  VN799_in0 <= VN_sign_in(4794) & VN_data_in(4794);
  VN799_in1 <= VN_sign_in(4795) & VN_data_in(4795);
  VN799_in2 <= VN_sign_in(4796) & VN_data_in(4796);
  VN799_in3 <= VN_sign_in(4797) & VN_data_in(4797);
  VN799_in4 <= VN_sign_in(4798) & VN_data_in(4798);
  VN799_in5 <= VN_sign_in(4799) & VN_data_in(4799);
  VN800_in0 <= VN_sign_in(4800) & VN_data_in(4800);
  VN800_in1 <= VN_sign_in(4801) & VN_data_in(4801);
  VN800_in2 <= VN_sign_in(4802) & VN_data_in(4802);
  VN800_in3 <= VN_sign_in(4803) & VN_data_in(4803);
  VN800_in4 <= VN_sign_in(4804) & VN_data_in(4804);
  VN800_in5 <= VN_sign_in(4805) & VN_data_in(4805);
  VN801_in0 <= VN_sign_in(4806) & VN_data_in(4806);
  VN801_in1 <= VN_sign_in(4807) & VN_data_in(4807);
  VN801_in2 <= VN_sign_in(4808) & VN_data_in(4808);
  VN801_in3 <= VN_sign_in(4809) & VN_data_in(4809);
  VN801_in4 <= VN_sign_in(4810) & VN_data_in(4810);
  VN801_in5 <= VN_sign_in(4811) & VN_data_in(4811);
  VN802_in0 <= VN_sign_in(4812) & VN_data_in(4812);
  VN802_in1 <= VN_sign_in(4813) & VN_data_in(4813);
  VN802_in2 <= VN_sign_in(4814) & VN_data_in(4814);
  VN802_in3 <= VN_sign_in(4815) & VN_data_in(4815);
  VN802_in4 <= VN_sign_in(4816) & VN_data_in(4816);
  VN802_in5 <= VN_sign_in(4817) & VN_data_in(4817);
  VN803_in0 <= VN_sign_in(4818) & VN_data_in(4818);
  VN803_in1 <= VN_sign_in(4819) & VN_data_in(4819);
  VN803_in2 <= VN_sign_in(4820) & VN_data_in(4820);
  VN803_in3 <= VN_sign_in(4821) & VN_data_in(4821);
  VN803_in4 <= VN_sign_in(4822) & VN_data_in(4822);
  VN803_in5 <= VN_sign_in(4823) & VN_data_in(4823);
  VN804_in0 <= VN_sign_in(4824) & VN_data_in(4824);
  VN804_in1 <= VN_sign_in(4825) & VN_data_in(4825);
  VN804_in2 <= VN_sign_in(4826) & VN_data_in(4826);
  VN804_in3 <= VN_sign_in(4827) & VN_data_in(4827);
  VN804_in4 <= VN_sign_in(4828) & VN_data_in(4828);
  VN804_in5 <= VN_sign_in(4829) & VN_data_in(4829);
  VN805_in0 <= VN_sign_in(4830) & VN_data_in(4830);
  VN805_in1 <= VN_sign_in(4831) & VN_data_in(4831);
  VN805_in2 <= VN_sign_in(4832) & VN_data_in(4832);
  VN805_in3 <= VN_sign_in(4833) & VN_data_in(4833);
  VN805_in4 <= VN_sign_in(4834) & VN_data_in(4834);
  VN805_in5 <= VN_sign_in(4835) & VN_data_in(4835);
  VN806_in0 <= VN_sign_in(4836) & VN_data_in(4836);
  VN806_in1 <= VN_sign_in(4837) & VN_data_in(4837);
  VN806_in2 <= VN_sign_in(4838) & VN_data_in(4838);
  VN806_in3 <= VN_sign_in(4839) & VN_data_in(4839);
  VN806_in4 <= VN_sign_in(4840) & VN_data_in(4840);
  VN806_in5 <= VN_sign_in(4841) & VN_data_in(4841);
  VN807_in0 <= VN_sign_in(4842) & VN_data_in(4842);
  VN807_in1 <= VN_sign_in(4843) & VN_data_in(4843);
  VN807_in2 <= VN_sign_in(4844) & VN_data_in(4844);
  VN807_in3 <= VN_sign_in(4845) & VN_data_in(4845);
  VN807_in4 <= VN_sign_in(4846) & VN_data_in(4846);
  VN807_in5 <= VN_sign_in(4847) & VN_data_in(4847);
  VN808_in0 <= VN_sign_in(4848) & VN_data_in(4848);
  VN808_in1 <= VN_sign_in(4849) & VN_data_in(4849);
  VN808_in2 <= VN_sign_in(4850) & VN_data_in(4850);
  VN808_in3 <= VN_sign_in(4851) & VN_data_in(4851);
  VN808_in4 <= VN_sign_in(4852) & VN_data_in(4852);
  VN808_in5 <= VN_sign_in(4853) & VN_data_in(4853);
  VN809_in0 <= VN_sign_in(4854) & VN_data_in(4854);
  VN809_in1 <= VN_sign_in(4855) & VN_data_in(4855);
  VN809_in2 <= VN_sign_in(4856) & VN_data_in(4856);
  VN809_in3 <= VN_sign_in(4857) & VN_data_in(4857);
  VN809_in4 <= VN_sign_in(4858) & VN_data_in(4858);
  VN809_in5 <= VN_sign_in(4859) & VN_data_in(4859);
  VN810_in0 <= VN_sign_in(4860) & VN_data_in(4860);
  VN810_in1 <= VN_sign_in(4861) & VN_data_in(4861);
  VN810_in2 <= VN_sign_in(4862) & VN_data_in(4862);
  VN810_in3 <= VN_sign_in(4863) & VN_data_in(4863);
  VN810_in4 <= VN_sign_in(4864) & VN_data_in(4864);
  VN810_in5 <= VN_sign_in(4865) & VN_data_in(4865);
  VN811_in0 <= VN_sign_in(4866) & VN_data_in(4866);
  VN811_in1 <= VN_sign_in(4867) & VN_data_in(4867);
  VN811_in2 <= VN_sign_in(4868) & VN_data_in(4868);
  VN811_in3 <= VN_sign_in(4869) & VN_data_in(4869);
  VN811_in4 <= VN_sign_in(4870) & VN_data_in(4870);
  VN811_in5 <= VN_sign_in(4871) & VN_data_in(4871);
  VN812_in0 <= VN_sign_in(4872) & VN_data_in(4872);
  VN812_in1 <= VN_sign_in(4873) & VN_data_in(4873);
  VN812_in2 <= VN_sign_in(4874) & VN_data_in(4874);
  VN812_in3 <= VN_sign_in(4875) & VN_data_in(4875);
  VN812_in4 <= VN_sign_in(4876) & VN_data_in(4876);
  VN812_in5 <= VN_sign_in(4877) & VN_data_in(4877);
  VN813_in0 <= VN_sign_in(4878) & VN_data_in(4878);
  VN813_in1 <= VN_sign_in(4879) & VN_data_in(4879);
  VN813_in2 <= VN_sign_in(4880) & VN_data_in(4880);
  VN813_in3 <= VN_sign_in(4881) & VN_data_in(4881);
  VN813_in4 <= VN_sign_in(4882) & VN_data_in(4882);
  VN813_in5 <= VN_sign_in(4883) & VN_data_in(4883);
  VN814_in0 <= VN_sign_in(4884) & VN_data_in(4884);
  VN814_in1 <= VN_sign_in(4885) & VN_data_in(4885);
  VN814_in2 <= VN_sign_in(4886) & VN_data_in(4886);
  VN814_in3 <= VN_sign_in(4887) & VN_data_in(4887);
  VN814_in4 <= VN_sign_in(4888) & VN_data_in(4888);
  VN814_in5 <= VN_sign_in(4889) & VN_data_in(4889);
  VN815_in0 <= VN_sign_in(4890) & VN_data_in(4890);
  VN815_in1 <= VN_sign_in(4891) & VN_data_in(4891);
  VN815_in2 <= VN_sign_in(4892) & VN_data_in(4892);
  VN815_in3 <= VN_sign_in(4893) & VN_data_in(4893);
  VN815_in4 <= VN_sign_in(4894) & VN_data_in(4894);
  VN815_in5 <= VN_sign_in(4895) & VN_data_in(4895);
  VN816_in0 <= VN_sign_in(4896) & VN_data_in(4896);
  VN816_in1 <= VN_sign_in(4897) & VN_data_in(4897);
  VN816_in2 <= VN_sign_in(4898) & VN_data_in(4898);
  VN816_in3 <= VN_sign_in(4899) & VN_data_in(4899);
  VN816_in4 <= VN_sign_in(4900) & VN_data_in(4900);
  VN816_in5 <= VN_sign_in(4901) & VN_data_in(4901);
  VN817_in0 <= VN_sign_in(4902) & VN_data_in(4902);
  VN817_in1 <= VN_sign_in(4903) & VN_data_in(4903);
  VN817_in2 <= VN_sign_in(4904) & VN_data_in(4904);
  VN817_in3 <= VN_sign_in(4905) & VN_data_in(4905);
  VN817_in4 <= VN_sign_in(4906) & VN_data_in(4906);
  VN817_in5 <= VN_sign_in(4907) & VN_data_in(4907);
  VN818_in0 <= VN_sign_in(4908) & VN_data_in(4908);
  VN818_in1 <= VN_sign_in(4909) & VN_data_in(4909);
  VN818_in2 <= VN_sign_in(4910) & VN_data_in(4910);
  VN818_in3 <= VN_sign_in(4911) & VN_data_in(4911);
  VN818_in4 <= VN_sign_in(4912) & VN_data_in(4912);
  VN818_in5 <= VN_sign_in(4913) & VN_data_in(4913);
  VN819_in0 <= VN_sign_in(4914) & VN_data_in(4914);
  VN819_in1 <= VN_sign_in(4915) & VN_data_in(4915);
  VN819_in2 <= VN_sign_in(4916) & VN_data_in(4916);
  VN819_in3 <= VN_sign_in(4917) & VN_data_in(4917);
  VN819_in4 <= VN_sign_in(4918) & VN_data_in(4918);
  VN819_in5 <= VN_sign_in(4919) & VN_data_in(4919);
  VN820_in0 <= VN_sign_in(4920) & VN_data_in(4920);
  VN820_in1 <= VN_sign_in(4921) & VN_data_in(4921);
  VN820_in2 <= VN_sign_in(4922) & VN_data_in(4922);
  VN820_in3 <= VN_sign_in(4923) & VN_data_in(4923);
  VN820_in4 <= VN_sign_in(4924) & VN_data_in(4924);
  VN820_in5 <= VN_sign_in(4925) & VN_data_in(4925);
  VN821_in0 <= VN_sign_in(4926) & VN_data_in(4926);
  VN821_in1 <= VN_sign_in(4927) & VN_data_in(4927);
  VN821_in2 <= VN_sign_in(4928) & VN_data_in(4928);
  VN821_in3 <= VN_sign_in(4929) & VN_data_in(4929);
  VN821_in4 <= VN_sign_in(4930) & VN_data_in(4930);
  VN821_in5 <= VN_sign_in(4931) & VN_data_in(4931);
  VN822_in0 <= VN_sign_in(4932) & VN_data_in(4932);
  VN822_in1 <= VN_sign_in(4933) & VN_data_in(4933);
  VN822_in2 <= VN_sign_in(4934) & VN_data_in(4934);
  VN822_in3 <= VN_sign_in(4935) & VN_data_in(4935);
  VN822_in4 <= VN_sign_in(4936) & VN_data_in(4936);
  VN822_in5 <= VN_sign_in(4937) & VN_data_in(4937);
  VN823_in0 <= VN_sign_in(4938) & VN_data_in(4938);
  VN823_in1 <= VN_sign_in(4939) & VN_data_in(4939);
  VN823_in2 <= VN_sign_in(4940) & VN_data_in(4940);
  VN823_in3 <= VN_sign_in(4941) & VN_data_in(4941);
  VN823_in4 <= VN_sign_in(4942) & VN_data_in(4942);
  VN823_in5 <= VN_sign_in(4943) & VN_data_in(4943);
  VN824_in0 <= VN_sign_in(4944) & VN_data_in(4944);
  VN824_in1 <= VN_sign_in(4945) & VN_data_in(4945);
  VN824_in2 <= VN_sign_in(4946) & VN_data_in(4946);
  VN824_in3 <= VN_sign_in(4947) & VN_data_in(4947);
  VN824_in4 <= VN_sign_in(4948) & VN_data_in(4948);
  VN824_in5 <= VN_sign_in(4949) & VN_data_in(4949);
  VN825_in0 <= VN_sign_in(4950) & VN_data_in(4950);
  VN825_in1 <= VN_sign_in(4951) & VN_data_in(4951);
  VN825_in2 <= VN_sign_in(4952) & VN_data_in(4952);
  VN825_in3 <= VN_sign_in(4953) & VN_data_in(4953);
  VN825_in4 <= VN_sign_in(4954) & VN_data_in(4954);
  VN825_in5 <= VN_sign_in(4955) & VN_data_in(4955);
  VN826_in0 <= VN_sign_in(4956) & VN_data_in(4956);
  VN826_in1 <= VN_sign_in(4957) & VN_data_in(4957);
  VN826_in2 <= VN_sign_in(4958) & VN_data_in(4958);
  VN826_in3 <= VN_sign_in(4959) & VN_data_in(4959);
  VN826_in4 <= VN_sign_in(4960) & VN_data_in(4960);
  VN826_in5 <= VN_sign_in(4961) & VN_data_in(4961);
  VN827_in0 <= VN_sign_in(4962) & VN_data_in(4962);
  VN827_in1 <= VN_sign_in(4963) & VN_data_in(4963);
  VN827_in2 <= VN_sign_in(4964) & VN_data_in(4964);
  VN827_in3 <= VN_sign_in(4965) & VN_data_in(4965);
  VN827_in4 <= VN_sign_in(4966) & VN_data_in(4966);
  VN827_in5 <= VN_sign_in(4967) & VN_data_in(4967);
  VN828_in0 <= VN_sign_in(4968) & VN_data_in(4968);
  VN828_in1 <= VN_sign_in(4969) & VN_data_in(4969);
  VN828_in2 <= VN_sign_in(4970) & VN_data_in(4970);
  VN828_in3 <= VN_sign_in(4971) & VN_data_in(4971);
  VN828_in4 <= VN_sign_in(4972) & VN_data_in(4972);
  VN828_in5 <= VN_sign_in(4973) & VN_data_in(4973);
  VN829_in0 <= VN_sign_in(4974) & VN_data_in(4974);
  VN829_in1 <= VN_sign_in(4975) & VN_data_in(4975);
  VN829_in2 <= VN_sign_in(4976) & VN_data_in(4976);
  VN829_in3 <= VN_sign_in(4977) & VN_data_in(4977);
  VN829_in4 <= VN_sign_in(4978) & VN_data_in(4978);
  VN829_in5 <= VN_sign_in(4979) & VN_data_in(4979);
  VN830_in0 <= VN_sign_in(4980) & VN_data_in(4980);
  VN830_in1 <= VN_sign_in(4981) & VN_data_in(4981);
  VN830_in2 <= VN_sign_in(4982) & VN_data_in(4982);
  VN830_in3 <= VN_sign_in(4983) & VN_data_in(4983);
  VN830_in4 <= VN_sign_in(4984) & VN_data_in(4984);
  VN830_in5 <= VN_sign_in(4985) & VN_data_in(4985);
  VN831_in0 <= VN_sign_in(4986) & VN_data_in(4986);
  VN831_in1 <= VN_sign_in(4987) & VN_data_in(4987);
  VN831_in2 <= VN_sign_in(4988) & VN_data_in(4988);
  VN831_in3 <= VN_sign_in(4989) & VN_data_in(4989);
  VN831_in4 <= VN_sign_in(4990) & VN_data_in(4990);
  VN831_in5 <= VN_sign_in(4991) & VN_data_in(4991);
  VN832_in0 <= VN_sign_in(4992) & VN_data_in(4992);
  VN832_in1 <= VN_sign_in(4993) & VN_data_in(4993);
  VN832_in2 <= VN_sign_in(4994) & VN_data_in(4994);
  VN832_in3 <= VN_sign_in(4995) & VN_data_in(4995);
  VN832_in4 <= VN_sign_in(4996) & VN_data_in(4996);
  VN832_in5 <= VN_sign_in(4997) & VN_data_in(4997);
  VN833_in0 <= VN_sign_in(4998) & VN_data_in(4998);
  VN833_in1 <= VN_sign_in(4999) & VN_data_in(4999);
  VN833_in2 <= VN_sign_in(5000) & VN_data_in(5000);
  VN833_in3 <= VN_sign_in(5001) & VN_data_in(5001);
  VN833_in4 <= VN_sign_in(5002) & VN_data_in(5002);
  VN833_in5 <= VN_sign_in(5003) & VN_data_in(5003);
  VN834_in0 <= VN_sign_in(5004) & VN_data_in(5004);
  VN834_in1 <= VN_sign_in(5005) & VN_data_in(5005);
  VN834_in2 <= VN_sign_in(5006) & VN_data_in(5006);
  VN834_in3 <= VN_sign_in(5007) & VN_data_in(5007);
  VN834_in4 <= VN_sign_in(5008) & VN_data_in(5008);
  VN834_in5 <= VN_sign_in(5009) & VN_data_in(5009);
  VN835_in0 <= VN_sign_in(5010) & VN_data_in(5010);
  VN835_in1 <= VN_sign_in(5011) & VN_data_in(5011);
  VN835_in2 <= VN_sign_in(5012) & VN_data_in(5012);
  VN835_in3 <= VN_sign_in(5013) & VN_data_in(5013);
  VN835_in4 <= VN_sign_in(5014) & VN_data_in(5014);
  VN835_in5 <= VN_sign_in(5015) & VN_data_in(5015);
  VN836_in0 <= VN_sign_in(5016) & VN_data_in(5016);
  VN836_in1 <= VN_sign_in(5017) & VN_data_in(5017);
  VN836_in2 <= VN_sign_in(5018) & VN_data_in(5018);
  VN836_in3 <= VN_sign_in(5019) & VN_data_in(5019);
  VN836_in4 <= VN_sign_in(5020) & VN_data_in(5020);
  VN836_in5 <= VN_sign_in(5021) & VN_data_in(5021);
  VN837_in0 <= VN_sign_in(5022) & VN_data_in(5022);
  VN837_in1 <= VN_sign_in(5023) & VN_data_in(5023);
  VN837_in2 <= VN_sign_in(5024) & VN_data_in(5024);
  VN837_in3 <= VN_sign_in(5025) & VN_data_in(5025);
  VN837_in4 <= VN_sign_in(5026) & VN_data_in(5026);
  VN837_in5 <= VN_sign_in(5027) & VN_data_in(5027);
  VN838_in0 <= VN_sign_in(5028) & VN_data_in(5028);
  VN838_in1 <= VN_sign_in(5029) & VN_data_in(5029);
  VN838_in2 <= VN_sign_in(5030) & VN_data_in(5030);
  VN838_in3 <= VN_sign_in(5031) & VN_data_in(5031);
  VN838_in4 <= VN_sign_in(5032) & VN_data_in(5032);
  VN838_in5 <= VN_sign_in(5033) & VN_data_in(5033);
  VN839_in0 <= VN_sign_in(5034) & VN_data_in(5034);
  VN839_in1 <= VN_sign_in(5035) & VN_data_in(5035);
  VN839_in2 <= VN_sign_in(5036) & VN_data_in(5036);
  VN839_in3 <= VN_sign_in(5037) & VN_data_in(5037);
  VN839_in4 <= VN_sign_in(5038) & VN_data_in(5038);
  VN839_in5 <= VN_sign_in(5039) & VN_data_in(5039);
  VN840_in0 <= VN_sign_in(5040) & VN_data_in(5040);
  VN840_in1 <= VN_sign_in(5041) & VN_data_in(5041);
  VN840_in2 <= VN_sign_in(5042) & VN_data_in(5042);
  VN840_in3 <= VN_sign_in(5043) & VN_data_in(5043);
  VN840_in4 <= VN_sign_in(5044) & VN_data_in(5044);
  VN840_in5 <= VN_sign_in(5045) & VN_data_in(5045);
  VN841_in0 <= VN_sign_in(5046) & VN_data_in(5046);
  VN841_in1 <= VN_sign_in(5047) & VN_data_in(5047);
  VN841_in2 <= VN_sign_in(5048) & VN_data_in(5048);
  VN841_in3 <= VN_sign_in(5049) & VN_data_in(5049);
  VN841_in4 <= VN_sign_in(5050) & VN_data_in(5050);
  VN841_in5 <= VN_sign_in(5051) & VN_data_in(5051);
  VN842_in0 <= VN_sign_in(5052) & VN_data_in(5052);
  VN842_in1 <= VN_sign_in(5053) & VN_data_in(5053);
  VN842_in2 <= VN_sign_in(5054) & VN_data_in(5054);
  VN842_in3 <= VN_sign_in(5055) & VN_data_in(5055);
  VN842_in4 <= VN_sign_in(5056) & VN_data_in(5056);
  VN842_in5 <= VN_sign_in(5057) & VN_data_in(5057);
  VN843_in0 <= VN_sign_in(5058) & VN_data_in(5058);
  VN843_in1 <= VN_sign_in(5059) & VN_data_in(5059);
  VN843_in2 <= VN_sign_in(5060) & VN_data_in(5060);
  VN843_in3 <= VN_sign_in(5061) & VN_data_in(5061);
  VN843_in4 <= VN_sign_in(5062) & VN_data_in(5062);
  VN843_in5 <= VN_sign_in(5063) & VN_data_in(5063);
  VN844_in0 <= VN_sign_in(5064) & VN_data_in(5064);
  VN844_in1 <= VN_sign_in(5065) & VN_data_in(5065);
  VN844_in2 <= VN_sign_in(5066) & VN_data_in(5066);
  VN844_in3 <= VN_sign_in(5067) & VN_data_in(5067);
  VN844_in4 <= VN_sign_in(5068) & VN_data_in(5068);
  VN844_in5 <= VN_sign_in(5069) & VN_data_in(5069);
  VN845_in0 <= VN_sign_in(5070) & VN_data_in(5070);
  VN845_in1 <= VN_sign_in(5071) & VN_data_in(5071);
  VN845_in2 <= VN_sign_in(5072) & VN_data_in(5072);
  VN845_in3 <= VN_sign_in(5073) & VN_data_in(5073);
  VN845_in4 <= VN_sign_in(5074) & VN_data_in(5074);
  VN845_in5 <= VN_sign_in(5075) & VN_data_in(5075);
  VN846_in0 <= VN_sign_in(5076) & VN_data_in(5076);
  VN846_in1 <= VN_sign_in(5077) & VN_data_in(5077);
  VN846_in2 <= VN_sign_in(5078) & VN_data_in(5078);
  VN846_in3 <= VN_sign_in(5079) & VN_data_in(5079);
  VN846_in4 <= VN_sign_in(5080) & VN_data_in(5080);
  VN846_in5 <= VN_sign_in(5081) & VN_data_in(5081);
  VN847_in0 <= VN_sign_in(5082) & VN_data_in(5082);
  VN847_in1 <= VN_sign_in(5083) & VN_data_in(5083);
  VN847_in2 <= VN_sign_in(5084) & VN_data_in(5084);
  VN847_in3 <= VN_sign_in(5085) & VN_data_in(5085);
  VN847_in4 <= VN_sign_in(5086) & VN_data_in(5086);
  VN847_in5 <= VN_sign_in(5087) & VN_data_in(5087);
  VN848_in0 <= VN_sign_in(5088) & VN_data_in(5088);
  VN848_in1 <= VN_sign_in(5089) & VN_data_in(5089);
  VN848_in2 <= VN_sign_in(5090) & VN_data_in(5090);
  VN848_in3 <= VN_sign_in(5091) & VN_data_in(5091);
  VN848_in4 <= VN_sign_in(5092) & VN_data_in(5092);
  VN848_in5 <= VN_sign_in(5093) & VN_data_in(5093);
  VN849_in0 <= VN_sign_in(5094) & VN_data_in(5094);
  VN849_in1 <= VN_sign_in(5095) & VN_data_in(5095);
  VN849_in2 <= VN_sign_in(5096) & VN_data_in(5096);
  VN849_in3 <= VN_sign_in(5097) & VN_data_in(5097);
  VN849_in4 <= VN_sign_in(5098) & VN_data_in(5098);
  VN849_in5 <= VN_sign_in(5099) & VN_data_in(5099);
  VN850_in0 <= VN_sign_in(5100) & VN_data_in(5100);
  VN850_in1 <= VN_sign_in(5101) & VN_data_in(5101);
  VN850_in2 <= VN_sign_in(5102) & VN_data_in(5102);
  VN850_in3 <= VN_sign_in(5103) & VN_data_in(5103);
  VN850_in4 <= VN_sign_in(5104) & VN_data_in(5104);
  VN850_in5 <= VN_sign_in(5105) & VN_data_in(5105);
  VN851_in0 <= VN_sign_in(5106) & VN_data_in(5106);
  VN851_in1 <= VN_sign_in(5107) & VN_data_in(5107);
  VN851_in2 <= VN_sign_in(5108) & VN_data_in(5108);
  VN851_in3 <= VN_sign_in(5109) & VN_data_in(5109);
  VN851_in4 <= VN_sign_in(5110) & VN_data_in(5110);
  VN851_in5 <= VN_sign_in(5111) & VN_data_in(5111);
  VN852_in0 <= VN_sign_in(5112) & VN_data_in(5112);
  VN852_in1 <= VN_sign_in(5113) & VN_data_in(5113);
  VN852_in2 <= VN_sign_in(5114) & VN_data_in(5114);
  VN852_in3 <= VN_sign_in(5115) & VN_data_in(5115);
  VN852_in4 <= VN_sign_in(5116) & VN_data_in(5116);
  VN852_in5 <= VN_sign_in(5117) & VN_data_in(5117);
  VN853_in0 <= VN_sign_in(5118) & VN_data_in(5118);
  VN853_in1 <= VN_sign_in(5119) & VN_data_in(5119);
  VN853_in2 <= VN_sign_in(5120) & VN_data_in(5120);
  VN853_in3 <= VN_sign_in(5121) & VN_data_in(5121);
  VN853_in4 <= VN_sign_in(5122) & VN_data_in(5122);
  VN853_in5 <= VN_sign_in(5123) & VN_data_in(5123);
  VN854_in0 <= VN_sign_in(5124) & VN_data_in(5124);
  VN854_in1 <= VN_sign_in(5125) & VN_data_in(5125);
  VN854_in2 <= VN_sign_in(5126) & VN_data_in(5126);
  VN854_in3 <= VN_sign_in(5127) & VN_data_in(5127);
  VN854_in4 <= VN_sign_in(5128) & VN_data_in(5128);
  VN854_in5 <= VN_sign_in(5129) & VN_data_in(5129);
  VN855_in0 <= VN_sign_in(5130) & VN_data_in(5130);
  VN855_in1 <= VN_sign_in(5131) & VN_data_in(5131);
  VN855_in2 <= VN_sign_in(5132) & VN_data_in(5132);
  VN855_in3 <= VN_sign_in(5133) & VN_data_in(5133);
  VN855_in4 <= VN_sign_in(5134) & VN_data_in(5134);
  VN855_in5 <= VN_sign_in(5135) & VN_data_in(5135);
  VN856_in0 <= VN_sign_in(5136) & VN_data_in(5136);
  VN856_in1 <= VN_sign_in(5137) & VN_data_in(5137);
  VN856_in2 <= VN_sign_in(5138) & VN_data_in(5138);
  VN856_in3 <= VN_sign_in(5139) & VN_data_in(5139);
  VN856_in4 <= VN_sign_in(5140) & VN_data_in(5140);
  VN856_in5 <= VN_sign_in(5141) & VN_data_in(5141);
  VN857_in0 <= VN_sign_in(5142) & VN_data_in(5142);
  VN857_in1 <= VN_sign_in(5143) & VN_data_in(5143);
  VN857_in2 <= VN_sign_in(5144) & VN_data_in(5144);
  VN857_in3 <= VN_sign_in(5145) & VN_data_in(5145);
  VN857_in4 <= VN_sign_in(5146) & VN_data_in(5146);
  VN857_in5 <= VN_sign_in(5147) & VN_data_in(5147);
  VN858_in0 <= VN_sign_in(5148) & VN_data_in(5148);
  VN858_in1 <= VN_sign_in(5149) & VN_data_in(5149);
  VN858_in2 <= VN_sign_in(5150) & VN_data_in(5150);
  VN858_in3 <= VN_sign_in(5151) & VN_data_in(5151);
  VN858_in4 <= VN_sign_in(5152) & VN_data_in(5152);
  VN858_in5 <= VN_sign_in(5153) & VN_data_in(5153);
  VN859_in0 <= VN_sign_in(5154) & VN_data_in(5154);
  VN859_in1 <= VN_sign_in(5155) & VN_data_in(5155);
  VN859_in2 <= VN_sign_in(5156) & VN_data_in(5156);
  VN859_in3 <= VN_sign_in(5157) & VN_data_in(5157);
  VN859_in4 <= VN_sign_in(5158) & VN_data_in(5158);
  VN859_in5 <= VN_sign_in(5159) & VN_data_in(5159);
  VN860_in0 <= VN_sign_in(5160) & VN_data_in(5160);
  VN860_in1 <= VN_sign_in(5161) & VN_data_in(5161);
  VN860_in2 <= VN_sign_in(5162) & VN_data_in(5162);
  VN860_in3 <= VN_sign_in(5163) & VN_data_in(5163);
  VN860_in4 <= VN_sign_in(5164) & VN_data_in(5164);
  VN860_in5 <= VN_sign_in(5165) & VN_data_in(5165);
  VN861_in0 <= VN_sign_in(5166) & VN_data_in(5166);
  VN861_in1 <= VN_sign_in(5167) & VN_data_in(5167);
  VN861_in2 <= VN_sign_in(5168) & VN_data_in(5168);
  VN861_in3 <= VN_sign_in(5169) & VN_data_in(5169);
  VN861_in4 <= VN_sign_in(5170) & VN_data_in(5170);
  VN861_in5 <= VN_sign_in(5171) & VN_data_in(5171);
  VN862_in0 <= VN_sign_in(5172) & VN_data_in(5172);
  VN862_in1 <= VN_sign_in(5173) & VN_data_in(5173);
  VN862_in2 <= VN_sign_in(5174) & VN_data_in(5174);
  VN862_in3 <= VN_sign_in(5175) & VN_data_in(5175);
  VN862_in4 <= VN_sign_in(5176) & VN_data_in(5176);
  VN862_in5 <= VN_sign_in(5177) & VN_data_in(5177);
  VN863_in0 <= VN_sign_in(5178) & VN_data_in(5178);
  VN863_in1 <= VN_sign_in(5179) & VN_data_in(5179);
  VN863_in2 <= VN_sign_in(5180) & VN_data_in(5180);
  VN863_in3 <= VN_sign_in(5181) & VN_data_in(5181);
  VN863_in4 <= VN_sign_in(5182) & VN_data_in(5182);
  VN863_in5 <= VN_sign_in(5183) & VN_data_in(5183);
  VN864_in0 <= VN_sign_in(5184) & VN_data_in(5184);
  VN864_in1 <= VN_sign_in(5185) & VN_data_in(5185);
  VN864_in2 <= VN_sign_in(5186) & VN_data_in(5186);
  VN864_in3 <= VN_sign_in(5187) & VN_data_in(5187);
  VN864_in4 <= VN_sign_in(5188) & VN_data_in(5188);
  VN864_in5 <= VN_sign_in(5189) & VN_data_in(5189);
  VN865_in0 <= VN_sign_in(5190) & VN_data_in(5190);
  VN865_in1 <= VN_sign_in(5191) & VN_data_in(5191);
  VN865_in2 <= VN_sign_in(5192) & VN_data_in(5192);
  VN865_in3 <= VN_sign_in(5193) & VN_data_in(5193);
  VN865_in4 <= VN_sign_in(5194) & VN_data_in(5194);
  VN865_in5 <= VN_sign_in(5195) & VN_data_in(5195);
  VN866_in0 <= VN_sign_in(5196) & VN_data_in(5196);
  VN866_in1 <= VN_sign_in(5197) & VN_data_in(5197);
  VN866_in2 <= VN_sign_in(5198) & VN_data_in(5198);
  VN866_in3 <= VN_sign_in(5199) & VN_data_in(5199);
  VN866_in4 <= VN_sign_in(5200) & VN_data_in(5200);
  VN866_in5 <= VN_sign_in(5201) & VN_data_in(5201);
  VN867_in0 <= VN_sign_in(5202) & VN_data_in(5202);
  VN867_in1 <= VN_sign_in(5203) & VN_data_in(5203);
  VN867_in2 <= VN_sign_in(5204) & VN_data_in(5204);
  VN867_in3 <= VN_sign_in(5205) & VN_data_in(5205);
  VN867_in4 <= VN_sign_in(5206) & VN_data_in(5206);
  VN867_in5 <= VN_sign_in(5207) & VN_data_in(5207);
  VN868_in0 <= VN_sign_in(5208) & VN_data_in(5208);
  VN868_in1 <= VN_sign_in(5209) & VN_data_in(5209);
  VN868_in2 <= VN_sign_in(5210) & VN_data_in(5210);
  VN868_in3 <= VN_sign_in(5211) & VN_data_in(5211);
  VN868_in4 <= VN_sign_in(5212) & VN_data_in(5212);
  VN868_in5 <= VN_sign_in(5213) & VN_data_in(5213);
  VN869_in0 <= VN_sign_in(5214) & VN_data_in(5214);
  VN869_in1 <= VN_sign_in(5215) & VN_data_in(5215);
  VN869_in2 <= VN_sign_in(5216) & VN_data_in(5216);
  VN869_in3 <= VN_sign_in(5217) & VN_data_in(5217);
  VN869_in4 <= VN_sign_in(5218) & VN_data_in(5218);
  VN869_in5 <= VN_sign_in(5219) & VN_data_in(5219);
  VN870_in0 <= VN_sign_in(5220) & VN_data_in(5220);
  VN870_in1 <= VN_sign_in(5221) & VN_data_in(5221);
  VN870_in2 <= VN_sign_in(5222) & VN_data_in(5222);
  VN870_in3 <= VN_sign_in(5223) & VN_data_in(5223);
  VN870_in4 <= VN_sign_in(5224) & VN_data_in(5224);
  VN870_in5 <= VN_sign_in(5225) & VN_data_in(5225);
  VN871_in0 <= VN_sign_in(5226) & VN_data_in(5226);
  VN871_in1 <= VN_sign_in(5227) & VN_data_in(5227);
  VN871_in2 <= VN_sign_in(5228) & VN_data_in(5228);
  VN871_in3 <= VN_sign_in(5229) & VN_data_in(5229);
  VN871_in4 <= VN_sign_in(5230) & VN_data_in(5230);
  VN871_in5 <= VN_sign_in(5231) & VN_data_in(5231);
  VN872_in0 <= VN_sign_in(5232) & VN_data_in(5232);
  VN872_in1 <= VN_sign_in(5233) & VN_data_in(5233);
  VN872_in2 <= VN_sign_in(5234) & VN_data_in(5234);
  VN872_in3 <= VN_sign_in(5235) & VN_data_in(5235);
  VN872_in4 <= VN_sign_in(5236) & VN_data_in(5236);
  VN872_in5 <= VN_sign_in(5237) & VN_data_in(5237);
  VN873_in0 <= VN_sign_in(5238) & VN_data_in(5238);
  VN873_in1 <= VN_sign_in(5239) & VN_data_in(5239);
  VN873_in2 <= VN_sign_in(5240) & VN_data_in(5240);
  VN873_in3 <= VN_sign_in(5241) & VN_data_in(5241);
  VN873_in4 <= VN_sign_in(5242) & VN_data_in(5242);
  VN873_in5 <= VN_sign_in(5243) & VN_data_in(5243);
  VN874_in0 <= VN_sign_in(5244) & VN_data_in(5244);
  VN874_in1 <= VN_sign_in(5245) & VN_data_in(5245);
  VN874_in2 <= VN_sign_in(5246) & VN_data_in(5246);
  VN874_in3 <= VN_sign_in(5247) & VN_data_in(5247);
  VN874_in4 <= VN_sign_in(5248) & VN_data_in(5248);
  VN874_in5 <= VN_sign_in(5249) & VN_data_in(5249);
  VN875_in0 <= VN_sign_in(5250) & VN_data_in(5250);
  VN875_in1 <= VN_sign_in(5251) & VN_data_in(5251);
  VN875_in2 <= VN_sign_in(5252) & VN_data_in(5252);
  VN875_in3 <= VN_sign_in(5253) & VN_data_in(5253);
  VN875_in4 <= VN_sign_in(5254) & VN_data_in(5254);
  VN875_in5 <= VN_sign_in(5255) & VN_data_in(5255);
  VN876_in0 <= VN_sign_in(5256) & VN_data_in(5256);
  VN876_in1 <= VN_sign_in(5257) & VN_data_in(5257);
  VN876_in2 <= VN_sign_in(5258) & VN_data_in(5258);
  VN876_in3 <= VN_sign_in(5259) & VN_data_in(5259);
  VN876_in4 <= VN_sign_in(5260) & VN_data_in(5260);
  VN876_in5 <= VN_sign_in(5261) & VN_data_in(5261);
  VN877_in0 <= VN_sign_in(5262) & VN_data_in(5262);
  VN877_in1 <= VN_sign_in(5263) & VN_data_in(5263);
  VN877_in2 <= VN_sign_in(5264) & VN_data_in(5264);
  VN877_in3 <= VN_sign_in(5265) & VN_data_in(5265);
  VN877_in4 <= VN_sign_in(5266) & VN_data_in(5266);
  VN877_in5 <= VN_sign_in(5267) & VN_data_in(5267);
  VN878_in0 <= VN_sign_in(5268) & VN_data_in(5268);
  VN878_in1 <= VN_sign_in(5269) & VN_data_in(5269);
  VN878_in2 <= VN_sign_in(5270) & VN_data_in(5270);
  VN878_in3 <= VN_sign_in(5271) & VN_data_in(5271);
  VN878_in4 <= VN_sign_in(5272) & VN_data_in(5272);
  VN878_in5 <= VN_sign_in(5273) & VN_data_in(5273);
  VN879_in0 <= VN_sign_in(5274) & VN_data_in(5274);
  VN879_in1 <= VN_sign_in(5275) & VN_data_in(5275);
  VN879_in2 <= VN_sign_in(5276) & VN_data_in(5276);
  VN879_in3 <= VN_sign_in(5277) & VN_data_in(5277);
  VN879_in4 <= VN_sign_in(5278) & VN_data_in(5278);
  VN879_in5 <= VN_sign_in(5279) & VN_data_in(5279);
  VN880_in0 <= VN_sign_in(5280) & VN_data_in(5280);
  VN880_in1 <= VN_sign_in(5281) & VN_data_in(5281);
  VN880_in2 <= VN_sign_in(5282) & VN_data_in(5282);
  VN880_in3 <= VN_sign_in(5283) & VN_data_in(5283);
  VN880_in4 <= VN_sign_in(5284) & VN_data_in(5284);
  VN880_in5 <= VN_sign_in(5285) & VN_data_in(5285);
  VN881_in0 <= VN_sign_in(5286) & VN_data_in(5286);
  VN881_in1 <= VN_sign_in(5287) & VN_data_in(5287);
  VN881_in2 <= VN_sign_in(5288) & VN_data_in(5288);
  VN881_in3 <= VN_sign_in(5289) & VN_data_in(5289);
  VN881_in4 <= VN_sign_in(5290) & VN_data_in(5290);
  VN881_in5 <= VN_sign_in(5291) & VN_data_in(5291);
  VN882_in0 <= VN_sign_in(5292) & VN_data_in(5292);
  VN882_in1 <= VN_sign_in(5293) & VN_data_in(5293);
  VN882_in2 <= VN_sign_in(5294) & VN_data_in(5294);
  VN882_in3 <= VN_sign_in(5295) & VN_data_in(5295);
  VN882_in4 <= VN_sign_in(5296) & VN_data_in(5296);
  VN882_in5 <= VN_sign_in(5297) & VN_data_in(5297);
  VN883_in0 <= VN_sign_in(5298) & VN_data_in(5298);
  VN883_in1 <= VN_sign_in(5299) & VN_data_in(5299);
  VN883_in2 <= VN_sign_in(5300) & VN_data_in(5300);
  VN883_in3 <= VN_sign_in(5301) & VN_data_in(5301);
  VN883_in4 <= VN_sign_in(5302) & VN_data_in(5302);
  VN883_in5 <= VN_sign_in(5303) & VN_data_in(5303);
  VN884_in0 <= VN_sign_in(5304) & VN_data_in(5304);
  VN884_in1 <= VN_sign_in(5305) & VN_data_in(5305);
  VN884_in2 <= VN_sign_in(5306) & VN_data_in(5306);
  VN884_in3 <= VN_sign_in(5307) & VN_data_in(5307);
  VN884_in4 <= VN_sign_in(5308) & VN_data_in(5308);
  VN884_in5 <= VN_sign_in(5309) & VN_data_in(5309);
  VN885_in0 <= VN_sign_in(5310) & VN_data_in(5310);
  VN885_in1 <= VN_sign_in(5311) & VN_data_in(5311);
  VN885_in2 <= VN_sign_in(5312) & VN_data_in(5312);
  VN885_in3 <= VN_sign_in(5313) & VN_data_in(5313);
  VN885_in4 <= VN_sign_in(5314) & VN_data_in(5314);
  VN885_in5 <= VN_sign_in(5315) & VN_data_in(5315);
  VN886_in0 <= VN_sign_in(5316) & VN_data_in(5316);
  VN886_in1 <= VN_sign_in(5317) & VN_data_in(5317);
  VN886_in2 <= VN_sign_in(5318) & VN_data_in(5318);
  VN886_in3 <= VN_sign_in(5319) & VN_data_in(5319);
  VN886_in4 <= VN_sign_in(5320) & VN_data_in(5320);
  VN886_in5 <= VN_sign_in(5321) & VN_data_in(5321);
  VN887_in0 <= VN_sign_in(5322) & VN_data_in(5322);
  VN887_in1 <= VN_sign_in(5323) & VN_data_in(5323);
  VN887_in2 <= VN_sign_in(5324) & VN_data_in(5324);
  VN887_in3 <= VN_sign_in(5325) & VN_data_in(5325);
  VN887_in4 <= VN_sign_in(5326) & VN_data_in(5326);
  VN887_in5 <= VN_sign_in(5327) & VN_data_in(5327);
  VN888_in0 <= VN_sign_in(5328) & VN_data_in(5328);
  VN888_in1 <= VN_sign_in(5329) & VN_data_in(5329);
  VN888_in2 <= VN_sign_in(5330) & VN_data_in(5330);
  VN888_in3 <= VN_sign_in(5331) & VN_data_in(5331);
  VN888_in4 <= VN_sign_in(5332) & VN_data_in(5332);
  VN888_in5 <= VN_sign_in(5333) & VN_data_in(5333);
  VN889_in0 <= VN_sign_in(5334) & VN_data_in(5334);
  VN889_in1 <= VN_sign_in(5335) & VN_data_in(5335);
  VN889_in2 <= VN_sign_in(5336) & VN_data_in(5336);
  VN889_in3 <= VN_sign_in(5337) & VN_data_in(5337);
  VN889_in4 <= VN_sign_in(5338) & VN_data_in(5338);
  VN889_in5 <= VN_sign_in(5339) & VN_data_in(5339);
  VN890_in0 <= VN_sign_in(5340) & VN_data_in(5340);
  VN890_in1 <= VN_sign_in(5341) & VN_data_in(5341);
  VN890_in2 <= VN_sign_in(5342) & VN_data_in(5342);
  VN890_in3 <= VN_sign_in(5343) & VN_data_in(5343);
  VN890_in4 <= VN_sign_in(5344) & VN_data_in(5344);
  VN890_in5 <= VN_sign_in(5345) & VN_data_in(5345);
  VN891_in0 <= VN_sign_in(5346) & VN_data_in(5346);
  VN891_in1 <= VN_sign_in(5347) & VN_data_in(5347);
  VN891_in2 <= VN_sign_in(5348) & VN_data_in(5348);
  VN891_in3 <= VN_sign_in(5349) & VN_data_in(5349);
  VN891_in4 <= VN_sign_in(5350) & VN_data_in(5350);
  VN891_in5 <= VN_sign_in(5351) & VN_data_in(5351);
  VN892_in0 <= VN_sign_in(5352) & VN_data_in(5352);
  VN892_in1 <= VN_sign_in(5353) & VN_data_in(5353);
  VN892_in2 <= VN_sign_in(5354) & VN_data_in(5354);
  VN892_in3 <= VN_sign_in(5355) & VN_data_in(5355);
  VN892_in4 <= VN_sign_in(5356) & VN_data_in(5356);
  VN892_in5 <= VN_sign_in(5357) & VN_data_in(5357);
  VN893_in0 <= VN_sign_in(5358) & VN_data_in(5358);
  VN893_in1 <= VN_sign_in(5359) & VN_data_in(5359);
  VN893_in2 <= VN_sign_in(5360) & VN_data_in(5360);
  VN893_in3 <= VN_sign_in(5361) & VN_data_in(5361);
  VN893_in4 <= VN_sign_in(5362) & VN_data_in(5362);
  VN893_in5 <= VN_sign_in(5363) & VN_data_in(5363);
  VN894_in0 <= VN_sign_in(5364) & VN_data_in(5364);
  VN894_in1 <= VN_sign_in(5365) & VN_data_in(5365);
  VN894_in2 <= VN_sign_in(5366) & VN_data_in(5366);
  VN894_in3 <= VN_sign_in(5367) & VN_data_in(5367);
  VN894_in4 <= VN_sign_in(5368) & VN_data_in(5368);
  VN894_in5 <= VN_sign_in(5369) & VN_data_in(5369);
  VN895_in0 <= VN_sign_in(5370) & VN_data_in(5370);
  VN895_in1 <= VN_sign_in(5371) & VN_data_in(5371);
  VN895_in2 <= VN_sign_in(5372) & VN_data_in(5372);
  VN895_in3 <= VN_sign_in(5373) & VN_data_in(5373);
  VN895_in4 <= VN_sign_in(5374) & VN_data_in(5374);
  VN895_in5 <= VN_sign_in(5375) & VN_data_in(5375);
  VN896_in0 <= VN_sign_in(5376) & VN_data_in(5376);
  VN896_in1 <= VN_sign_in(5377) & VN_data_in(5377);
  VN896_in2 <= VN_sign_in(5378) & VN_data_in(5378);
  VN896_in3 <= VN_sign_in(5379) & VN_data_in(5379);
  VN896_in4 <= VN_sign_in(5380) & VN_data_in(5380);
  VN896_in5 <= VN_sign_in(5381) & VN_data_in(5381);
  VN897_in0 <= VN_sign_in(5382) & VN_data_in(5382);
  VN897_in1 <= VN_sign_in(5383) & VN_data_in(5383);
  VN897_in2 <= VN_sign_in(5384) & VN_data_in(5384);
  VN897_in3 <= VN_sign_in(5385) & VN_data_in(5385);
  VN897_in4 <= VN_sign_in(5386) & VN_data_in(5386);
  VN897_in5 <= VN_sign_in(5387) & VN_data_in(5387);
  VN898_in0 <= VN_sign_in(5388) & VN_data_in(5388);
  VN898_in1 <= VN_sign_in(5389) & VN_data_in(5389);
  VN898_in2 <= VN_sign_in(5390) & VN_data_in(5390);
  VN898_in3 <= VN_sign_in(5391) & VN_data_in(5391);
  VN898_in4 <= VN_sign_in(5392) & VN_data_in(5392);
  VN898_in5 <= VN_sign_in(5393) & VN_data_in(5393);
  VN899_in0 <= VN_sign_in(5394) & VN_data_in(5394);
  VN899_in1 <= VN_sign_in(5395) & VN_data_in(5395);
  VN899_in2 <= VN_sign_in(5396) & VN_data_in(5396);
  VN899_in3 <= VN_sign_in(5397) & VN_data_in(5397);
  VN899_in4 <= VN_sign_in(5398) & VN_data_in(5398);
  VN899_in5 <= VN_sign_in(5399) & VN_data_in(5399);
  VN900_in0 <= VN_sign_in(5400) & VN_data_in(5400);
  VN900_in1 <= VN_sign_in(5401) & VN_data_in(5401);
  VN900_in2 <= VN_sign_in(5402) & VN_data_in(5402);
  VN900_in3 <= VN_sign_in(5403) & VN_data_in(5403);
  VN900_in4 <= VN_sign_in(5404) & VN_data_in(5404);
  VN900_in5 <= VN_sign_in(5405) & VN_data_in(5405);
  VN901_in0 <= VN_sign_in(5406) & VN_data_in(5406);
  VN901_in1 <= VN_sign_in(5407) & VN_data_in(5407);
  VN901_in2 <= VN_sign_in(5408) & VN_data_in(5408);
  VN901_in3 <= VN_sign_in(5409) & VN_data_in(5409);
  VN901_in4 <= VN_sign_in(5410) & VN_data_in(5410);
  VN901_in5 <= VN_sign_in(5411) & VN_data_in(5411);
  VN902_in0 <= VN_sign_in(5412) & VN_data_in(5412);
  VN902_in1 <= VN_sign_in(5413) & VN_data_in(5413);
  VN902_in2 <= VN_sign_in(5414) & VN_data_in(5414);
  VN902_in3 <= VN_sign_in(5415) & VN_data_in(5415);
  VN902_in4 <= VN_sign_in(5416) & VN_data_in(5416);
  VN902_in5 <= VN_sign_in(5417) & VN_data_in(5417);
  VN903_in0 <= VN_sign_in(5418) & VN_data_in(5418);
  VN903_in1 <= VN_sign_in(5419) & VN_data_in(5419);
  VN903_in2 <= VN_sign_in(5420) & VN_data_in(5420);
  VN903_in3 <= VN_sign_in(5421) & VN_data_in(5421);
  VN903_in4 <= VN_sign_in(5422) & VN_data_in(5422);
  VN903_in5 <= VN_sign_in(5423) & VN_data_in(5423);
  VN904_in0 <= VN_sign_in(5424) & VN_data_in(5424);
  VN904_in1 <= VN_sign_in(5425) & VN_data_in(5425);
  VN904_in2 <= VN_sign_in(5426) & VN_data_in(5426);
  VN904_in3 <= VN_sign_in(5427) & VN_data_in(5427);
  VN904_in4 <= VN_sign_in(5428) & VN_data_in(5428);
  VN904_in5 <= VN_sign_in(5429) & VN_data_in(5429);
  VN905_in0 <= VN_sign_in(5430) & VN_data_in(5430);
  VN905_in1 <= VN_sign_in(5431) & VN_data_in(5431);
  VN905_in2 <= VN_sign_in(5432) & VN_data_in(5432);
  VN905_in3 <= VN_sign_in(5433) & VN_data_in(5433);
  VN905_in4 <= VN_sign_in(5434) & VN_data_in(5434);
  VN905_in5 <= VN_sign_in(5435) & VN_data_in(5435);
  VN906_in0 <= VN_sign_in(5436) & VN_data_in(5436);
  VN906_in1 <= VN_sign_in(5437) & VN_data_in(5437);
  VN906_in2 <= VN_sign_in(5438) & VN_data_in(5438);
  VN906_in3 <= VN_sign_in(5439) & VN_data_in(5439);
  VN906_in4 <= VN_sign_in(5440) & VN_data_in(5440);
  VN906_in5 <= VN_sign_in(5441) & VN_data_in(5441);
  VN907_in0 <= VN_sign_in(5442) & VN_data_in(5442);
  VN907_in1 <= VN_sign_in(5443) & VN_data_in(5443);
  VN907_in2 <= VN_sign_in(5444) & VN_data_in(5444);
  VN907_in3 <= VN_sign_in(5445) & VN_data_in(5445);
  VN907_in4 <= VN_sign_in(5446) & VN_data_in(5446);
  VN907_in5 <= VN_sign_in(5447) & VN_data_in(5447);
  VN908_in0 <= VN_sign_in(5448) & VN_data_in(5448);
  VN908_in1 <= VN_sign_in(5449) & VN_data_in(5449);
  VN908_in2 <= VN_sign_in(5450) & VN_data_in(5450);
  VN908_in3 <= VN_sign_in(5451) & VN_data_in(5451);
  VN908_in4 <= VN_sign_in(5452) & VN_data_in(5452);
  VN908_in5 <= VN_sign_in(5453) & VN_data_in(5453);
  VN909_in0 <= VN_sign_in(5454) & VN_data_in(5454);
  VN909_in1 <= VN_sign_in(5455) & VN_data_in(5455);
  VN909_in2 <= VN_sign_in(5456) & VN_data_in(5456);
  VN909_in3 <= VN_sign_in(5457) & VN_data_in(5457);
  VN909_in4 <= VN_sign_in(5458) & VN_data_in(5458);
  VN909_in5 <= VN_sign_in(5459) & VN_data_in(5459);
  VN910_in0 <= VN_sign_in(5460) & VN_data_in(5460);
  VN910_in1 <= VN_sign_in(5461) & VN_data_in(5461);
  VN910_in2 <= VN_sign_in(5462) & VN_data_in(5462);
  VN910_in3 <= VN_sign_in(5463) & VN_data_in(5463);
  VN910_in4 <= VN_sign_in(5464) & VN_data_in(5464);
  VN910_in5 <= VN_sign_in(5465) & VN_data_in(5465);
  VN911_in0 <= VN_sign_in(5466) & VN_data_in(5466);
  VN911_in1 <= VN_sign_in(5467) & VN_data_in(5467);
  VN911_in2 <= VN_sign_in(5468) & VN_data_in(5468);
  VN911_in3 <= VN_sign_in(5469) & VN_data_in(5469);
  VN911_in4 <= VN_sign_in(5470) & VN_data_in(5470);
  VN911_in5 <= VN_sign_in(5471) & VN_data_in(5471);
  VN912_in0 <= VN_sign_in(5472) & VN_data_in(5472);
  VN912_in1 <= VN_sign_in(5473) & VN_data_in(5473);
  VN912_in2 <= VN_sign_in(5474) & VN_data_in(5474);
  VN912_in3 <= VN_sign_in(5475) & VN_data_in(5475);
  VN912_in4 <= VN_sign_in(5476) & VN_data_in(5476);
  VN912_in5 <= VN_sign_in(5477) & VN_data_in(5477);
  VN913_in0 <= VN_sign_in(5478) & VN_data_in(5478);
  VN913_in1 <= VN_sign_in(5479) & VN_data_in(5479);
  VN913_in2 <= VN_sign_in(5480) & VN_data_in(5480);
  VN913_in3 <= VN_sign_in(5481) & VN_data_in(5481);
  VN913_in4 <= VN_sign_in(5482) & VN_data_in(5482);
  VN913_in5 <= VN_sign_in(5483) & VN_data_in(5483);
  VN914_in0 <= VN_sign_in(5484) & VN_data_in(5484);
  VN914_in1 <= VN_sign_in(5485) & VN_data_in(5485);
  VN914_in2 <= VN_sign_in(5486) & VN_data_in(5486);
  VN914_in3 <= VN_sign_in(5487) & VN_data_in(5487);
  VN914_in4 <= VN_sign_in(5488) & VN_data_in(5488);
  VN914_in5 <= VN_sign_in(5489) & VN_data_in(5489);
  VN915_in0 <= VN_sign_in(5490) & VN_data_in(5490);
  VN915_in1 <= VN_sign_in(5491) & VN_data_in(5491);
  VN915_in2 <= VN_sign_in(5492) & VN_data_in(5492);
  VN915_in3 <= VN_sign_in(5493) & VN_data_in(5493);
  VN915_in4 <= VN_sign_in(5494) & VN_data_in(5494);
  VN915_in5 <= VN_sign_in(5495) & VN_data_in(5495);
  VN916_in0 <= VN_sign_in(5496) & VN_data_in(5496);
  VN916_in1 <= VN_sign_in(5497) & VN_data_in(5497);
  VN916_in2 <= VN_sign_in(5498) & VN_data_in(5498);
  VN916_in3 <= VN_sign_in(5499) & VN_data_in(5499);
  VN916_in4 <= VN_sign_in(5500) & VN_data_in(5500);
  VN916_in5 <= VN_sign_in(5501) & VN_data_in(5501);
  VN917_in0 <= VN_sign_in(5502) & VN_data_in(5502);
  VN917_in1 <= VN_sign_in(5503) & VN_data_in(5503);
  VN917_in2 <= VN_sign_in(5504) & VN_data_in(5504);
  VN917_in3 <= VN_sign_in(5505) & VN_data_in(5505);
  VN917_in4 <= VN_sign_in(5506) & VN_data_in(5506);
  VN917_in5 <= VN_sign_in(5507) & VN_data_in(5507);
  VN918_in0 <= VN_sign_in(5508) & VN_data_in(5508);
  VN918_in1 <= VN_sign_in(5509) & VN_data_in(5509);
  VN918_in2 <= VN_sign_in(5510) & VN_data_in(5510);
  VN918_in3 <= VN_sign_in(5511) & VN_data_in(5511);
  VN918_in4 <= VN_sign_in(5512) & VN_data_in(5512);
  VN918_in5 <= VN_sign_in(5513) & VN_data_in(5513);
  VN919_in0 <= VN_sign_in(5514) & VN_data_in(5514);
  VN919_in1 <= VN_sign_in(5515) & VN_data_in(5515);
  VN919_in2 <= VN_sign_in(5516) & VN_data_in(5516);
  VN919_in3 <= VN_sign_in(5517) & VN_data_in(5517);
  VN919_in4 <= VN_sign_in(5518) & VN_data_in(5518);
  VN919_in5 <= VN_sign_in(5519) & VN_data_in(5519);
  VN920_in0 <= VN_sign_in(5520) & VN_data_in(5520);
  VN920_in1 <= VN_sign_in(5521) & VN_data_in(5521);
  VN920_in2 <= VN_sign_in(5522) & VN_data_in(5522);
  VN920_in3 <= VN_sign_in(5523) & VN_data_in(5523);
  VN920_in4 <= VN_sign_in(5524) & VN_data_in(5524);
  VN920_in5 <= VN_sign_in(5525) & VN_data_in(5525);
  VN921_in0 <= VN_sign_in(5526) & VN_data_in(5526);
  VN921_in1 <= VN_sign_in(5527) & VN_data_in(5527);
  VN921_in2 <= VN_sign_in(5528) & VN_data_in(5528);
  VN921_in3 <= VN_sign_in(5529) & VN_data_in(5529);
  VN921_in4 <= VN_sign_in(5530) & VN_data_in(5530);
  VN921_in5 <= VN_sign_in(5531) & VN_data_in(5531);
  VN922_in0 <= VN_sign_in(5532) & VN_data_in(5532);
  VN922_in1 <= VN_sign_in(5533) & VN_data_in(5533);
  VN922_in2 <= VN_sign_in(5534) & VN_data_in(5534);
  VN922_in3 <= VN_sign_in(5535) & VN_data_in(5535);
  VN922_in4 <= VN_sign_in(5536) & VN_data_in(5536);
  VN922_in5 <= VN_sign_in(5537) & VN_data_in(5537);
  VN923_in0 <= VN_sign_in(5538) & VN_data_in(5538);
  VN923_in1 <= VN_sign_in(5539) & VN_data_in(5539);
  VN923_in2 <= VN_sign_in(5540) & VN_data_in(5540);
  VN923_in3 <= VN_sign_in(5541) & VN_data_in(5541);
  VN923_in4 <= VN_sign_in(5542) & VN_data_in(5542);
  VN923_in5 <= VN_sign_in(5543) & VN_data_in(5543);
  VN924_in0 <= VN_sign_in(5544) & VN_data_in(5544);
  VN924_in1 <= VN_sign_in(5545) & VN_data_in(5545);
  VN924_in2 <= VN_sign_in(5546) & VN_data_in(5546);
  VN924_in3 <= VN_sign_in(5547) & VN_data_in(5547);
  VN924_in4 <= VN_sign_in(5548) & VN_data_in(5548);
  VN924_in5 <= VN_sign_in(5549) & VN_data_in(5549);
  VN925_in0 <= VN_sign_in(5550) & VN_data_in(5550);
  VN925_in1 <= VN_sign_in(5551) & VN_data_in(5551);
  VN925_in2 <= VN_sign_in(5552) & VN_data_in(5552);
  VN925_in3 <= VN_sign_in(5553) & VN_data_in(5553);
  VN925_in4 <= VN_sign_in(5554) & VN_data_in(5554);
  VN925_in5 <= VN_sign_in(5555) & VN_data_in(5555);
  VN926_in0 <= VN_sign_in(5556) & VN_data_in(5556);
  VN926_in1 <= VN_sign_in(5557) & VN_data_in(5557);
  VN926_in2 <= VN_sign_in(5558) & VN_data_in(5558);
  VN926_in3 <= VN_sign_in(5559) & VN_data_in(5559);
  VN926_in4 <= VN_sign_in(5560) & VN_data_in(5560);
  VN926_in5 <= VN_sign_in(5561) & VN_data_in(5561);
  VN927_in0 <= VN_sign_in(5562) & VN_data_in(5562);
  VN927_in1 <= VN_sign_in(5563) & VN_data_in(5563);
  VN927_in2 <= VN_sign_in(5564) & VN_data_in(5564);
  VN927_in3 <= VN_sign_in(5565) & VN_data_in(5565);
  VN927_in4 <= VN_sign_in(5566) & VN_data_in(5566);
  VN927_in5 <= VN_sign_in(5567) & VN_data_in(5567);
  VN928_in0 <= VN_sign_in(5568) & VN_data_in(5568);
  VN928_in1 <= VN_sign_in(5569) & VN_data_in(5569);
  VN928_in2 <= VN_sign_in(5570) & VN_data_in(5570);
  VN928_in3 <= VN_sign_in(5571) & VN_data_in(5571);
  VN928_in4 <= VN_sign_in(5572) & VN_data_in(5572);
  VN928_in5 <= VN_sign_in(5573) & VN_data_in(5573);
  VN929_in0 <= VN_sign_in(5574) & VN_data_in(5574);
  VN929_in1 <= VN_sign_in(5575) & VN_data_in(5575);
  VN929_in2 <= VN_sign_in(5576) & VN_data_in(5576);
  VN929_in3 <= VN_sign_in(5577) & VN_data_in(5577);
  VN929_in4 <= VN_sign_in(5578) & VN_data_in(5578);
  VN929_in5 <= VN_sign_in(5579) & VN_data_in(5579);
  VN930_in0 <= VN_sign_in(5580) & VN_data_in(5580);
  VN930_in1 <= VN_sign_in(5581) & VN_data_in(5581);
  VN930_in2 <= VN_sign_in(5582) & VN_data_in(5582);
  VN930_in3 <= VN_sign_in(5583) & VN_data_in(5583);
  VN930_in4 <= VN_sign_in(5584) & VN_data_in(5584);
  VN930_in5 <= VN_sign_in(5585) & VN_data_in(5585);
  VN931_in0 <= VN_sign_in(5586) & VN_data_in(5586);
  VN931_in1 <= VN_sign_in(5587) & VN_data_in(5587);
  VN931_in2 <= VN_sign_in(5588) & VN_data_in(5588);
  VN931_in3 <= VN_sign_in(5589) & VN_data_in(5589);
  VN931_in4 <= VN_sign_in(5590) & VN_data_in(5590);
  VN931_in5 <= VN_sign_in(5591) & VN_data_in(5591);
  VN932_in0 <= VN_sign_in(5592) & VN_data_in(5592);
  VN932_in1 <= VN_sign_in(5593) & VN_data_in(5593);
  VN932_in2 <= VN_sign_in(5594) & VN_data_in(5594);
  VN932_in3 <= VN_sign_in(5595) & VN_data_in(5595);
  VN932_in4 <= VN_sign_in(5596) & VN_data_in(5596);
  VN932_in5 <= VN_sign_in(5597) & VN_data_in(5597);
  VN933_in0 <= VN_sign_in(5598) & VN_data_in(5598);
  VN933_in1 <= VN_sign_in(5599) & VN_data_in(5599);
  VN933_in2 <= VN_sign_in(5600) & VN_data_in(5600);
  VN933_in3 <= VN_sign_in(5601) & VN_data_in(5601);
  VN933_in4 <= VN_sign_in(5602) & VN_data_in(5602);
  VN933_in5 <= VN_sign_in(5603) & VN_data_in(5603);
  VN934_in0 <= VN_sign_in(5604) & VN_data_in(5604);
  VN934_in1 <= VN_sign_in(5605) & VN_data_in(5605);
  VN934_in2 <= VN_sign_in(5606) & VN_data_in(5606);
  VN934_in3 <= VN_sign_in(5607) & VN_data_in(5607);
  VN934_in4 <= VN_sign_in(5608) & VN_data_in(5608);
  VN934_in5 <= VN_sign_in(5609) & VN_data_in(5609);
  VN935_in0 <= VN_sign_in(5610) & VN_data_in(5610);
  VN935_in1 <= VN_sign_in(5611) & VN_data_in(5611);
  VN935_in2 <= VN_sign_in(5612) & VN_data_in(5612);
  VN935_in3 <= VN_sign_in(5613) & VN_data_in(5613);
  VN935_in4 <= VN_sign_in(5614) & VN_data_in(5614);
  VN935_in5 <= VN_sign_in(5615) & VN_data_in(5615);
  VN936_in0 <= VN_sign_in(5616) & VN_data_in(5616);
  VN936_in1 <= VN_sign_in(5617) & VN_data_in(5617);
  VN936_in2 <= VN_sign_in(5618) & VN_data_in(5618);
  VN936_in3 <= VN_sign_in(5619) & VN_data_in(5619);
  VN936_in4 <= VN_sign_in(5620) & VN_data_in(5620);
  VN936_in5 <= VN_sign_in(5621) & VN_data_in(5621);
  VN937_in0 <= VN_sign_in(5622) & VN_data_in(5622);
  VN937_in1 <= VN_sign_in(5623) & VN_data_in(5623);
  VN937_in2 <= VN_sign_in(5624) & VN_data_in(5624);
  VN937_in3 <= VN_sign_in(5625) & VN_data_in(5625);
  VN937_in4 <= VN_sign_in(5626) & VN_data_in(5626);
  VN937_in5 <= VN_sign_in(5627) & VN_data_in(5627);
  VN938_in0 <= VN_sign_in(5628) & VN_data_in(5628);
  VN938_in1 <= VN_sign_in(5629) & VN_data_in(5629);
  VN938_in2 <= VN_sign_in(5630) & VN_data_in(5630);
  VN938_in3 <= VN_sign_in(5631) & VN_data_in(5631);
  VN938_in4 <= VN_sign_in(5632) & VN_data_in(5632);
  VN938_in5 <= VN_sign_in(5633) & VN_data_in(5633);
  VN939_in0 <= VN_sign_in(5634) & VN_data_in(5634);
  VN939_in1 <= VN_sign_in(5635) & VN_data_in(5635);
  VN939_in2 <= VN_sign_in(5636) & VN_data_in(5636);
  VN939_in3 <= VN_sign_in(5637) & VN_data_in(5637);
  VN939_in4 <= VN_sign_in(5638) & VN_data_in(5638);
  VN939_in5 <= VN_sign_in(5639) & VN_data_in(5639);
  VN940_in0 <= VN_sign_in(5640) & VN_data_in(5640);
  VN940_in1 <= VN_sign_in(5641) & VN_data_in(5641);
  VN940_in2 <= VN_sign_in(5642) & VN_data_in(5642);
  VN940_in3 <= VN_sign_in(5643) & VN_data_in(5643);
  VN940_in4 <= VN_sign_in(5644) & VN_data_in(5644);
  VN940_in5 <= VN_sign_in(5645) & VN_data_in(5645);
  VN941_in0 <= VN_sign_in(5646) & VN_data_in(5646);
  VN941_in1 <= VN_sign_in(5647) & VN_data_in(5647);
  VN941_in2 <= VN_sign_in(5648) & VN_data_in(5648);
  VN941_in3 <= VN_sign_in(5649) & VN_data_in(5649);
  VN941_in4 <= VN_sign_in(5650) & VN_data_in(5650);
  VN941_in5 <= VN_sign_in(5651) & VN_data_in(5651);
  VN942_in0 <= VN_sign_in(5652) & VN_data_in(5652);
  VN942_in1 <= VN_sign_in(5653) & VN_data_in(5653);
  VN942_in2 <= VN_sign_in(5654) & VN_data_in(5654);
  VN942_in3 <= VN_sign_in(5655) & VN_data_in(5655);
  VN942_in4 <= VN_sign_in(5656) & VN_data_in(5656);
  VN942_in5 <= VN_sign_in(5657) & VN_data_in(5657);
  VN943_in0 <= VN_sign_in(5658) & VN_data_in(5658);
  VN943_in1 <= VN_sign_in(5659) & VN_data_in(5659);
  VN943_in2 <= VN_sign_in(5660) & VN_data_in(5660);
  VN943_in3 <= VN_sign_in(5661) & VN_data_in(5661);
  VN943_in4 <= VN_sign_in(5662) & VN_data_in(5662);
  VN943_in5 <= VN_sign_in(5663) & VN_data_in(5663);
  VN944_in0 <= VN_sign_in(5664) & VN_data_in(5664);
  VN944_in1 <= VN_sign_in(5665) & VN_data_in(5665);
  VN944_in2 <= VN_sign_in(5666) & VN_data_in(5666);
  VN944_in3 <= VN_sign_in(5667) & VN_data_in(5667);
  VN944_in4 <= VN_sign_in(5668) & VN_data_in(5668);
  VN944_in5 <= VN_sign_in(5669) & VN_data_in(5669);
  VN945_in0 <= VN_sign_in(5670) & VN_data_in(5670);
  VN945_in1 <= VN_sign_in(5671) & VN_data_in(5671);
  VN945_in2 <= VN_sign_in(5672) & VN_data_in(5672);
  VN945_in3 <= VN_sign_in(5673) & VN_data_in(5673);
  VN945_in4 <= VN_sign_in(5674) & VN_data_in(5674);
  VN945_in5 <= VN_sign_in(5675) & VN_data_in(5675);
  VN946_in0 <= VN_sign_in(5676) & VN_data_in(5676);
  VN946_in1 <= VN_sign_in(5677) & VN_data_in(5677);
  VN946_in2 <= VN_sign_in(5678) & VN_data_in(5678);
  VN946_in3 <= VN_sign_in(5679) & VN_data_in(5679);
  VN946_in4 <= VN_sign_in(5680) & VN_data_in(5680);
  VN946_in5 <= VN_sign_in(5681) & VN_data_in(5681);
  VN947_in0 <= VN_sign_in(5682) & VN_data_in(5682);
  VN947_in1 <= VN_sign_in(5683) & VN_data_in(5683);
  VN947_in2 <= VN_sign_in(5684) & VN_data_in(5684);
  VN947_in3 <= VN_sign_in(5685) & VN_data_in(5685);
  VN947_in4 <= VN_sign_in(5686) & VN_data_in(5686);
  VN947_in5 <= VN_sign_in(5687) & VN_data_in(5687);
  VN948_in0 <= VN_sign_in(5688) & VN_data_in(5688);
  VN948_in1 <= VN_sign_in(5689) & VN_data_in(5689);
  VN948_in2 <= VN_sign_in(5690) & VN_data_in(5690);
  VN948_in3 <= VN_sign_in(5691) & VN_data_in(5691);
  VN948_in4 <= VN_sign_in(5692) & VN_data_in(5692);
  VN948_in5 <= VN_sign_in(5693) & VN_data_in(5693);
  VN949_in0 <= VN_sign_in(5694) & VN_data_in(5694);
  VN949_in1 <= VN_sign_in(5695) & VN_data_in(5695);
  VN949_in2 <= VN_sign_in(5696) & VN_data_in(5696);
  VN949_in3 <= VN_sign_in(5697) & VN_data_in(5697);
  VN949_in4 <= VN_sign_in(5698) & VN_data_in(5698);
  VN949_in5 <= VN_sign_in(5699) & VN_data_in(5699);
  VN950_in0 <= VN_sign_in(5700) & VN_data_in(5700);
  VN950_in1 <= VN_sign_in(5701) & VN_data_in(5701);
  VN950_in2 <= VN_sign_in(5702) & VN_data_in(5702);
  VN950_in3 <= VN_sign_in(5703) & VN_data_in(5703);
  VN950_in4 <= VN_sign_in(5704) & VN_data_in(5704);
  VN950_in5 <= VN_sign_in(5705) & VN_data_in(5705);
  VN951_in0 <= VN_sign_in(5706) & VN_data_in(5706);
  VN951_in1 <= VN_sign_in(5707) & VN_data_in(5707);
  VN951_in2 <= VN_sign_in(5708) & VN_data_in(5708);
  VN951_in3 <= VN_sign_in(5709) & VN_data_in(5709);
  VN951_in4 <= VN_sign_in(5710) & VN_data_in(5710);
  VN951_in5 <= VN_sign_in(5711) & VN_data_in(5711);
  VN952_in0 <= VN_sign_in(5712) & VN_data_in(5712);
  VN952_in1 <= VN_sign_in(5713) & VN_data_in(5713);
  VN952_in2 <= VN_sign_in(5714) & VN_data_in(5714);
  VN952_in3 <= VN_sign_in(5715) & VN_data_in(5715);
  VN952_in4 <= VN_sign_in(5716) & VN_data_in(5716);
  VN952_in5 <= VN_sign_in(5717) & VN_data_in(5717);
  VN953_in0 <= VN_sign_in(5718) & VN_data_in(5718);
  VN953_in1 <= VN_sign_in(5719) & VN_data_in(5719);
  VN953_in2 <= VN_sign_in(5720) & VN_data_in(5720);
  VN953_in3 <= VN_sign_in(5721) & VN_data_in(5721);
  VN953_in4 <= VN_sign_in(5722) & VN_data_in(5722);
  VN953_in5 <= VN_sign_in(5723) & VN_data_in(5723);
  VN954_in0 <= VN_sign_in(5724) & VN_data_in(5724);
  VN954_in1 <= VN_sign_in(5725) & VN_data_in(5725);
  VN954_in2 <= VN_sign_in(5726) & VN_data_in(5726);
  VN954_in3 <= VN_sign_in(5727) & VN_data_in(5727);
  VN954_in4 <= VN_sign_in(5728) & VN_data_in(5728);
  VN954_in5 <= VN_sign_in(5729) & VN_data_in(5729);
  VN955_in0 <= VN_sign_in(5730) & VN_data_in(5730);
  VN955_in1 <= VN_sign_in(5731) & VN_data_in(5731);
  VN955_in2 <= VN_sign_in(5732) & VN_data_in(5732);
  VN955_in3 <= VN_sign_in(5733) & VN_data_in(5733);
  VN955_in4 <= VN_sign_in(5734) & VN_data_in(5734);
  VN955_in5 <= VN_sign_in(5735) & VN_data_in(5735);
  VN956_in0 <= VN_sign_in(5736) & VN_data_in(5736);
  VN956_in1 <= VN_sign_in(5737) & VN_data_in(5737);
  VN956_in2 <= VN_sign_in(5738) & VN_data_in(5738);
  VN956_in3 <= VN_sign_in(5739) & VN_data_in(5739);
  VN956_in4 <= VN_sign_in(5740) & VN_data_in(5740);
  VN956_in5 <= VN_sign_in(5741) & VN_data_in(5741);
  VN957_in0 <= VN_sign_in(5742) & VN_data_in(5742);
  VN957_in1 <= VN_sign_in(5743) & VN_data_in(5743);
  VN957_in2 <= VN_sign_in(5744) & VN_data_in(5744);
  VN957_in3 <= VN_sign_in(5745) & VN_data_in(5745);
  VN957_in4 <= VN_sign_in(5746) & VN_data_in(5746);
  VN957_in5 <= VN_sign_in(5747) & VN_data_in(5747);
  VN958_in0 <= VN_sign_in(5748) & VN_data_in(5748);
  VN958_in1 <= VN_sign_in(5749) & VN_data_in(5749);
  VN958_in2 <= VN_sign_in(5750) & VN_data_in(5750);
  VN958_in3 <= VN_sign_in(5751) & VN_data_in(5751);
  VN958_in4 <= VN_sign_in(5752) & VN_data_in(5752);
  VN958_in5 <= VN_sign_in(5753) & VN_data_in(5753);
  VN959_in0 <= VN_sign_in(5754) & VN_data_in(5754);
  VN959_in1 <= VN_sign_in(5755) & VN_data_in(5755);
  VN959_in2 <= VN_sign_in(5756) & VN_data_in(5756);
  VN959_in3 <= VN_sign_in(5757) & VN_data_in(5757);
  VN959_in4 <= VN_sign_in(5758) & VN_data_in(5758);
  VN959_in5 <= VN_sign_in(5759) & VN_data_in(5759);
  VN960_in0 <= VN_sign_in(5760) & VN_data_in(5760);
  VN960_in1 <= VN_sign_in(5761) & VN_data_in(5761);
  VN960_in2 <= VN_sign_in(5762) & VN_data_in(5762);
  VN960_in3 <= VN_sign_in(5763) & VN_data_in(5763);
  VN960_in4 <= VN_sign_in(5764) & VN_data_in(5764);
  VN960_in5 <= VN_sign_in(5765) & VN_data_in(5765);
  VN961_in0 <= VN_sign_in(5766) & VN_data_in(5766);
  VN961_in1 <= VN_sign_in(5767) & VN_data_in(5767);
  VN961_in2 <= VN_sign_in(5768) & VN_data_in(5768);
  VN961_in3 <= VN_sign_in(5769) & VN_data_in(5769);
  VN961_in4 <= VN_sign_in(5770) & VN_data_in(5770);
  VN961_in5 <= VN_sign_in(5771) & VN_data_in(5771);
  VN962_in0 <= VN_sign_in(5772) & VN_data_in(5772);
  VN962_in1 <= VN_sign_in(5773) & VN_data_in(5773);
  VN962_in2 <= VN_sign_in(5774) & VN_data_in(5774);
  VN962_in3 <= VN_sign_in(5775) & VN_data_in(5775);
  VN962_in4 <= VN_sign_in(5776) & VN_data_in(5776);
  VN962_in5 <= VN_sign_in(5777) & VN_data_in(5777);
  VN963_in0 <= VN_sign_in(5778) & VN_data_in(5778);
  VN963_in1 <= VN_sign_in(5779) & VN_data_in(5779);
  VN963_in2 <= VN_sign_in(5780) & VN_data_in(5780);
  VN963_in3 <= VN_sign_in(5781) & VN_data_in(5781);
  VN963_in4 <= VN_sign_in(5782) & VN_data_in(5782);
  VN963_in5 <= VN_sign_in(5783) & VN_data_in(5783);
  VN964_in0 <= VN_sign_in(5784) & VN_data_in(5784);
  VN964_in1 <= VN_sign_in(5785) & VN_data_in(5785);
  VN964_in2 <= VN_sign_in(5786) & VN_data_in(5786);
  VN964_in3 <= VN_sign_in(5787) & VN_data_in(5787);
  VN964_in4 <= VN_sign_in(5788) & VN_data_in(5788);
  VN964_in5 <= VN_sign_in(5789) & VN_data_in(5789);
  VN965_in0 <= VN_sign_in(5790) & VN_data_in(5790);
  VN965_in1 <= VN_sign_in(5791) & VN_data_in(5791);
  VN965_in2 <= VN_sign_in(5792) & VN_data_in(5792);
  VN965_in3 <= VN_sign_in(5793) & VN_data_in(5793);
  VN965_in4 <= VN_sign_in(5794) & VN_data_in(5794);
  VN965_in5 <= VN_sign_in(5795) & VN_data_in(5795);
  VN966_in0 <= VN_sign_in(5796) & VN_data_in(5796);
  VN966_in1 <= VN_sign_in(5797) & VN_data_in(5797);
  VN966_in2 <= VN_sign_in(5798) & VN_data_in(5798);
  VN966_in3 <= VN_sign_in(5799) & VN_data_in(5799);
  VN966_in4 <= VN_sign_in(5800) & VN_data_in(5800);
  VN966_in5 <= VN_sign_in(5801) & VN_data_in(5801);
  VN967_in0 <= VN_sign_in(5802) & VN_data_in(5802);
  VN967_in1 <= VN_sign_in(5803) & VN_data_in(5803);
  VN967_in2 <= VN_sign_in(5804) & VN_data_in(5804);
  VN967_in3 <= VN_sign_in(5805) & VN_data_in(5805);
  VN967_in4 <= VN_sign_in(5806) & VN_data_in(5806);
  VN967_in5 <= VN_sign_in(5807) & VN_data_in(5807);
  VN968_in0 <= VN_sign_in(5808) & VN_data_in(5808);
  VN968_in1 <= VN_sign_in(5809) & VN_data_in(5809);
  VN968_in2 <= VN_sign_in(5810) & VN_data_in(5810);
  VN968_in3 <= VN_sign_in(5811) & VN_data_in(5811);
  VN968_in4 <= VN_sign_in(5812) & VN_data_in(5812);
  VN968_in5 <= VN_sign_in(5813) & VN_data_in(5813);
  VN969_in0 <= VN_sign_in(5814) & VN_data_in(5814);
  VN969_in1 <= VN_sign_in(5815) & VN_data_in(5815);
  VN969_in2 <= VN_sign_in(5816) & VN_data_in(5816);
  VN969_in3 <= VN_sign_in(5817) & VN_data_in(5817);
  VN969_in4 <= VN_sign_in(5818) & VN_data_in(5818);
  VN969_in5 <= VN_sign_in(5819) & VN_data_in(5819);
  VN970_in0 <= VN_sign_in(5820) & VN_data_in(5820);
  VN970_in1 <= VN_sign_in(5821) & VN_data_in(5821);
  VN970_in2 <= VN_sign_in(5822) & VN_data_in(5822);
  VN970_in3 <= VN_sign_in(5823) & VN_data_in(5823);
  VN970_in4 <= VN_sign_in(5824) & VN_data_in(5824);
  VN970_in5 <= VN_sign_in(5825) & VN_data_in(5825);
  VN971_in0 <= VN_sign_in(5826) & VN_data_in(5826);
  VN971_in1 <= VN_sign_in(5827) & VN_data_in(5827);
  VN971_in2 <= VN_sign_in(5828) & VN_data_in(5828);
  VN971_in3 <= VN_sign_in(5829) & VN_data_in(5829);
  VN971_in4 <= VN_sign_in(5830) & VN_data_in(5830);
  VN971_in5 <= VN_sign_in(5831) & VN_data_in(5831);
  VN972_in0 <= VN_sign_in(5832) & VN_data_in(5832);
  VN972_in1 <= VN_sign_in(5833) & VN_data_in(5833);
  VN972_in2 <= VN_sign_in(5834) & VN_data_in(5834);
  VN972_in3 <= VN_sign_in(5835) & VN_data_in(5835);
  VN972_in4 <= VN_sign_in(5836) & VN_data_in(5836);
  VN972_in5 <= VN_sign_in(5837) & VN_data_in(5837);
  VN973_in0 <= VN_sign_in(5838) & VN_data_in(5838);
  VN973_in1 <= VN_sign_in(5839) & VN_data_in(5839);
  VN973_in2 <= VN_sign_in(5840) & VN_data_in(5840);
  VN973_in3 <= VN_sign_in(5841) & VN_data_in(5841);
  VN973_in4 <= VN_sign_in(5842) & VN_data_in(5842);
  VN973_in5 <= VN_sign_in(5843) & VN_data_in(5843);
  VN974_in0 <= VN_sign_in(5844) & VN_data_in(5844);
  VN974_in1 <= VN_sign_in(5845) & VN_data_in(5845);
  VN974_in2 <= VN_sign_in(5846) & VN_data_in(5846);
  VN974_in3 <= VN_sign_in(5847) & VN_data_in(5847);
  VN974_in4 <= VN_sign_in(5848) & VN_data_in(5848);
  VN974_in5 <= VN_sign_in(5849) & VN_data_in(5849);
  VN975_in0 <= VN_sign_in(5850) & VN_data_in(5850);
  VN975_in1 <= VN_sign_in(5851) & VN_data_in(5851);
  VN975_in2 <= VN_sign_in(5852) & VN_data_in(5852);
  VN975_in3 <= VN_sign_in(5853) & VN_data_in(5853);
  VN975_in4 <= VN_sign_in(5854) & VN_data_in(5854);
  VN975_in5 <= VN_sign_in(5855) & VN_data_in(5855);
  VN976_in0 <= VN_sign_in(5856) & VN_data_in(5856);
  VN976_in1 <= VN_sign_in(5857) & VN_data_in(5857);
  VN976_in2 <= VN_sign_in(5858) & VN_data_in(5858);
  VN976_in3 <= VN_sign_in(5859) & VN_data_in(5859);
  VN976_in4 <= VN_sign_in(5860) & VN_data_in(5860);
  VN976_in5 <= VN_sign_in(5861) & VN_data_in(5861);
  VN977_in0 <= VN_sign_in(5862) & VN_data_in(5862);
  VN977_in1 <= VN_sign_in(5863) & VN_data_in(5863);
  VN977_in2 <= VN_sign_in(5864) & VN_data_in(5864);
  VN977_in3 <= VN_sign_in(5865) & VN_data_in(5865);
  VN977_in4 <= VN_sign_in(5866) & VN_data_in(5866);
  VN977_in5 <= VN_sign_in(5867) & VN_data_in(5867);
  VN978_in0 <= VN_sign_in(5868) & VN_data_in(5868);
  VN978_in1 <= VN_sign_in(5869) & VN_data_in(5869);
  VN978_in2 <= VN_sign_in(5870) & VN_data_in(5870);
  VN978_in3 <= VN_sign_in(5871) & VN_data_in(5871);
  VN978_in4 <= VN_sign_in(5872) & VN_data_in(5872);
  VN978_in5 <= VN_sign_in(5873) & VN_data_in(5873);
  VN979_in0 <= VN_sign_in(5874) & VN_data_in(5874);
  VN979_in1 <= VN_sign_in(5875) & VN_data_in(5875);
  VN979_in2 <= VN_sign_in(5876) & VN_data_in(5876);
  VN979_in3 <= VN_sign_in(5877) & VN_data_in(5877);
  VN979_in4 <= VN_sign_in(5878) & VN_data_in(5878);
  VN979_in5 <= VN_sign_in(5879) & VN_data_in(5879);
  VN980_in0 <= VN_sign_in(5880) & VN_data_in(5880);
  VN980_in1 <= VN_sign_in(5881) & VN_data_in(5881);
  VN980_in2 <= VN_sign_in(5882) & VN_data_in(5882);
  VN980_in3 <= VN_sign_in(5883) & VN_data_in(5883);
  VN980_in4 <= VN_sign_in(5884) & VN_data_in(5884);
  VN980_in5 <= VN_sign_in(5885) & VN_data_in(5885);
  VN981_in0 <= VN_sign_in(5886) & VN_data_in(5886);
  VN981_in1 <= VN_sign_in(5887) & VN_data_in(5887);
  VN981_in2 <= VN_sign_in(5888) & VN_data_in(5888);
  VN981_in3 <= VN_sign_in(5889) & VN_data_in(5889);
  VN981_in4 <= VN_sign_in(5890) & VN_data_in(5890);
  VN981_in5 <= VN_sign_in(5891) & VN_data_in(5891);
  VN982_in0 <= VN_sign_in(5892) & VN_data_in(5892);
  VN982_in1 <= VN_sign_in(5893) & VN_data_in(5893);
  VN982_in2 <= VN_sign_in(5894) & VN_data_in(5894);
  VN982_in3 <= VN_sign_in(5895) & VN_data_in(5895);
  VN982_in4 <= VN_sign_in(5896) & VN_data_in(5896);
  VN982_in5 <= VN_sign_in(5897) & VN_data_in(5897);
  VN983_in0 <= VN_sign_in(5898) & VN_data_in(5898);
  VN983_in1 <= VN_sign_in(5899) & VN_data_in(5899);
  VN983_in2 <= VN_sign_in(5900) & VN_data_in(5900);
  VN983_in3 <= VN_sign_in(5901) & VN_data_in(5901);
  VN983_in4 <= VN_sign_in(5902) & VN_data_in(5902);
  VN983_in5 <= VN_sign_in(5903) & VN_data_in(5903);
  VN984_in0 <= VN_sign_in(5904) & VN_data_in(5904);
  VN984_in1 <= VN_sign_in(5905) & VN_data_in(5905);
  VN984_in2 <= VN_sign_in(5906) & VN_data_in(5906);
  VN984_in3 <= VN_sign_in(5907) & VN_data_in(5907);
  VN984_in4 <= VN_sign_in(5908) & VN_data_in(5908);
  VN984_in5 <= VN_sign_in(5909) & VN_data_in(5909);
  VN985_in0 <= VN_sign_in(5910) & VN_data_in(5910);
  VN985_in1 <= VN_sign_in(5911) & VN_data_in(5911);
  VN985_in2 <= VN_sign_in(5912) & VN_data_in(5912);
  VN985_in3 <= VN_sign_in(5913) & VN_data_in(5913);
  VN985_in4 <= VN_sign_in(5914) & VN_data_in(5914);
  VN985_in5 <= VN_sign_in(5915) & VN_data_in(5915);
  VN986_in0 <= VN_sign_in(5916) & VN_data_in(5916);
  VN986_in1 <= VN_sign_in(5917) & VN_data_in(5917);
  VN986_in2 <= VN_sign_in(5918) & VN_data_in(5918);
  VN986_in3 <= VN_sign_in(5919) & VN_data_in(5919);
  VN986_in4 <= VN_sign_in(5920) & VN_data_in(5920);
  VN986_in5 <= VN_sign_in(5921) & VN_data_in(5921);
  VN987_in0 <= VN_sign_in(5922) & VN_data_in(5922);
  VN987_in1 <= VN_sign_in(5923) & VN_data_in(5923);
  VN987_in2 <= VN_sign_in(5924) & VN_data_in(5924);
  VN987_in3 <= VN_sign_in(5925) & VN_data_in(5925);
  VN987_in4 <= VN_sign_in(5926) & VN_data_in(5926);
  VN987_in5 <= VN_sign_in(5927) & VN_data_in(5927);
  VN988_in0 <= VN_sign_in(5928) & VN_data_in(5928);
  VN988_in1 <= VN_sign_in(5929) & VN_data_in(5929);
  VN988_in2 <= VN_sign_in(5930) & VN_data_in(5930);
  VN988_in3 <= VN_sign_in(5931) & VN_data_in(5931);
  VN988_in4 <= VN_sign_in(5932) & VN_data_in(5932);
  VN988_in5 <= VN_sign_in(5933) & VN_data_in(5933);
  VN989_in0 <= VN_sign_in(5934) & VN_data_in(5934);
  VN989_in1 <= VN_sign_in(5935) & VN_data_in(5935);
  VN989_in2 <= VN_sign_in(5936) & VN_data_in(5936);
  VN989_in3 <= VN_sign_in(5937) & VN_data_in(5937);
  VN989_in4 <= VN_sign_in(5938) & VN_data_in(5938);
  VN989_in5 <= VN_sign_in(5939) & VN_data_in(5939);
  VN990_in0 <= VN_sign_in(5940) & VN_data_in(5940);
  VN990_in1 <= VN_sign_in(5941) & VN_data_in(5941);
  VN990_in2 <= VN_sign_in(5942) & VN_data_in(5942);
  VN990_in3 <= VN_sign_in(5943) & VN_data_in(5943);
  VN990_in4 <= VN_sign_in(5944) & VN_data_in(5944);
  VN990_in5 <= VN_sign_in(5945) & VN_data_in(5945);
  VN991_in0 <= VN_sign_in(5946) & VN_data_in(5946);
  VN991_in1 <= VN_sign_in(5947) & VN_data_in(5947);
  VN991_in2 <= VN_sign_in(5948) & VN_data_in(5948);
  VN991_in3 <= VN_sign_in(5949) & VN_data_in(5949);
  VN991_in4 <= VN_sign_in(5950) & VN_data_in(5950);
  VN991_in5 <= VN_sign_in(5951) & VN_data_in(5951);
  VN992_in0 <= VN_sign_in(5952) & VN_data_in(5952);
  VN992_in1 <= VN_sign_in(5953) & VN_data_in(5953);
  VN992_in2 <= VN_sign_in(5954) & VN_data_in(5954);
  VN992_in3 <= VN_sign_in(5955) & VN_data_in(5955);
  VN992_in4 <= VN_sign_in(5956) & VN_data_in(5956);
  VN992_in5 <= VN_sign_in(5957) & VN_data_in(5957);
  VN993_in0 <= VN_sign_in(5958) & VN_data_in(5958);
  VN993_in1 <= VN_sign_in(5959) & VN_data_in(5959);
  VN993_in2 <= VN_sign_in(5960) & VN_data_in(5960);
  VN993_in3 <= VN_sign_in(5961) & VN_data_in(5961);
  VN993_in4 <= VN_sign_in(5962) & VN_data_in(5962);
  VN993_in5 <= VN_sign_in(5963) & VN_data_in(5963);
  VN994_in0 <= VN_sign_in(5964) & VN_data_in(5964);
  VN994_in1 <= VN_sign_in(5965) & VN_data_in(5965);
  VN994_in2 <= VN_sign_in(5966) & VN_data_in(5966);
  VN994_in3 <= VN_sign_in(5967) & VN_data_in(5967);
  VN994_in4 <= VN_sign_in(5968) & VN_data_in(5968);
  VN994_in5 <= VN_sign_in(5969) & VN_data_in(5969);
  VN995_in0 <= VN_sign_in(5970) & VN_data_in(5970);
  VN995_in1 <= VN_sign_in(5971) & VN_data_in(5971);
  VN995_in2 <= VN_sign_in(5972) & VN_data_in(5972);
  VN995_in3 <= VN_sign_in(5973) & VN_data_in(5973);
  VN995_in4 <= VN_sign_in(5974) & VN_data_in(5974);
  VN995_in5 <= VN_sign_in(5975) & VN_data_in(5975);
  VN996_in0 <= VN_sign_in(5976) & VN_data_in(5976);
  VN996_in1 <= VN_sign_in(5977) & VN_data_in(5977);
  VN996_in2 <= VN_sign_in(5978) & VN_data_in(5978);
  VN996_in3 <= VN_sign_in(5979) & VN_data_in(5979);
  VN996_in4 <= VN_sign_in(5980) & VN_data_in(5980);
  VN996_in5 <= VN_sign_in(5981) & VN_data_in(5981);
  VN997_in0 <= VN_sign_in(5982) & VN_data_in(5982);
  VN997_in1 <= VN_sign_in(5983) & VN_data_in(5983);
  VN997_in2 <= VN_sign_in(5984) & VN_data_in(5984);
  VN997_in3 <= VN_sign_in(5985) & VN_data_in(5985);
  VN997_in4 <= VN_sign_in(5986) & VN_data_in(5986);
  VN997_in5 <= VN_sign_in(5987) & VN_data_in(5987);
  VN998_in0 <= VN_sign_in(5988) & VN_data_in(5988);
  VN998_in1 <= VN_sign_in(5989) & VN_data_in(5989);
  VN998_in2 <= VN_sign_in(5990) & VN_data_in(5990);
  VN998_in3 <= VN_sign_in(5991) & VN_data_in(5991);
  VN998_in4 <= VN_sign_in(5992) & VN_data_in(5992);
  VN998_in5 <= VN_sign_in(5993) & VN_data_in(5993);
  VN999_in0 <= VN_sign_in(5994) & VN_data_in(5994);
  VN999_in1 <= VN_sign_in(5995) & VN_data_in(5995);
  VN999_in2 <= VN_sign_in(5996) & VN_data_in(5996);
  VN999_in3 <= VN_sign_in(5997) & VN_data_in(5997);
  VN999_in4 <= VN_sign_in(5998) & VN_data_in(5998);
  VN999_in5 <= VN_sign_in(5999) & VN_data_in(5999);
  VN1000_in0 <= VN_sign_in(6000) & VN_data_in(6000);
  VN1000_in1 <= VN_sign_in(6001) & VN_data_in(6001);
  VN1000_in2 <= VN_sign_in(6002) & VN_data_in(6002);
  VN1000_in3 <= VN_sign_in(6003) & VN_data_in(6003);
  VN1000_in4 <= VN_sign_in(6004) & VN_data_in(6004);
  VN1000_in5 <= VN_sign_in(6005) & VN_data_in(6005);
  VN1001_in0 <= VN_sign_in(6006) & VN_data_in(6006);
  VN1001_in1 <= VN_sign_in(6007) & VN_data_in(6007);
  VN1001_in2 <= VN_sign_in(6008) & VN_data_in(6008);
  VN1001_in3 <= VN_sign_in(6009) & VN_data_in(6009);
  VN1001_in4 <= VN_sign_in(6010) & VN_data_in(6010);
  VN1001_in5 <= VN_sign_in(6011) & VN_data_in(6011);
  VN1002_in0 <= VN_sign_in(6012) & VN_data_in(6012);
  VN1002_in1 <= VN_sign_in(6013) & VN_data_in(6013);
  VN1002_in2 <= VN_sign_in(6014) & VN_data_in(6014);
  VN1002_in3 <= VN_sign_in(6015) & VN_data_in(6015);
  VN1002_in4 <= VN_sign_in(6016) & VN_data_in(6016);
  VN1002_in5 <= VN_sign_in(6017) & VN_data_in(6017);
  VN1003_in0 <= VN_sign_in(6018) & VN_data_in(6018);
  VN1003_in1 <= VN_sign_in(6019) & VN_data_in(6019);
  VN1003_in2 <= VN_sign_in(6020) & VN_data_in(6020);
  VN1003_in3 <= VN_sign_in(6021) & VN_data_in(6021);
  VN1003_in4 <= VN_sign_in(6022) & VN_data_in(6022);
  VN1003_in5 <= VN_sign_in(6023) & VN_data_in(6023);
  VN1004_in0 <= VN_sign_in(6024) & VN_data_in(6024);
  VN1004_in1 <= VN_sign_in(6025) & VN_data_in(6025);
  VN1004_in2 <= VN_sign_in(6026) & VN_data_in(6026);
  VN1004_in3 <= VN_sign_in(6027) & VN_data_in(6027);
  VN1004_in4 <= VN_sign_in(6028) & VN_data_in(6028);
  VN1004_in5 <= VN_sign_in(6029) & VN_data_in(6029);
  VN1005_in0 <= VN_sign_in(6030) & VN_data_in(6030);
  VN1005_in1 <= VN_sign_in(6031) & VN_data_in(6031);
  VN1005_in2 <= VN_sign_in(6032) & VN_data_in(6032);
  VN1005_in3 <= VN_sign_in(6033) & VN_data_in(6033);
  VN1005_in4 <= VN_sign_in(6034) & VN_data_in(6034);
  VN1005_in5 <= VN_sign_in(6035) & VN_data_in(6035);
  VN1006_in0 <= VN_sign_in(6036) & VN_data_in(6036);
  VN1006_in1 <= VN_sign_in(6037) & VN_data_in(6037);
  VN1006_in2 <= VN_sign_in(6038) & VN_data_in(6038);
  VN1006_in3 <= VN_sign_in(6039) & VN_data_in(6039);
  VN1006_in4 <= VN_sign_in(6040) & VN_data_in(6040);
  VN1006_in5 <= VN_sign_in(6041) & VN_data_in(6041);
  VN1007_in0 <= VN_sign_in(6042) & VN_data_in(6042);
  VN1007_in1 <= VN_sign_in(6043) & VN_data_in(6043);
  VN1007_in2 <= VN_sign_in(6044) & VN_data_in(6044);
  VN1007_in3 <= VN_sign_in(6045) & VN_data_in(6045);
  VN1007_in4 <= VN_sign_in(6046) & VN_data_in(6046);
  VN1007_in5 <= VN_sign_in(6047) & VN_data_in(6047);
  VN1008_in0 <= VN_sign_in(6048) & VN_data_in(6048);
  VN1008_in1 <= VN_sign_in(6049) & VN_data_in(6049);
  VN1008_in2 <= VN_sign_in(6050) & VN_data_in(6050);
  VN1008_in3 <= VN_sign_in(6051) & VN_data_in(6051);
  VN1008_in4 <= VN_sign_in(6052) & VN_data_in(6052);
  VN1008_in5 <= VN_sign_in(6053) & VN_data_in(6053);
  VN1009_in0 <= VN_sign_in(6054) & VN_data_in(6054);
  VN1009_in1 <= VN_sign_in(6055) & VN_data_in(6055);
  VN1009_in2 <= VN_sign_in(6056) & VN_data_in(6056);
  VN1009_in3 <= VN_sign_in(6057) & VN_data_in(6057);
  VN1009_in4 <= VN_sign_in(6058) & VN_data_in(6058);
  VN1009_in5 <= VN_sign_in(6059) & VN_data_in(6059);
  VN1010_in0 <= VN_sign_in(6060) & VN_data_in(6060);
  VN1010_in1 <= VN_sign_in(6061) & VN_data_in(6061);
  VN1010_in2 <= VN_sign_in(6062) & VN_data_in(6062);
  VN1010_in3 <= VN_sign_in(6063) & VN_data_in(6063);
  VN1010_in4 <= VN_sign_in(6064) & VN_data_in(6064);
  VN1010_in5 <= VN_sign_in(6065) & VN_data_in(6065);
  VN1011_in0 <= VN_sign_in(6066) & VN_data_in(6066);
  VN1011_in1 <= VN_sign_in(6067) & VN_data_in(6067);
  VN1011_in2 <= VN_sign_in(6068) & VN_data_in(6068);
  VN1011_in3 <= VN_sign_in(6069) & VN_data_in(6069);
  VN1011_in4 <= VN_sign_in(6070) & VN_data_in(6070);
  VN1011_in5 <= VN_sign_in(6071) & VN_data_in(6071);
  VN1012_in0 <= VN_sign_in(6072) & VN_data_in(6072);
  VN1012_in1 <= VN_sign_in(6073) & VN_data_in(6073);
  VN1012_in2 <= VN_sign_in(6074) & VN_data_in(6074);
  VN1012_in3 <= VN_sign_in(6075) & VN_data_in(6075);
  VN1012_in4 <= VN_sign_in(6076) & VN_data_in(6076);
  VN1012_in5 <= VN_sign_in(6077) & VN_data_in(6077);
  VN1013_in0 <= VN_sign_in(6078) & VN_data_in(6078);
  VN1013_in1 <= VN_sign_in(6079) & VN_data_in(6079);
  VN1013_in2 <= VN_sign_in(6080) & VN_data_in(6080);
  VN1013_in3 <= VN_sign_in(6081) & VN_data_in(6081);
  VN1013_in4 <= VN_sign_in(6082) & VN_data_in(6082);
  VN1013_in5 <= VN_sign_in(6083) & VN_data_in(6083);
  VN1014_in0 <= VN_sign_in(6084) & VN_data_in(6084);
  VN1014_in1 <= VN_sign_in(6085) & VN_data_in(6085);
  VN1014_in2 <= VN_sign_in(6086) & VN_data_in(6086);
  VN1014_in3 <= VN_sign_in(6087) & VN_data_in(6087);
  VN1014_in4 <= VN_sign_in(6088) & VN_data_in(6088);
  VN1014_in5 <= VN_sign_in(6089) & VN_data_in(6089);
  VN1015_in0 <= VN_sign_in(6090) & VN_data_in(6090);
  VN1015_in1 <= VN_sign_in(6091) & VN_data_in(6091);
  VN1015_in2 <= VN_sign_in(6092) & VN_data_in(6092);
  VN1015_in3 <= VN_sign_in(6093) & VN_data_in(6093);
  VN1015_in4 <= VN_sign_in(6094) & VN_data_in(6094);
  VN1015_in5 <= VN_sign_in(6095) & VN_data_in(6095);
  VN1016_in0 <= VN_sign_in(6096) & VN_data_in(6096);
  VN1016_in1 <= VN_sign_in(6097) & VN_data_in(6097);
  VN1016_in2 <= VN_sign_in(6098) & VN_data_in(6098);
  VN1016_in3 <= VN_sign_in(6099) & VN_data_in(6099);
  VN1016_in4 <= VN_sign_in(6100) & VN_data_in(6100);
  VN1016_in5 <= VN_sign_in(6101) & VN_data_in(6101);
  VN1017_in0 <= VN_sign_in(6102) & VN_data_in(6102);
  VN1017_in1 <= VN_sign_in(6103) & VN_data_in(6103);
  VN1017_in2 <= VN_sign_in(6104) & VN_data_in(6104);
  VN1017_in3 <= VN_sign_in(6105) & VN_data_in(6105);
  VN1017_in4 <= VN_sign_in(6106) & VN_data_in(6106);
  VN1017_in5 <= VN_sign_in(6107) & VN_data_in(6107);
  VN1018_in0 <= VN_sign_in(6108) & VN_data_in(6108);
  VN1018_in1 <= VN_sign_in(6109) & VN_data_in(6109);
  VN1018_in2 <= VN_sign_in(6110) & VN_data_in(6110);
  VN1018_in3 <= VN_sign_in(6111) & VN_data_in(6111);
  VN1018_in4 <= VN_sign_in(6112) & VN_data_in(6112);
  VN1018_in5 <= VN_sign_in(6113) & VN_data_in(6113);
  VN1019_in0 <= VN_sign_in(6114) & VN_data_in(6114);
  VN1019_in1 <= VN_sign_in(6115) & VN_data_in(6115);
  VN1019_in2 <= VN_sign_in(6116) & VN_data_in(6116);
  VN1019_in3 <= VN_sign_in(6117) & VN_data_in(6117);
  VN1019_in4 <= VN_sign_in(6118) & VN_data_in(6118);
  VN1019_in5 <= VN_sign_in(6119) & VN_data_in(6119);
  VN1020_in0 <= VN_sign_in(6120) & VN_data_in(6120);
  VN1020_in1 <= VN_sign_in(6121) & VN_data_in(6121);
  VN1020_in2 <= VN_sign_in(6122) & VN_data_in(6122);
  VN1020_in3 <= VN_sign_in(6123) & VN_data_in(6123);
  VN1020_in4 <= VN_sign_in(6124) & VN_data_in(6124);
  VN1020_in5 <= VN_sign_in(6125) & VN_data_in(6125);
  VN1021_in0 <= VN_sign_in(6126) & VN_data_in(6126);
  VN1021_in1 <= VN_sign_in(6127) & VN_data_in(6127);
  VN1021_in2 <= VN_sign_in(6128) & VN_data_in(6128);
  VN1021_in3 <= VN_sign_in(6129) & VN_data_in(6129);
  VN1021_in4 <= VN_sign_in(6130) & VN_data_in(6130);
  VN1021_in5 <= VN_sign_in(6131) & VN_data_in(6131);
  VN1022_in0 <= VN_sign_in(6132) & VN_data_in(6132);
  VN1022_in1 <= VN_sign_in(6133) & VN_data_in(6133);
  VN1022_in2 <= VN_sign_in(6134) & VN_data_in(6134);
  VN1022_in3 <= VN_sign_in(6135) & VN_data_in(6135);
  VN1022_in4 <= VN_sign_in(6136) & VN_data_in(6136);
  VN1022_in5 <= VN_sign_in(6137) & VN_data_in(6137);
  VN1023_in0 <= VN_sign_in(6138) & VN_data_in(6138);
  VN1023_in1 <= VN_sign_in(6139) & VN_data_in(6139);
  VN1023_in2 <= VN_sign_in(6140) & VN_data_in(6140);
  VN1023_in3 <= VN_sign_in(6141) & VN_data_in(6141);
  VN1023_in4 <= VN_sign_in(6142) & VN_data_in(6142);
  VN1023_in5 <= VN_sign_in(6143) & VN_data_in(6143);
  VN1024_in0 <= VN_sign_in(6144) & VN_data_in(6144);
  VN1024_in1 <= VN_sign_in(6145) & VN_data_in(6145);
  VN1024_in2 <= VN_sign_in(6146) & VN_data_in(6146);
  VN1024_in3 <= VN_sign_in(6147) & VN_data_in(6147);
  VN1024_in4 <= VN_sign_in(6148) & VN_data_in(6148);
  VN1024_in5 <= VN_sign_in(6149) & VN_data_in(6149);
  VN1025_in0 <= VN_sign_in(6150) & VN_data_in(6150);
  VN1025_in1 <= VN_sign_in(6151) & VN_data_in(6151);
  VN1025_in2 <= VN_sign_in(6152) & VN_data_in(6152);
  VN1025_in3 <= VN_sign_in(6153) & VN_data_in(6153);
  VN1025_in4 <= VN_sign_in(6154) & VN_data_in(6154);
  VN1025_in5 <= VN_sign_in(6155) & VN_data_in(6155);
  VN1026_in0 <= VN_sign_in(6156) & VN_data_in(6156);
  VN1026_in1 <= VN_sign_in(6157) & VN_data_in(6157);
  VN1026_in2 <= VN_sign_in(6158) & VN_data_in(6158);
  VN1026_in3 <= VN_sign_in(6159) & VN_data_in(6159);
  VN1026_in4 <= VN_sign_in(6160) & VN_data_in(6160);
  VN1026_in5 <= VN_sign_in(6161) & VN_data_in(6161);
  VN1027_in0 <= VN_sign_in(6162) & VN_data_in(6162);
  VN1027_in1 <= VN_sign_in(6163) & VN_data_in(6163);
  VN1027_in2 <= VN_sign_in(6164) & VN_data_in(6164);
  VN1027_in3 <= VN_sign_in(6165) & VN_data_in(6165);
  VN1027_in4 <= VN_sign_in(6166) & VN_data_in(6166);
  VN1027_in5 <= VN_sign_in(6167) & VN_data_in(6167);
  VN1028_in0 <= VN_sign_in(6168) & VN_data_in(6168);
  VN1028_in1 <= VN_sign_in(6169) & VN_data_in(6169);
  VN1028_in2 <= VN_sign_in(6170) & VN_data_in(6170);
  VN1028_in3 <= VN_sign_in(6171) & VN_data_in(6171);
  VN1028_in4 <= VN_sign_in(6172) & VN_data_in(6172);
  VN1028_in5 <= VN_sign_in(6173) & VN_data_in(6173);
  VN1029_in0 <= VN_sign_in(6174) & VN_data_in(6174);
  VN1029_in1 <= VN_sign_in(6175) & VN_data_in(6175);
  VN1029_in2 <= VN_sign_in(6176) & VN_data_in(6176);
  VN1029_in3 <= VN_sign_in(6177) & VN_data_in(6177);
  VN1029_in4 <= VN_sign_in(6178) & VN_data_in(6178);
  VN1029_in5 <= VN_sign_in(6179) & VN_data_in(6179);
  VN1030_in0 <= VN_sign_in(6180) & VN_data_in(6180);
  VN1030_in1 <= VN_sign_in(6181) & VN_data_in(6181);
  VN1030_in2 <= VN_sign_in(6182) & VN_data_in(6182);
  VN1030_in3 <= VN_sign_in(6183) & VN_data_in(6183);
  VN1030_in4 <= VN_sign_in(6184) & VN_data_in(6184);
  VN1030_in5 <= VN_sign_in(6185) & VN_data_in(6185);
  VN1031_in0 <= VN_sign_in(6186) & VN_data_in(6186);
  VN1031_in1 <= VN_sign_in(6187) & VN_data_in(6187);
  VN1031_in2 <= VN_sign_in(6188) & VN_data_in(6188);
  VN1031_in3 <= VN_sign_in(6189) & VN_data_in(6189);
  VN1031_in4 <= VN_sign_in(6190) & VN_data_in(6190);
  VN1031_in5 <= VN_sign_in(6191) & VN_data_in(6191);
  VN1032_in0 <= VN_sign_in(6192) & VN_data_in(6192);
  VN1032_in1 <= VN_sign_in(6193) & VN_data_in(6193);
  VN1032_in2 <= VN_sign_in(6194) & VN_data_in(6194);
  VN1032_in3 <= VN_sign_in(6195) & VN_data_in(6195);
  VN1032_in4 <= VN_sign_in(6196) & VN_data_in(6196);
  VN1032_in5 <= VN_sign_in(6197) & VN_data_in(6197);
  VN1033_in0 <= VN_sign_in(6198) & VN_data_in(6198);
  VN1033_in1 <= VN_sign_in(6199) & VN_data_in(6199);
  VN1033_in2 <= VN_sign_in(6200) & VN_data_in(6200);
  VN1033_in3 <= VN_sign_in(6201) & VN_data_in(6201);
  VN1033_in4 <= VN_sign_in(6202) & VN_data_in(6202);
  VN1033_in5 <= VN_sign_in(6203) & VN_data_in(6203);
  VN1034_in0 <= VN_sign_in(6204) & VN_data_in(6204);
  VN1034_in1 <= VN_sign_in(6205) & VN_data_in(6205);
  VN1034_in2 <= VN_sign_in(6206) & VN_data_in(6206);
  VN1034_in3 <= VN_sign_in(6207) & VN_data_in(6207);
  VN1034_in4 <= VN_sign_in(6208) & VN_data_in(6208);
  VN1034_in5 <= VN_sign_in(6209) & VN_data_in(6209);
  VN1035_in0 <= VN_sign_in(6210) & VN_data_in(6210);
  VN1035_in1 <= VN_sign_in(6211) & VN_data_in(6211);
  VN1035_in2 <= VN_sign_in(6212) & VN_data_in(6212);
  VN1035_in3 <= VN_sign_in(6213) & VN_data_in(6213);
  VN1035_in4 <= VN_sign_in(6214) & VN_data_in(6214);
  VN1035_in5 <= VN_sign_in(6215) & VN_data_in(6215);
  VN1036_in0 <= VN_sign_in(6216) & VN_data_in(6216);
  VN1036_in1 <= VN_sign_in(6217) & VN_data_in(6217);
  VN1036_in2 <= VN_sign_in(6218) & VN_data_in(6218);
  VN1036_in3 <= VN_sign_in(6219) & VN_data_in(6219);
  VN1036_in4 <= VN_sign_in(6220) & VN_data_in(6220);
  VN1036_in5 <= VN_sign_in(6221) & VN_data_in(6221);
  VN1037_in0 <= VN_sign_in(6222) & VN_data_in(6222);
  VN1037_in1 <= VN_sign_in(6223) & VN_data_in(6223);
  VN1037_in2 <= VN_sign_in(6224) & VN_data_in(6224);
  VN1037_in3 <= VN_sign_in(6225) & VN_data_in(6225);
  VN1037_in4 <= VN_sign_in(6226) & VN_data_in(6226);
  VN1037_in5 <= VN_sign_in(6227) & VN_data_in(6227);
  VN1038_in0 <= VN_sign_in(6228) & VN_data_in(6228);
  VN1038_in1 <= VN_sign_in(6229) & VN_data_in(6229);
  VN1038_in2 <= VN_sign_in(6230) & VN_data_in(6230);
  VN1038_in3 <= VN_sign_in(6231) & VN_data_in(6231);
  VN1038_in4 <= VN_sign_in(6232) & VN_data_in(6232);
  VN1038_in5 <= VN_sign_in(6233) & VN_data_in(6233);
  VN1039_in0 <= VN_sign_in(6234) & VN_data_in(6234);
  VN1039_in1 <= VN_sign_in(6235) & VN_data_in(6235);
  VN1039_in2 <= VN_sign_in(6236) & VN_data_in(6236);
  VN1039_in3 <= VN_sign_in(6237) & VN_data_in(6237);
  VN1039_in4 <= VN_sign_in(6238) & VN_data_in(6238);
  VN1039_in5 <= VN_sign_in(6239) & VN_data_in(6239);
  VN1040_in0 <= VN_sign_in(6240) & VN_data_in(6240);
  VN1040_in1 <= VN_sign_in(6241) & VN_data_in(6241);
  VN1040_in2 <= VN_sign_in(6242) & VN_data_in(6242);
  VN1040_in3 <= VN_sign_in(6243) & VN_data_in(6243);
  VN1040_in4 <= VN_sign_in(6244) & VN_data_in(6244);
  VN1040_in5 <= VN_sign_in(6245) & VN_data_in(6245);
  VN1041_in0 <= VN_sign_in(6246) & VN_data_in(6246);
  VN1041_in1 <= VN_sign_in(6247) & VN_data_in(6247);
  VN1041_in2 <= VN_sign_in(6248) & VN_data_in(6248);
  VN1041_in3 <= VN_sign_in(6249) & VN_data_in(6249);
  VN1041_in4 <= VN_sign_in(6250) & VN_data_in(6250);
  VN1041_in5 <= VN_sign_in(6251) & VN_data_in(6251);
  VN1042_in0 <= VN_sign_in(6252) & VN_data_in(6252);
  VN1042_in1 <= VN_sign_in(6253) & VN_data_in(6253);
  VN1042_in2 <= VN_sign_in(6254) & VN_data_in(6254);
  VN1042_in3 <= VN_sign_in(6255) & VN_data_in(6255);
  VN1042_in4 <= VN_sign_in(6256) & VN_data_in(6256);
  VN1042_in5 <= VN_sign_in(6257) & VN_data_in(6257);
  VN1043_in0 <= VN_sign_in(6258) & VN_data_in(6258);
  VN1043_in1 <= VN_sign_in(6259) & VN_data_in(6259);
  VN1043_in2 <= VN_sign_in(6260) & VN_data_in(6260);
  VN1043_in3 <= VN_sign_in(6261) & VN_data_in(6261);
  VN1043_in4 <= VN_sign_in(6262) & VN_data_in(6262);
  VN1043_in5 <= VN_sign_in(6263) & VN_data_in(6263);
  VN1044_in0 <= VN_sign_in(6264) & VN_data_in(6264);
  VN1044_in1 <= VN_sign_in(6265) & VN_data_in(6265);
  VN1044_in2 <= VN_sign_in(6266) & VN_data_in(6266);
  VN1044_in3 <= VN_sign_in(6267) & VN_data_in(6267);
  VN1044_in4 <= VN_sign_in(6268) & VN_data_in(6268);
  VN1044_in5 <= VN_sign_in(6269) & VN_data_in(6269);
  VN1045_in0 <= VN_sign_in(6270) & VN_data_in(6270);
  VN1045_in1 <= VN_sign_in(6271) & VN_data_in(6271);
  VN1045_in2 <= VN_sign_in(6272) & VN_data_in(6272);
  VN1045_in3 <= VN_sign_in(6273) & VN_data_in(6273);
  VN1045_in4 <= VN_sign_in(6274) & VN_data_in(6274);
  VN1045_in5 <= VN_sign_in(6275) & VN_data_in(6275);
  VN1046_in0 <= VN_sign_in(6276) & VN_data_in(6276);
  VN1046_in1 <= VN_sign_in(6277) & VN_data_in(6277);
  VN1046_in2 <= VN_sign_in(6278) & VN_data_in(6278);
  VN1046_in3 <= VN_sign_in(6279) & VN_data_in(6279);
  VN1046_in4 <= VN_sign_in(6280) & VN_data_in(6280);
  VN1046_in5 <= VN_sign_in(6281) & VN_data_in(6281);
  VN1047_in0 <= VN_sign_in(6282) & VN_data_in(6282);
  VN1047_in1 <= VN_sign_in(6283) & VN_data_in(6283);
  VN1047_in2 <= VN_sign_in(6284) & VN_data_in(6284);
  VN1047_in3 <= VN_sign_in(6285) & VN_data_in(6285);
  VN1047_in4 <= VN_sign_in(6286) & VN_data_in(6286);
  VN1047_in5 <= VN_sign_in(6287) & VN_data_in(6287);
  VN1048_in0 <= VN_sign_in(6288) & VN_data_in(6288);
  VN1048_in1 <= VN_sign_in(6289) & VN_data_in(6289);
  VN1048_in2 <= VN_sign_in(6290) & VN_data_in(6290);
  VN1048_in3 <= VN_sign_in(6291) & VN_data_in(6291);
  VN1048_in4 <= VN_sign_in(6292) & VN_data_in(6292);
  VN1048_in5 <= VN_sign_in(6293) & VN_data_in(6293);
  VN1049_in0 <= VN_sign_in(6294) & VN_data_in(6294);
  VN1049_in1 <= VN_sign_in(6295) & VN_data_in(6295);
  VN1049_in2 <= VN_sign_in(6296) & VN_data_in(6296);
  VN1049_in3 <= VN_sign_in(6297) & VN_data_in(6297);
  VN1049_in4 <= VN_sign_in(6298) & VN_data_in(6298);
  VN1049_in5 <= VN_sign_in(6299) & VN_data_in(6299);
  VN1050_in0 <= VN_sign_in(6300) & VN_data_in(6300);
  VN1050_in1 <= VN_sign_in(6301) & VN_data_in(6301);
  VN1050_in2 <= VN_sign_in(6302) & VN_data_in(6302);
  VN1050_in3 <= VN_sign_in(6303) & VN_data_in(6303);
  VN1050_in4 <= VN_sign_in(6304) & VN_data_in(6304);
  VN1050_in5 <= VN_sign_in(6305) & VN_data_in(6305);
  VN1051_in0 <= VN_sign_in(6306) & VN_data_in(6306);
  VN1051_in1 <= VN_sign_in(6307) & VN_data_in(6307);
  VN1051_in2 <= VN_sign_in(6308) & VN_data_in(6308);
  VN1051_in3 <= VN_sign_in(6309) & VN_data_in(6309);
  VN1051_in4 <= VN_sign_in(6310) & VN_data_in(6310);
  VN1051_in5 <= VN_sign_in(6311) & VN_data_in(6311);
  VN1052_in0 <= VN_sign_in(6312) & VN_data_in(6312);
  VN1052_in1 <= VN_sign_in(6313) & VN_data_in(6313);
  VN1052_in2 <= VN_sign_in(6314) & VN_data_in(6314);
  VN1052_in3 <= VN_sign_in(6315) & VN_data_in(6315);
  VN1052_in4 <= VN_sign_in(6316) & VN_data_in(6316);
  VN1052_in5 <= VN_sign_in(6317) & VN_data_in(6317);
  VN1053_in0 <= VN_sign_in(6318) & VN_data_in(6318);
  VN1053_in1 <= VN_sign_in(6319) & VN_data_in(6319);
  VN1053_in2 <= VN_sign_in(6320) & VN_data_in(6320);
  VN1053_in3 <= VN_sign_in(6321) & VN_data_in(6321);
  VN1053_in4 <= VN_sign_in(6322) & VN_data_in(6322);
  VN1053_in5 <= VN_sign_in(6323) & VN_data_in(6323);
  VN1054_in0 <= VN_sign_in(6324) & VN_data_in(6324);
  VN1054_in1 <= VN_sign_in(6325) & VN_data_in(6325);
  VN1054_in2 <= VN_sign_in(6326) & VN_data_in(6326);
  VN1054_in3 <= VN_sign_in(6327) & VN_data_in(6327);
  VN1054_in4 <= VN_sign_in(6328) & VN_data_in(6328);
  VN1054_in5 <= VN_sign_in(6329) & VN_data_in(6329);
  VN1055_in0 <= VN_sign_in(6330) & VN_data_in(6330);
  VN1055_in1 <= VN_sign_in(6331) & VN_data_in(6331);
  VN1055_in2 <= VN_sign_in(6332) & VN_data_in(6332);
  VN1055_in3 <= VN_sign_in(6333) & VN_data_in(6333);
  VN1055_in4 <= VN_sign_in(6334) & VN_data_in(6334);
  VN1055_in5 <= VN_sign_in(6335) & VN_data_in(6335);
  VN1056_in0 <= VN_sign_in(6336) & VN_data_in(6336);
  VN1056_in1 <= VN_sign_in(6337) & VN_data_in(6337);
  VN1056_in2 <= VN_sign_in(6338) & VN_data_in(6338);
  VN1056_in3 <= VN_sign_in(6339) & VN_data_in(6339);
  VN1056_in4 <= VN_sign_in(6340) & VN_data_in(6340);
  VN1056_in5 <= VN_sign_in(6341) & VN_data_in(6341);
  VN1057_in0 <= VN_sign_in(6342) & VN_data_in(6342);
  VN1057_in1 <= VN_sign_in(6343) & VN_data_in(6343);
  VN1057_in2 <= VN_sign_in(6344) & VN_data_in(6344);
  VN1057_in3 <= VN_sign_in(6345) & VN_data_in(6345);
  VN1057_in4 <= VN_sign_in(6346) & VN_data_in(6346);
  VN1057_in5 <= VN_sign_in(6347) & VN_data_in(6347);
  VN1058_in0 <= VN_sign_in(6348) & VN_data_in(6348);
  VN1058_in1 <= VN_sign_in(6349) & VN_data_in(6349);
  VN1058_in2 <= VN_sign_in(6350) & VN_data_in(6350);
  VN1058_in3 <= VN_sign_in(6351) & VN_data_in(6351);
  VN1058_in4 <= VN_sign_in(6352) & VN_data_in(6352);
  VN1058_in5 <= VN_sign_in(6353) & VN_data_in(6353);
  VN1059_in0 <= VN_sign_in(6354) & VN_data_in(6354);
  VN1059_in1 <= VN_sign_in(6355) & VN_data_in(6355);
  VN1059_in2 <= VN_sign_in(6356) & VN_data_in(6356);
  VN1059_in3 <= VN_sign_in(6357) & VN_data_in(6357);
  VN1059_in4 <= VN_sign_in(6358) & VN_data_in(6358);
  VN1059_in5 <= VN_sign_in(6359) & VN_data_in(6359);
  VN1060_in0 <= VN_sign_in(6360) & VN_data_in(6360);
  VN1060_in1 <= VN_sign_in(6361) & VN_data_in(6361);
  VN1060_in2 <= VN_sign_in(6362) & VN_data_in(6362);
  VN1060_in3 <= VN_sign_in(6363) & VN_data_in(6363);
  VN1060_in4 <= VN_sign_in(6364) & VN_data_in(6364);
  VN1060_in5 <= VN_sign_in(6365) & VN_data_in(6365);
  VN1061_in0 <= VN_sign_in(6366) & VN_data_in(6366);
  VN1061_in1 <= VN_sign_in(6367) & VN_data_in(6367);
  VN1061_in2 <= VN_sign_in(6368) & VN_data_in(6368);
  VN1061_in3 <= VN_sign_in(6369) & VN_data_in(6369);
  VN1061_in4 <= VN_sign_in(6370) & VN_data_in(6370);
  VN1061_in5 <= VN_sign_in(6371) & VN_data_in(6371);
  VN1062_in0 <= VN_sign_in(6372) & VN_data_in(6372);
  VN1062_in1 <= VN_sign_in(6373) & VN_data_in(6373);
  VN1062_in2 <= VN_sign_in(6374) & VN_data_in(6374);
  VN1062_in3 <= VN_sign_in(6375) & VN_data_in(6375);
  VN1062_in4 <= VN_sign_in(6376) & VN_data_in(6376);
  VN1062_in5 <= VN_sign_in(6377) & VN_data_in(6377);
  VN1063_in0 <= VN_sign_in(6378) & VN_data_in(6378);
  VN1063_in1 <= VN_sign_in(6379) & VN_data_in(6379);
  VN1063_in2 <= VN_sign_in(6380) & VN_data_in(6380);
  VN1063_in3 <= VN_sign_in(6381) & VN_data_in(6381);
  VN1063_in4 <= VN_sign_in(6382) & VN_data_in(6382);
  VN1063_in5 <= VN_sign_in(6383) & VN_data_in(6383);
  VN1064_in0 <= VN_sign_in(6384) & VN_data_in(6384);
  VN1064_in1 <= VN_sign_in(6385) & VN_data_in(6385);
  VN1064_in2 <= VN_sign_in(6386) & VN_data_in(6386);
  VN1064_in3 <= VN_sign_in(6387) & VN_data_in(6387);
  VN1064_in4 <= VN_sign_in(6388) & VN_data_in(6388);
  VN1064_in5 <= VN_sign_in(6389) & VN_data_in(6389);
  VN1065_in0 <= VN_sign_in(6390) & VN_data_in(6390);
  VN1065_in1 <= VN_sign_in(6391) & VN_data_in(6391);
  VN1065_in2 <= VN_sign_in(6392) & VN_data_in(6392);
  VN1065_in3 <= VN_sign_in(6393) & VN_data_in(6393);
  VN1065_in4 <= VN_sign_in(6394) & VN_data_in(6394);
  VN1065_in5 <= VN_sign_in(6395) & VN_data_in(6395);
  VN1066_in0 <= VN_sign_in(6396) & VN_data_in(6396);
  VN1066_in1 <= VN_sign_in(6397) & VN_data_in(6397);
  VN1066_in2 <= VN_sign_in(6398) & VN_data_in(6398);
  VN1066_in3 <= VN_sign_in(6399) & VN_data_in(6399);
  VN1066_in4 <= VN_sign_in(6400) & VN_data_in(6400);
  VN1066_in5 <= VN_sign_in(6401) & VN_data_in(6401);
  VN1067_in0 <= VN_sign_in(6402) & VN_data_in(6402);
  VN1067_in1 <= VN_sign_in(6403) & VN_data_in(6403);
  VN1067_in2 <= VN_sign_in(6404) & VN_data_in(6404);
  VN1067_in3 <= VN_sign_in(6405) & VN_data_in(6405);
  VN1067_in4 <= VN_sign_in(6406) & VN_data_in(6406);
  VN1067_in5 <= VN_sign_in(6407) & VN_data_in(6407);
  VN1068_in0 <= VN_sign_in(6408) & VN_data_in(6408);
  VN1068_in1 <= VN_sign_in(6409) & VN_data_in(6409);
  VN1068_in2 <= VN_sign_in(6410) & VN_data_in(6410);
  VN1068_in3 <= VN_sign_in(6411) & VN_data_in(6411);
  VN1068_in4 <= VN_sign_in(6412) & VN_data_in(6412);
  VN1068_in5 <= VN_sign_in(6413) & VN_data_in(6413);
  VN1069_in0 <= VN_sign_in(6414) & VN_data_in(6414);
  VN1069_in1 <= VN_sign_in(6415) & VN_data_in(6415);
  VN1069_in2 <= VN_sign_in(6416) & VN_data_in(6416);
  VN1069_in3 <= VN_sign_in(6417) & VN_data_in(6417);
  VN1069_in4 <= VN_sign_in(6418) & VN_data_in(6418);
  VN1069_in5 <= VN_sign_in(6419) & VN_data_in(6419);
  VN1070_in0 <= VN_sign_in(6420) & VN_data_in(6420);
  VN1070_in1 <= VN_sign_in(6421) & VN_data_in(6421);
  VN1070_in2 <= VN_sign_in(6422) & VN_data_in(6422);
  VN1070_in3 <= VN_sign_in(6423) & VN_data_in(6423);
  VN1070_in4 <= VN_sign_in(6424) & VN_data_in(6424);
  VN1070_in5 <= VN_sign_in(6425) & VN_data_in(6425);
  VN1071_in0 <= VN_sign_in(6426) & VN_data_in(6426);
  VN1071_in1 <= VN_sign_in(6427) & VN_data_in(6427);
  VN1071_in2 <= VN_sign_in(6428) & VN_data_in(6428);
  VN1071_in3 <= VN_sign_in(6429) & VN_data_in(6429);
  VN1071_in4 <= VN_sign_in(6430) & VN_data_in(6430);
  VN1071_in5 <= VN_sign_in(6431) & VN_data_in(6431);
  VN1072_in0 <= VN_sign_in(6432) & VN_data_in(6432);
  VN1072_in1 <= VN_sign_in(6433) & VN_data_in(6433);
  VN1072_in2 <= VN_sign_in(6434) & VN_data_in(6434);
  VN1072_in3 <= VN_sign_in(6435) & VN_data_in(6435);
  VN1072_in4 <= VN_sign_in(6436) & VN_data_in(6436);
  VN1072_in5 <= VN_sign_in(6437) & VN_data_in(6437);
  VN1073_in0 <= VN_sign_in(6438) & VN_data_in(6438);
  VN1073_in1 <= VN_sign_in(6439) & VN_data_in(6439);
  VN1073_in2 <= VN_sign_in(6440) & VN_data_in(6440);
  VN1073_in3 <= VN_sign_in(6441) & VN_data_in(6441);
  VN1073_in4 <= VN_sign_in(6442) & VN_data_in(6442);
  VN1073_in5 <= VN_sign_in(6443) & VN_data_in(6443);
  VN1074_in0 <= VN_sign_in(6444) & VN_data_in(6444);
  VN1074_in1 <= VN_sign_in(6445) & VN_data_in(6445);
  VN1074_in2 <= VN_sign_in(6446) & VN_data_in(6446);
  VN1074_in3 <= VN_sign_in(6447) & VN_data_in(6447);
  VN1074_in4 <= VN_sign_in(6448) & VN_data_in(6448);
  VN1074_in5 <= VN_sign_in(6449) & VN_data_in(6449);
  VN1075_in0 <= VN_sign_in(6450) & VN_data_in(6450);
  VN1075_in1 <= VN_sign_in(6451) & VN_data_in(6451);
  VN1075_in2 <= VN_sign_in(6452) & VN_data_in(6452);
  VN1075_in3 <= VN_sign_in(6453) & VN_data_in(6453);
  VN1075_in4 <= VN_sign_in(6454) & VN_data_in(6454);
  VN1075_in5 <= VN_sign_in(6455) & VN_data_in(6455);
  VN1076_in0 <= VN_sign_in(6456) & VN_data_in(6456);
  VN1076_in1 <= VN_sign_in(6457) & VN_data_in(6457);
  VN1076_in2 <= VN_sign_in(6458) & VN_data_in(6458);
  VN1076_in3 <= VN_sign_in(6459) & VN_data_in(6459);
  VN1076_in4 <= VN_sign_in(6460) & VN_data_in(6460);
  VN1076_in5 <= VN_sign_in(6461) & VN_data_in(6461);
  VN1077_in0 <= VN_sign_in(6462) & VN_data_in(6462);
  VN1077_in1 <= VN_sign_in(6463) & VN_data_in(6463);
  VN1077_in2 <= VN_sign_in(6464) & VN_data_in(6464);
  VN1077_in3 <= VN_sign_in(6465) & VN_data_in(6465);
  VN1077_in4 <= VN_sign_in(6466) & VN_data_in(6466);
  VN1077_in5 <= VN_sign_in(6467) & VN_data_in(6467);
  VN1078_in0 <= VN_sign_in(6468) & VN_data_in(6468);
  VN1078_in1 <= VN_sign_in(6469) & VN_data_in(6469);
  VN1078_in2 <= VN_sign_in(6470) & VN_data_in(6470);
  VN1078_in3 <= VN_sign_in(6471) & VN_data_in(6471);
  VN1078_in4 <= VN_sign_in(6472) & VN_data_in(6472);
  VN1078_in5 <= VN_sign_in(6473) & VN_data_in(6473);
  VN1079_in0 <= VN_sign_in(6474) & VN_data_in(6474);
  VN1079_in1 <= VN_sign_in(6475) & VN_data_in(6475);
  VN1079_in2 <= VN_sign_in(6476) & VN_data_in(6476);
  VN1079_in3 <= VN_sign_in(6477) & VN_data_in(6477);
  VN1079_in4 <= VN_sign_in(6478) & VN_data_in(6478);
  VN1079_in5 <= VN_sign_in(6479) & VN_data_in(6479);
  VN1080_in0 <= VN_sign_in(6480) & VN_data_in(6480);
  VN1080_in1 <= VN_sign_in(6481) & VN_data_in(6481);
  VN1080_in2 <= VN_sign_in(6482) & VN_data_in(6482);
  VN1080_in3 <= VN_sign_in(6483) & VN_data_in(6483);
  VN1080_in4 <= VN_sign_in(6484) & VN_data_in(6484);
  VN1080_in5 <= VN_sign_in(6485) & VN_data_in(6485);
  VN1081_in0 <= VN_sign_in(6486) & VN_data_in(6486);
  VN1081_in1 <= VN_sign_in(6487) & VN_data_in(6487);
  VN1081_in2 <= VN_sign_in(6488) & VN_data_in(6488);
  VN1081_in3 <= VN_sign_in(6489) & VN_data_in(6489);
  VN1081_in4 <= VN_sign_in(6490) & VN_data_in(6490);
  VN1081_in5 <= VN_sign_in(6491) & VN_data_in(6491);
  VN1082_in0 <= VN_sign_in(6492) & VN_data_in(6492);
  VN1082_in1 <= VN_sign_in(6493) & VN_data_in(6493);
  VN1082_in2 <= VN_sign_in(6494) & VN_data_in(6494);
  VN1082_in3 <= VN_sign_in(6495) & VN_data_in(6495);
  VN1082_in4 <= VN_sign_in(6496) & VN_data_in(6496);
  VN1082_in5 <= VN_sign_in(6497) & VN_data_in(6497);
  VN1083_in0 <= VN_sign_in(6498) & VN_data_in(6498);
  VN1083_in1 <= VN_sign_in(6499) & VN_data_in(6499);
  VN1083_in2 <= VN_sign_in(6500) & VN_data_in(6500);
  VN1083_in3 <= VN_sign_in(6501) & VN_data_in(6501);
  VN1083_in4 <= VN_sign_in(6502) & VN_data_in(6502);
  VN1083_in5 <= VN_sign_in(6503) & VN_data_in(6503);
  VN1084_in0 <= VN_sign_in(6504) & VN_data_in(6504);
  VN1084_in1 <= VN_sign_in(6505) & VN_data_in(6505);
  VN1084_in2 <= VN_sign_in(6506) & VN_data_in(6506);
  VN1084_in3 <= VN_sign_in(6507) & VN_data_in(6507);
  VN1084_in4 <= VN_sign_in(6508) & VN_data_in(6508);
  VN1084_in5 <= VN_sign_in(6509) & VN_data_in(6509);
  VN1085_in0 <= VN_sign_in(6510) & VN_data_in(6510);
  VN1085_in1 <= VN_sign_in(6511) & VN_data_in(6511);
  VN1085_in2 <= VN_sign_in(6512) & VN_data_in(6512);
  VN1085_in3 <= VN_sign_in(6513) & VN_data_in(6513);
  VN1085_in4 <= VN_sign_in(6514) & VN_data_in(6514);
  VN1085_in5 <= VN_sign_in(6515) & VN_data_in(6515);
  VN1086_in0 <= VN_sign_in(6516) & VN_data_in(6516);
  VN1086_in1 <= VN_sign_in(6517) & VN_data_in(6517);
  VN1086_in2 <= VN_sign_in(6518) & VN_data_in(6518);
  VN1086_in3 <= VN_sign_in(6519) & VN_data_in(6519);
  VN1086_in4 <= VN_sign_in(6520) & VN_data_in(6520);
  VN1086_in5 <= VN_sign_in(6521) & VN_data_in(6521);
  VN1087_in0 <= VN_sign_in(6522) & VN_data_in(6522);
  VN1087_in1 <= VN_sign_in(6523) & VN_data_in(6523);
  VN1087_in2 <= VN_sign_in(6524) & VN_data_in(6524);
  VN1087_in3 <= VN_sign_in(6525) & VN_data_in(6525);
  VN1087_in4 <= VN_sign_in(6526) & VN_data_in(6526);
  VN1087_in5 <= VN_sign_in(6527) & VN_data_in(6527);
  VN1088_in0 <= VN_sign_in(6528) & VN_data_in(6528);
  VN1088_in1 <= VN_sign_in(6529) & VN_data_in(6529);
  VN1088_in2 <= VN_sign_in(6530) & VN_data_in(6530);
  VN1088_in3 <= VN_sign_in(6531) & VN_data_in(6531);
  VN1088_in4 <= VN_sign_in(6532) & VN_data_in(6532);
  VN1088_in5 <= VN_sign_in(6533) & VN_data_in(6533);
  VN1089_in0 <= VN_sign_in(6534) & VN_data_in(6534);
  VN1089_in1 <= VN_sign_in(6535) & VN_data_in(6535);
  VN1089_in2 <= VN_sign_in(6536) & VN_data_in(6536);
  VN1089_in3 <= VN_sign_in(6537) & VN_data_in(6537);
  VN1089_in4 <= VN_sign_in(6538) & VN_data_in(6538);
  VN1089_in5 <= VN_sign_in(6539) & VN_data_in(6539);
  VN1090_in0 <= VN_sign_in(6540) & VN_data_in(6540);
  VN1090_in1 <= VN_sign_in(6541) & VN_data_in(6541);
  VN1090_in2 <= VN_sign_in(6542) & VN_data_in(6542);
  VN1090_in3 <= VN_sign_in(6543) & VN_data_in(6543);
  VN1090_in4 <= VN_sign_in(6544) & VN_data_in(6544);
  VN1090_in5 <= VN_sign_in(6545) & VN_data_in(6545);
  VN1091_in0 <= VN_sign_in(6546) & VN_data_in(6546);
  VN1091_in1 <= VN_sign_in(6547) & VN_data_in(6547);
  VN1091_in2 <= VN_sign_in(6548) & VN_data_in(6548);
  VN1091_in3 <= VN_sign_in(6549) & VN_data_in(6549);
  VN1091_in4 <= VN_sign_in(6550) & VN_data_in(6550);
  VN1091_in5 <= VN_sign_in(6551) & VN_data_in(6551);
  VN1092_in0 <= VN_sign_in(6552) & VN_data_in(6552);
  VN1092_in1 <= VN_sign_in(6553) & VN_data_in(6553);
  VN1092_in2 <= VN_sign_in(6554) & VN_data_in(6554);
  VN1092_in3 <= VN_sign_in(6555) & VN_data_in(6555);
  VN1092_in4 <= VN_sign_in(6556) & VN_data_in(6556);
  VN1092_in5 <= VN_sign_in(6557) & VN_data_in(6557);
  VN1093_in0 <= VN_sign_in(6558) & VN_data_in(6558);
  VN1093_in1 <= VN_sign_in(6559) & VN_data_in(6559);
  VN1093_in2 <= VN_sign_in(6560) & VN_data_in(6560);
  VN1093_in3 <= VN_sign_in(6561) & VN_data_in(6561);
  VN1093_in4 <= VN_sign_in(6562) & VN_data_in(6562);
  VN1093_in5 <= VN_sign_in(6563) & VN_data_in(6563);
  VN1094_in0 <= VN_sign_in(6564) & VN_data_in(6564);
  VN1094_in1 <= VN_sign_in(6565) & VN_data_in(6565);
  VN1094_in2 <= VN_sign_in(6566) & VN_data_in(6566);
  VN1094_in3 <= VN_sign_in(6567) & VN_data_in(6567);
  VN1094_in4 <= VN_sign_in(6568) & VN_data_in(6568);
  VN1094_in5 <= VN_sign_in(6569) & VN_data_in(6569);
  VN1095_in0 <= VN_sign_in(6570) & VN_data_in(6570);
  VN1095_in1 <= VN_sign_in(6571) & VN_data_in(6571);
  VN1095_in2 <= VN_sign_in(6572) & VN_data_in(6572);
  VN1095_in3 <= VN_sign_in(6573) & VN_data_in(6573);
  VN1095_in4 <= VN_sign_in(6574) & VN_data_in(6574);
  VN1095_in5 <= VN_sign_in(6575) & VN_data_in(6575);
  VN1096_in0 <= VN_sign_in(6576) & VN_data_in(6576);
  VN1096_in1 <= VN_sign_in(6577) & VN_data_in(6577);
  VN1096_in2 <= VN_sign_in(6578) & VN_data_in(6578);
  VN1096_in3 <= VN_sign_in(6579) & VN_data_in(6579);
  VN1096_in4 <= VN_sign_in(6580) & VN_data_in(6580);
  VN1096_in5 <= VN_sign_in(6581) & VN_data_in(6581);
  VN1097_in0 <= VN_sign_in(6582) & VN_data_in(6582);
  VN1097_in1 <= VN_sign_in(6583) & VN_data_in(6583);
  VN1097_in2 <= VN_sign_in(6584) & VN_data_in(6584);
  VN1097_in3 <= VN_sign_in(6585) & VN_data_in(6585);
  VN1097_in4 <= VN_sign_in(6586) & VN_data_in(6586);
  VN1097_in5 <= VN_sign_in(6587) & VN_data_in(6587);
  VN1098_in0 <= VN_sign_in(6588) & VN_data_in(6588);
  VN1098_in1 <= VN_sign_in(6589) & VN_data_in(6589);
  VN1098_in2 <= VN_sign_in(6590) & VN_data_in(6590);
  VN1098_in3 <= VN_sign_in(6591) & VN_data_in(6591);
  VN1098_in4 <= VN_sign_in(6592) & VN_data_in(6592);
  VN1098_in5 <= VN_sign_in(6593) & VN_data_in(6593);
  VN1099_in0 <= VN_sign_in(6594) & VN_data_in(6594);
  VN1099_in1 <= VN_sign_in(6595) & VN_data_in(6595);
  VN1099_in2 <= VN_sign_in(6596) & VN_data_in(6596);
  VN1099_in3 <= VN_sign_in(6597) & VN_data_in(6597);
  VN1099_in4 <= VN_sign_in(6598) & VN_data_in(6598);
  VN1099_in5 <= VN_sign_in(6599) & VN_data_in(6599);
  VN1100_in0 <= VN_sign_in(6600) & VN_data_in(6600);
  VN1100_in1 <= VN_sign_in(6601) & VN_data_in(6601);
  VN1100_in2 <= VN_sign_in(6602) & VN_data_in(6602);
  VN1100_in3 <= VN_sign_in(6603) & VN_data_in(6603);
  VN1100_in4 <= VN_sign_in(6604) & VN_data_in(6604);
  VN1100_in5 <= VN_sign_in(6605) & VN_data_in(6605);
  VN1101_in0 <= VN_sign_in(6606) & VN_data_in(6606);
  VN1101_in1 <= VN_sign_in(6607) & VN_data_in(6607);
  VN1101_in2 <= VN_sign_in(6608) & VN_data_in(6608);
  VN1101_in3 <= VN_sign_in(6609) & VN_data_in(6609);
  VN1101_in4 <= VN_sign_in(6610) & VN_data_in(6610);
  VN1101_in5 <= VN_sign_in(6611) & VN_data_in(6611);
  VN1102_in0 <= VN_sign_in(6612) & VN_data_in(6612);
  VN1102_in1 <= VN_sign_in(6613) & VN_data_in(6613);
  VN1102_in2 <= VN_sign_in(6614) & VN_data_in(6614);
  VN1102_in3 <= VN_sign_in(6615) & VN_data_in(6615);
  VN1102_in4 <= VN_sign_in(6616) & VN_data_in(6616);
  VN1102_in5 <= VN_sign_in(6617) & VN_data_in(6617);
  VN1103_in0 <= VN_sign_in(6618) & VN_data_in(6618);
  VN1103_in1 <= VN_sign_in(6619) & VN_data_in(6619);
  VN1103_in2 <= VN_sign_in(6620) & VN_data_in(6620);
  VN1103_in3 <= VN_sign_in(6621) & VN_data_in(6621);
  VN1103_in4 <= VN_sign_in(6622) & VN_data_in(6622);
  VN1103_in5 <= VN_sign_in(6623) & VN_data_in(6623);
  VN1104_in0 <= VN_sign_in(6624) & VN_data_in(6624);
  VN1104_in1 <= VN_sign_in(6625) & VN_data_in(6625);
  VN1104_in2 <= VN_sign_in(6626) & VN_data_in(6626);
  VN1104_in3 <= VN_sign_in(6627) & VN_data_in(6627);
  VN1104_in4 <= VN_sign_in(6628) & VN_data_in(6628);
  VN1104_in5 <= VN_sign_in(6629) & VN_data_in(6629);
  VN1105_in0 <= VN_sign_in(6630) & VN_data_in(6630);
  VN1105_in1 <= VN_sign_in(6631) & VN_data_in(6631);
  VN1105_in2 <= VN_sign_in(6632) & VN_data_in(6632);
  VN1105_in3 <= VN_sign_in(6633) & VN_data_in(6633);
  VN1105_in4 <= VN_sign_in(6634) & VN_data_in(6634);
  VN1105_in5 <= VN_sign_in(6635) & VN_data_in(6635);
  VN1106_in0 <= VN_sign_in(6636) & VN_data_in(6636);
  VN1106_in1 <= VN_sign_in(6637) & VN_data_in(6637);
  VN1106_in2 <= VN_sign_in(6638) & VN_data_in(6638);
  VN1106_in3 <= VN_sign_in(6639) & VN_data_in(6639);
  VN1106_in4 <= VN_sign_in(6640) & VN_data_in(6640);
  VN1106_in5 <= VN_sign_in(6641) & VN_data_in(6641);
  VN1107_in0 <= VN_sign_in(6642) & VN_data_in(6642);
  VN1107_in1 <= VN_sign_in(6643) & VN_data_in(6643);
  VN1107_in2 <= VN_sign_in(6644) & VN_data_in(6644);
  VN1107_in3 <= VN_sign_in(6645) & VN_data_in(6645);
  VN1107_in4 <= VN_sign_in(6646) & VN_data_in(6646);
  VN1107_in5 <= VN_sign_in(6647) & VN_data_in(6647);
  VN1108_in0 <= VN_sign_in(6648) & VN_data_in(6648);
  VN1108_in1 <= VN_sign_in(6649) & VN_data_in(6649);
  VN1108_in2 <= VN_sign_in(6650) & VN_data_in(6650);
  VN1108_in3 <= VN_sign_in(6651) & VN_data_in(6651);
  VN1108_in4 <= VN_sign_in(6652) & VN_data_in(6652);
  VN1108_in5 <= VN_sign_in(6653) & VN_data_in(6653);
  VN1109_in0 <= VN_sign_in(6654) & VN_data_in(6654);
  VN1109_in1 <= VN_sign_in(6655) & VN_data_in(6655);
  VN1109_in2 <= VN_sign_in(6656) & VN_data_in(6656);
  VN1109_in3 <= VN_sign_in(6657) & VN_data_in(6657);
  VN1109_in4 <= VN_sign_in(6658) & VN_data_in(6658);
  VN1109_in5 <= VN_sign_in(6659) & VN_data_in(6659);
  VN1110_in0 <= VN_sign_in(6660) & VN_data_in(6660);
  VN1110_in1 <= VN_sign_in(6661) & VN_data_in(6661);
  VN1110_in2 <= VN_sign_in(6662) & VN_data_in(6662);
  VN1110_in3 <= VN_sign_in(6663) & VN_data_in(6663);
  VN1110_in4 <= VN_sign_in(6664) & VN_data_in(6664);
  VN1110_in5 <= VN_sign_in(6665) & VN_data_in(6665);
  VN1111_in0 <= VN_sign_in(6666) & VN_data_in(6666);
  VN1111_in1 <= VN_sign_in(6667) & VN_data_in(6667);
  VN1111_in2 <= VN_sign_in(6668) & VN_data_in(6668);
  VN1111_in3 <= VN_sign_in(6669) & VN_data_in(6669);
  VN1111_in4 <= VN_sign_in(6670) & VN_data_in(6670);
  VN1111_in5 <= VN_sign_in(6671) & VN_data_in(6671);
  VN1112_in0 <= VN_sign_in(6672) & VN_data_in(6672);
  VN1112_in1 <= VN_sign_in(6673) & VN_data_in(6673);
  VN1112_in2 <= VN_sign_in(6674) & VN_data_in(6674);
  VN1112_in3 <= VN_sign_in(6675) & VN_data_in(6675);
  VN1112_in4 <= VN_sign_in(6676) & VN_data_in(6676);
  VN1112_in5 <= VN_sign_in(6677) & VN_data_in(6677);
  VN1113_in0 <= VN_sign_in(6678) & VN_data_in(6678);
  VN1113_in1 <= VN_sign_in(6679) & VN_data_in(6679);
  VN1113_in2 <= VN_sign_in(6680) & VN_data_in(6680);
  VN1113_in3 <= VN_sign_in(6681) & VN_data_in(6681);
  VN1113_in4 <= VN_sign_in(6682) & VN_data_in(6682);
  VN1113_in5 <= VN_sign_in(6683) & VN_data_in(6683);
  VN1114_in0 <= VN_sign_in(6684) & VN_data_in(6684);
  VN1114_in1 <= VN_sign_in(6685) & VN_data_in(6685);
  VN1114_in2 <= VN_sign_in(6686) & VN_data_in(6686);
  VN1114_in3 <= VN_sign_in(6687) & VN_data_in(6687);
  VN1114_in4 <= VN_sign_in(6688) & VN_data_in(6688);
  VN1114_in5 <= VN_sign_in(6689) & VN_data_in(6689);
  VN1115_in0 <= VN_sign_in(6690) & VN_data_in(6690);
  VN1115_in1 <= VN_sign_in(6691) & VN_data_in(6691);
  VN1115_in2 <= VN_sign_in(6692) & VN_data_in(6692);
  VN1115_in3 <= VN_sign_in(6693) & VN_data_in(6693);
  VN1115_in4 <= VN_sign_in(6694) & VN_data_in(6694);
  VN1115_in5 <= VN_sign_in(6695) & VN_data_in(6695);
  VN1116_in0 <= VN_sign_in(6696) & VN_data_in(6696);
  VN1116_in1 <= VN_sign_in(6697) & VN_data_in(6697);
  VN1116_in2 <= VN_sign_in(6698) & VN_data_in(6698);
  VN1116_in3 <= VN_sign_in(6699) & VN_data_in(6699);
  VN1116_in4 <= VN_sign_in(6700) & VN_data_in(6700);
  VN1116_in5 <= VN_sign_in(6701) & VN_data_in(6701);
  VN1117_in0 <= VN_sign_in(6702) & VN_data_in(6702);
  VN1117_in1 <= VN_sign_in(6703) & VN_data_in(6703);
  VN1117_in2 <= VN_sign_in(6704) & VN_data_in(6704);
  VN1117_in3 <= VN_sign_in(6705) & VN_data_in(6705);
  VN1117_in4 <= VN_sign_in(6706) & VN_data_in(6706);
  VN1117_in5 <= VN_sign_in(6707) & VN_data_in(6707);
  VN1118_in0 <= VN_sign_in(6708) & VN_data_in(6708);
  VN1118_in1 <= VN_sign_in(6709) & VN_data_in(6709);
  VN1118_in2 <= VN_sign_in(6710) & VN_data_in(6710);
  VN1118_in3 <= VN_sign_in(6711) & VN_data_in(6711);
  VN1118_in4 <= VN_sign_in(6712) & VN_data_in(6712);
  VN1118_in5 <= VN_sign_in(6713) & VN_data_in(6713);
  VN1119_in0 <= VN_sign_in(6714) & VN_data_in(6714);
  VN1119_in1 <= VN_sign_in(6715) & VN_data_in(6715);
  VN1119_in2 <= VN_sign_in(6716) & VN_data_in(6716);
  VN1119_in3 <= VN_sign_in(6717) & VN_data_in(6717);
  VN1119_in4 <= VN_sign_in(6718) & VN_data_in(6718);
  VN1119_in5 <= VN_sign_in(6719) & VN_data_in(6719);
  VN1120_in0 <= VN_sign_in(6720) & VN_data_in(6720);
  VN1120_in1 <= VN_sign_in(6721) & VN_data_in(6721);
  VN1120_in2 <= VN_sign_in(6722) & VN_data_in(6722);
  VN1120_in3 <= VN_sign_in(6723) & VN_data_in(6723);
  VN1120_in4 <= VN_sign_in(6724) & VN_data_in(6724);
  VN1120_in5 <= VN_sign_in(6725) & VN_data_in(6725);
  VN1121_in0 <= VN_sign_in(6726) & VN_data_in(6726);
  VN1121_in1 <= VN_sign_in(6727) & VN_data_in(6727);
  VN1121_in2 <= VN_sign_in(6728) & VN_data_in(6728);
  VN1121_in3 <= VN_sign_in(6729) & VN_data_in(6729);
  VN1121_in4 <= VN_sign_in(6730) & VN_data_in(6730);
  VN1121_in5 <= VN_sign_in(6731) & VN_data_in(6731);
  VN1122_in0 <= VN_sign_in(6732) & VN_data_in(6732);
  VN1122_in1 <= VN_sign_in(6733) & VN_data_in(6733);
  VN1122_in2 <= VN_sign_in(6734) & VN_data_in(6734);
  VN1122_in3 <= VN_sign_in(6735) & VN_data_in(6735);
  VN1122_in4 <= VN_sign_in(6736) & VN_data_in(6736);
  VN1122_in5 <= VN_sign_in(6737) & VN_data_in(6737);
  VN1123_in0 <= VN_sign_in(6738) & VN_data_in(6738);
  VN1123_in1 <= VN_sign_in(6739) & VN_data_in(6739);
  VN1123_in2 <= VN_sign_in(6740) & VN_data_in(6740);
  VN1123_in3 <= VN_sign_in(6741) & VN_data_in(6741);
  VN1123_in4 <= VN_sign_in(6742) & VN_data_in(6742);
  VN1123_in5 <= VN_sign_in(6743) & VN_data_in(6743);
  VN1124_in0 <= VN_sign_in(6744) & VN_data_in(6744);
  VN1124_in1 <= VN_sign_in(6745) & VN_data_in(6745);
  VN1124_in2 <= VN_sign_in(6746) & VN_data_in(6746);
  VN1124_in3 <= VN_sign_in(6747) & VN_data_in(6747);
  VN1124_in4 <= VN_sign_in(6748) & VN_data_in(6748);
  VN1124_in5 <= VN_sign_in(6749) & VN_data_in(6749);
  VN1125_in0 <= VN_sign_in(6750) & VN_data_in(6750);
  VN1125_in1 <= VN_sign_in(6751) & VN_data_in(6751);
  VN1125_in2 <= VN_sign_in(6752) & VN_data_in(6752);
  VN1125_in3 <= VN_sign_in(6753) & VN_data_in(6753);
  VN1125_in4 <= VN_sign_in(6754) & VN_data_in(6754);
  VN1125_in5 <= VN_sign_in(6755) & VN_data_in(6755);
  VN1126_in0 <= VN_sign_in(6756) & VN_data_in(6756);
  VN1126_in1 <= VN_sign_in(6757) & VN_data_in(6757);
  VN1126_in2 <= VN_sign_in(6758) & VN_data_in(6758);
  VN1126_in3 <= VN_sign_in(6759) & VN_data_in(6759);
  VN1126_in4 <= VN_sign_in(6760) & VN_data_in(6760);
  VN1126_in5 <= VN_sign_in(6761) & VN_data_in(6761);
  VN1127_in0 <= VN_sign_in(6762) & VN_data_in(6762);
  VN1127_in1 <= VN_sign_in(6763) & VN_data_in(6763);
  VN1127_in2 <= VN_sign_in(6764) & VN_data_in(6764);
  VN1127_in3 <= VN_sign_in(6765) & VN_data_in(6765);
  VN1127_in4 <= VN_sign_in(6766) & VN_data_in(6766);
  VN1127_in5 <= VN_sign_in(6767) & VN_data_in(6767);
  VN1128_in0 <= VN_sign_in(6768) & VN_data_in(6768);
  VN1128_in1 <= VN_sign_in(6769) & VN_data_in(6769);
  VN1128_in2 <= VN_sign_in(6770) & VN_data_in(6770);
  VN1128_in3 <= VN_sign_in(6771) & VN_data_in(6771);
  VN1128_in4 <= VN_sign_in(6772) & VN_data_in(6772);
  VN1128_in5 <= VN_sign_in(6773) & VN_data_in(6773);
  VN1129_in0 <= VN_sign_in(6774) & VN_data_in(6774);
  VN1129_in1 <= VN_sign_in(6775) & VN_data_in(6775);
  VN1129_in2 <= VN_sign_in(6776) & VN_data_in(6776);
  VN1129_in3 <= VN_sign_in(6777) & VN_data_in(6777);
  VN1129_in4 <= VN_sign_in(6778) & VN_data_in(6778);
  VN1129_in5 <= VN_sign_in(6779) & VN_data_in(6779);
  VN1130_in0 <= VN_sign_in(6780) & VN_data_in(6780);
  VN1130_in1 <= VN_sign_in(6781) & VN_data_in(6781);
  VN1130_in2 <= VN_sign_in(6782) & VN_data_in(6782);
  VN1130_in3 <= VN_sign_in(6783) & VN_data_in(6783);
  VN1130_in4 <= VN_sign_in(6784) & VN_data_in(6784);
  VN1130_in5 <= VN_sign_in(6785) & VN_data_in(6785);
  VN1131_in0 <= VN_sign_in(6786) & VN_data_in(6786);
  VN1131_in1 <= VN_sign_in(6787) & VN_data_in(6787);
  VN1131_in2 <= VN_sign_in(6788) & VN_data_in(6788);
  VN1131_in3 <= VN_sign_in(6789) & VN_data_in(6789);
  VN1131_in4 <= VN_sign_in(6790) & VN_data_in(6790);
  VN1131_in5 <= VN_sign_in(6791) & VN_data_in(6791);
  VN1132_in0 <= VN_sign_in(6792) & VN_data_in(6792);
  VN1132_in1 <= VN_sign_in(6793) & VN_data_in(6793);
  VN1132_in2 <= VN_sign_in(6794) & VN_data_in(6794);
  VN1132_in3 <= VN_sign_in(6795) & VN_data_in(6795);
  VN1132_in4 <= VN_sign_in(6796) & VN_data_in(6796);
  VN1132_in5 <= VN_sign_in(6797) & VN_data_in(6797);
  VN1133_in0 <= VN_sign_in(6798) & VN_data_in(6798);
  VN1133_in1 <= VN_sign_in(6799) & VN_data_in(6799);
  VN1133_in2 <= VN_sign_in(6800) & VN_data_in(6800);
  VN1133_in3 <= VN_sign_in(6801) & VN_data_in(6801);
  VN1133_in4 <= VN_sign_in(6802) & VN_data_in(6802);
  VN1133_in5 <= VN_sign_in(6803) & VN_data_in(6803);
  VN1134_in0 <= VN_sign_in(6804) & VN_data_in(6804);
  VN1134_in1 <= VN_sign_in(6805) & VN_data_in(6805);
  VN1134_in2 <= VN_sign_in(6806) & VN_data_in(6806);
  VN1134_in3 <= VN_sign_in(6807) & VN_data_in(6807);
  VN1134_in4 <= VN_sign_in(6808) & VN_data_in(6808);
  VN1134_in5 <= VN_sign_in(6809) & VN_data_in(6809);
  VN1135_in0 <= VN_sign_in(6810) & VN_data_in(6810);
  VN1135_in1 <= VN_sign_in(6811) & VN_data_in(6811);
  VN1135_in2 <= VN_sign_in(6812) & VN_data_in(6812);
  VN1135_in3 <= VN_sign_in(6813) & VN_data_in(6813);
  VN1135_in4 <= VN_sign_in(6814) & VN_data_in(6814);
  VN1135_in5 <= VN_sign_in(6815) & VN_data_in(6815);
  VN1136_in0 <= VN_sign_in(6816) & VN_data_in(6816);
  VN1136_in1 <= VN_sign_in(6817) & VN_data_in(6817);
  VN1136_in2 <= VN_sign_in(6818) & VN_data_in(6818);
  VN1136_in3 <= VN_sign_in(6819) & VN_data_in(6819);
  VN1136_in4 <= VN_sign_in(6820) & VN_data_in(6820);
  VN1136_in5 <= VN_sign_in(6821) & VN_data_in(6821);
  VN1137_in0 <= VN_sign_in(6822) & VN_data_in(6822);
  VN1137_in1 <= VN_sign_in(6823) & VN_data_in(6823);
  VN1137_in2 <= VN_sign_in(6824) & VN_data_in(6824);
  VN1137_in3 <= VN_sign_in(6825) & VN_data_in(6825);
  VN1137_in4 <= VN_sign_in(6826) & VN_data_in(6826);
  VN1137_in5 <= VN_sign_in(6827) & VN_data_in(6827);
  VN1138_in0 <= VN_sign_in(6828) & VN_data_in(6828);
  VN1138_in1 <= VN_sign_in(6829) & VN_data_in(6829);
  VN1138_in2 <= VN_sign_in(6830) & VN_data_in(6830);
  VN1138_in3 <= VN_sign_in(6831) & VN_data_in(6831);
  VN1138_in4 <= VN_sign_in(6832) & VN_data_in(6832);
  VN1138_in5 <= VN_sign_in(6833) & VN_data_in(6833);
  VN1139_in0 <= VN_sign_in(6834) & VN_data_in(6834);
  VN1139_in1 <= VN_sign_in(6835) & VN_data_in(6835);
  VN1139_in2 <= VN_sign_in(6836) & VN_data_in(6836);
  VN1139_in3 <= VN_sign_in(6837) & VN_data_in(6837);
  VN1139_in4 <= VN_sign_in(6838) & VN_data_in(6838);
  VN1139_in5 <= VN_sign_in(6839) & VN_data_in(6839);
  VN1140_in0 <= VN_sign_in(6840) & VN_data_in(6840);
  VN1140_in1 <= VN_sign_in(6841) & VN_data_in(6841);
  VN1140_in2 <= VN_sign_in(6842) & VN_data_in(6842);
  VN1140_in3 <= VN_sign_in(6843) & VN_data_in(6843);
  VN1140_in4 <= VN_sign_in(6844) & VN_data_in(6844);
  VN1140_in5 <= VN_sign_in(6845) & VN_data_in(6845);
  VN1141_in0 <= VN_sign_in(6846) & VN_data_in(6846);
  VN1141_in1 <= VN_sign_in(6847) & VN_data_in(6847);
  VN1141_in2 <= VN_sign_in(6848) & VN_data_in(6848);
  VN1141_in3 <= VN_sign_in(6849) & VN_data_in(6849);
  VN1141_in4 <= VN_sign_in(6850) & VN_data_in(6850);
  VN1141_in5 <= VN_sign_in(6851) & VN_data_in(6851);
  VN1142_in0 <= VN_sign_in(6852) & VN_data_in(6852);
  VN1142_in1 <= VN_sign_in(6853) & VN_data_in(6853);
  VN1142_in2 <= VN_sign_in(6854) & VN_data_in(6854);
  VN1142_in3 <= VN_sign_in(6855) & VN_data_in(6855);
  VN1142_in4 <= VN_sign_in(6856) & VN_data_in(6856);
  VN1142_in5 <= VN_sign_in(6857) & VN_data_in(6857);
  VN1143_in0 <= VN_sign_in(6858) & VN_data_in(6858);
  VN1143_in1 <= VN_sign_in(6859) & VN_data_in(6859);
  VN1143_in2 <= VN_sign_in(6860) & VN_data_in(6860);
  VN1143_in3 <= VN_sign_in(6861) & VN_data_in(6861);
  VN1143_in4 <= VN_sign_in(6862) & VN_data_in(6862);
  VN1143_in5 <= VN_sign_in(6863) & VN_data_in(6863);
  VN1144_in0 <= VN_sign_in(6864) & VN_data_in(6864);
  VN1144_in1 <= VN_sign_in(6865) & VN_data_in(6865);
  VN1144_in2 <= VN_sign_in(6866) & VN_data_in(6866);
  VN1144_in3 <= VN_sign_in(6867) & VN_data_in(6867);
  VN1144_in4 <= VN_sign_in(6868) & VN_data_in(6868);
  VN1144_in5 <= VN_sign_in(6869) & VN_data_in(6869);
  VN1145_in0 <= VN_sign_in(6870) & VN_data_in(6870);
  VN1145_in1 <= VN_sign_in(6871) & VN_data_in(6871);
  VN1145_in2 <= VN_sign_in(6872) & VN_data_in(6872);
  VN1145_in3 <= VN_sign_in(6873) & VN_data_in(6873);
  VN1145_in4 <= VN_sign_in(6874) & VN_data_in(6874);
  VN1145_in5 <= VN_sign_in(6875) & VN_data_in(6875);
  VN1146_in0 <= VN_sign_in(6876) & VN_data_in(6876);
  VN1146_in1 <= VN_sign_in(6877) & VN_data_in(6877);
  VN1146_in2 <= VN_sign_in(6878) & VN_data_in(6878);
  VN1146_in3 <= VN_sign_in(6879) & VN_data_in(6879);
  VN1146_in4 <= VN_sign_in(6880) & VN_data_in(6880);
  VN1146_in5 <= VN_sign_in(6881) & VN_data_in(6881);
  VN1147_in0 <= VN_sign_in(6882) & VN_data_in(6882);
  VN1147_in1 <= VN_sign_in(6883) & VN_data_in(6883);
  VN1147_in2 <= VN_sign_in(6884) & VN_data_in(6884);
  VN1147_in3 <= VN_sign_in(6885) & VN_data_in(6885);
  VN1147_in4 <= VN_sign_in(6886) & VN_data_in(6886);
  VN1147_in5 <= VN_sign_in(6887) & VN_data_in(6887);
  VN1148_in0 <= VN_sign_in(6888) & VN_data_in(6888);
  VN1148_in1 <= VN_sign_in(6889) & VN_data_in(6889);
  VN1148_in2 <= VN_sign_in(6890) & VN_data_in(6890);
  VN1148_in3 <= VN_sign_in(6891) & VN_data_in(6891);
  VN1148_in4 <= VN_sign_in(6892) & VN_data_in(6892);
  VN1148_in5 <= VN_sign_in(6893) & VN_data_in(6893);
  VN1149_in0 <= VN_sign_in(6894) & VN_data_in(6894);
  VN1149_in1 <= VN_sign_in(6895) & VN_data_in(6895);
  VN1149_in2 <= VN_sign_in(6896) & VN_data_in(6896);
  VN1149_in3 <= VN_sign_in(6897) & VN_data_in(6897);
  VN1149_in4 <= VN_sign_in(6898) & VN_data_in(6898);
  VN1149_in5 <= VN_sign_in(6899) & VN_data_in(6899);
  VN1150_in0 <= VN_sign_in(6900) & VN_data_in(6900);
  VN1150_in1 <= VN_sign_in(6901) & VN_data_in(6901);
  VN1150_in2 <= VN_sign_in(6902) & VN_data_in(6902);
  VN1150_in3 <= VN_sign_in(6903) & VN_data_in(6903);
  VN1150_in4 <= VN_sign_in(6904) & VN_data_in(6904);
  VN1150_in5 <= VN_sign_in(6905) & VN_data_in(6905);
  VN1151_in0 <= VN_sign_in(6906) & VN_data_in(6906);
  VN1151_in1 <= VN_sign_in(6907) & VN_data_in(6907);
  VN1151_in2 <= VN_sign_in(6908) & VN_data_in(6908);
  VN1151_in3 <= VN_sign_in(6909) & VN_data_in(6909);
  VN1151_in4 <= VN_sign_in(6910) & VN_data_in(6910);
  VN1151_in5 <= VN_sign_in(6911) & VN_data_in(6911);
  VN1152_in0 <= VN_sign_in(6912) & VN_data_in(6912);
  VN1152_in1 <= VN_sign_in(6913) & VN_data_in(6913);
  VN1152_in2 <= VN_sign_in(6914) & VN_data_in(6914);
  VN1152_in3 <= VN_sign_in(6915) & VN_data_in(6915);
  VN1152_in4 <= VN_sign_in(6916) & VN_data_in(6916);
  VN1152_in5 <= VN_sign_in(6917) & VN_data_in(6917);
  VN1153_in0 <= VN_sign_in(6918) & VN_data_in(6918);
  VN1153_in1 <= VN_sign_in(6919) & VN_data_in(6919);
  VN1153_in2 <= VN_sign_in(6920) & VN_data_in(6920);
  VN1153_in3 <= VN_sign_in(6921) & VN_data_in(6921);
  VN1153_in4 <= VN_sign_in(6922) & VN_data_in(6922);
  VN1153_in5 <= VN_sign_in(6923) & VN_data_in(6923);
  VN1154_in0 <= VN_sign_in(6924) & VN_data_in(6924);
  VN1154_in1 <= VN_sign_in(6925) & VN_data_in(6925);
  VN1154_in2 <= VN_sign_in(6926) & VN_data_in(6926);
  VN1154_in3 <= VN_sign_in(6927) & VN_data_in(6927);
  VN1154_in4 <= VN_sign_in(6928) & VN_data_in(6928);
  VN1154_in5 <= VN_sign_in(6929) & VN_data_in(6929);
  VN1155_in0 <= VN_sign_in(6930) & VN_data_in(6930);
  VN1155_in1 <= VN_sign_in(6931) & VN_data_in(6931);
  VN1155_in2 <= VN_sign_in(6932) & VN_data_in(6932);
  VN1155_in3 <= VN_sign_in(6933) & VN_data_in(6933);
  VN1155_in4 <= VN_sign_in(6934) & VN_data_in(6934);
  VN1155_in5 <= VN_sign_in(6935) & VN_data_in(6935);
  VN1156_in0 <= VN_sign_in(6936) & VN_data_in(6936);
  VN1156_in1 <= VN_sign_in(6937) & VN_data_in(6937);
  VN1156_in2 <= VN_sign_in(6938) & VN_data_in(6938);
  VN1156_in3 <= VN_sign_in(6939) & VN_data_in(6939);
  VN1156_in4 <= VN_sign_in(6940) & VN_data_in(6940);
  VN1156_in5 <= VN_sign_in(6941) & VN_data_in(6941);
  VN1157_in0 <= VN_sign_in(6942) & VN_data_in(6942);
  VN1157_in1 <= VN_sign_in(6943) & VN_data_in(6943);
  VN1157_in2 <= VN_sign_in(6944) & VN_data_in(6944);
  VN1157_in3 <= VN_sign_in(6945) & VN_data_in(6945);
  VN1157_in4 <= VN_sign_in(6946) & VN_data_in(6946);
  VN1157_in5 <= VN_sign_in(6947) & VN_data_in(6947);
  VN1158_in0 <= VN_sign_in(6948) & VN_data_in(6948);
  VN1158_in1 <= VN_sign_in(6949) & VN_data_in(6949);
  VN1158_in2 <= VN_sign_in(6950) & VN_data_in(6950);
  VN1158_in3 <= VN_sign_in(6951) & VN_data_in(6951);
  VN1158_in4 <= VN_sign_in(6952) & VN_data_in(6952);
  VN1158_in5 <= VN_sign_in(6953) & VN_data_in(6953);
  VN1159_in0 <= VN_sign_in(6954) & VN_data_in(6954);
  VN1159_in1 <= VN_sign_in(6955) & VN_data_in(6955);
  VN1159_in2 <= VN_sign_in(6956) & VN_data_in(6956);
  VN1159_in3 <= VN_sign_in(6957) & VN_data_in(6957);
  VN1159_in4 <= VN_sign_in(6958) & VN_data_in(6958);
  VN1159_in5 <= VN_sign_in(6959) & VN_data_in(6959);
  VN1160_in0 <= VN_sign_in(6960) & VN_data_in(6960);
  VN1160_in1 <= VN_sign_in(6961) & VN_data_in(6961);
  VN1160_in2 <= VN_sign_in(6962) & VN_data_in(6962);
  VN1160_in3 <= VN_sign_in(6963) & VN_data_in(6963);
  VN1160_in4 <= VN_sign_in(6964) & VN_data_in(6964);
  VN1160_in5 <= VN_sign_in(6965) & VN_data_in(6965);
  VN1161_in0 <= VN_sign_in(6966) & VN_data_in(6966);
  VN1161_in1 <= VN_sign_in(6967) & VN_data_in(6967);
  VN1161_in2 <= VN_sign_in(6968) & VN_data_in(6968);
  VN1161_in3 <= VN_sign_in(6969) & VN_data_in(6969);
  VN1161_in4 <= VN_sign_in(6970) & VN_data_in(6970);
  VN1161_in5 <= VN_sign_in(6971) & VN_data_in(6971);
  VN1162_in0 <= VN_sign_in(6972) & VN_data_in(6972);
  VN1162_in1 <= VN_sign_in(6973) & VN_data_in(6973);
  VN1162_in2 <= VN_sign_in(6974) & VN_data_in(6974);
  VN1162_in3 <= VN_sign_in(6975) & VN_data_in(6975);
  VN1162_in4 <= VN_sign_in(6976) & VN_data_in(6976);
  VN1162_in5 <= VN_sign_in(6977) & VN_data_in(6977);
  VN1163_in0 <= VN_sign_in(6978) & VN_data_in(6978);
  VN1163_in1 <= VN_sign_in(6979) & VN_data_in(6979);
  VN1163_in2 <= VN_sign_in(6980) & VN_data_in(6980);
  VN1163_in3 <= VN_sign_in(6981) & VN_data_in(6981);
  VN1163_in4 <= VN_sign_in(6982) & VN_data_in(6982);
  VN1163_in5 <= VN_sign_in(6983) & VN_data_in(6983);
  VN1164_in0 <= VN_sign_in(6984) & VN_data_in(6984);
  VN1164_in1 <= VN_sign_in(6985) & VN_data_in(6985);
  VN1164_in2 <= VN_sign_in(6986) & VN_data_in(6986);
  VN1164_in3 <= VN_sign_in(6987) & VN_data_in(6987);
  VN1164_in4 <= VN_sign_in(6988) & VN_data_in(6988);
  VN1164_in5 <= VN_sign_in(6989) & VN_data_in(6989);
  VN1165_in0 <= VN_sign_in(6990) & VN_data_in(6990);
  VN1165_in1 <= VN_sign_in(6991) & VN_data_in(6991);
  VN1165_in2 <= VN_sign_in(6992) & VN_data_in(6992);
  VN1165_in3 <= VN_sign_in(6993) & VN_data_in(6993);
  VN1165_in4 <= VN_sign_in(6994) & VN_data_in(6994);
  VN1165_in5 <= VN_sign_in(6995) & VN_data_in(6995);
  VN1166_in0 <= VN_sign_in(6996) & VN_data_in(6996);
  VN1166_in1 <= VN_sign_in(6997) & VN_data_in(6997);
  VN1166_in2 <= VN_sign_in(6998) & VN_data_in(6998);
  VN1166_in3 <= VN_sign_in(6999) & VN_data_in(6999);
  VN1166_in4 <= VN_sign_in(7000) & VN_data_in(7000);
  VN1166_in5 <= VN_sign_in(7001) & VN_data_in(7001);
  VN1167_in0 <= VN_sign_in(7002) & VN_data_in(7002);
  VN1167_in1 <= VN_sign_in(7003) & VN_data_in(7003);
  VN1167_in2 <= VN_sign_in(7004) & VN_data_in(7004);
  VN1167_in3 <= VN_sign_in(7005) & VN_data_in(7005);
  VN1167_in4 <= VN_sign_in(7006) & VN_data_in(7006);
  VN1167_in5 <= VN_sign_in(7007) & VN_data_in(7007);
  VN1168_in0 <= VN_sign_in(7008) & VN_data_in(7008);
  VN1168_in1 <= VN_sign_in(7009) & VN_data_in(7009);
  VN1168_in2 <= VN_sign_in(7010) & VN_data_in(7010);
  VN1168_in3 <= VN_sign_in(7011) & VN_data_in(7011);
  VN1168_in4 <= VN_sign_in(7012) & VN_data_in(7012);
  VN1168_in5 <= VN_sign_in(7013) & VN_data_in(7013);
  VN1169_in0 <= VN_sign_in(7014) & VN_data_in(7014);
  VN1169_in1 <= VN_sign_in(7015) & VN_data_in(7015);
  VN1169_in2 <= VN_sign_in(7016) & VN_data_in(7016);
  VN1169_in3 <= VN_sign_in(7017) & VN_data_in(7017);
  VN1169_in4 <= VN_sign_in(7018) & VN_data_in(7018);
  VN1169_in5 <= VN_sign_in(7019) & VN_data_in(7019);
  VN1170_in0 <= VN_sign_in(7020) & VN_data_in(7020);
  VN1170_in1 <= VN_sign_in(7021) & VN_data_in(7021);
  VN1170_in2 <= VN_sign_in(7022) & VN_data_in(7022);
  VN1170_in3 <= VN_sign_in(7023) & VN_data_in(7023);
  VN1170_in4 <= VN_sign_in(7024) & VN_data_in(7024);
  VN1170_in5 <= VN_sign_in(7025) & VN_data_in(7025);
  VN1171_in0 <= VN_sign_in(7026) & VN_data_in(7026);
  VN1171_in1 <= VN_sign_in(7027) & VN_data_in(7027);
  VN1171_in2 <= VN_sign_in(7028) & VN_data_in(7028);
  VN1171_in3 <= VN_sign_in(7029) & VN_data_in(7029);
  VN1171_in4 <= VN_sign_in(7030) & VN_data_in(7030);
  VN1171_in5 <= VN_sign_in(7031) & VN_data_in(7031);
  VN1172_in0 <= VN_sign_in(7032) & VN_data_in(7032);
  VN1172_in1 <= VN_sign_in(7033) & VN_data_in(7033);
  VN1172_in2 <= VN_sign_in(7034) & VN_data_in(7034);
  VN1172_in3 <= VN_sign_in(7035) & VN_data_in(7035);
  VN1172_in4 <= VN_sign_in(7036) & VN_data_in(7036);
  VN1172_in5 <= VN_sign_in(7037) & VN_data_in(7037);
  VN1173_in0 <= VN_sign_in(7038) & VN_data_in(7038);
  VN1173_in1 <= VN_sign_in(7039) & VN_data_in(7039);
  VN1173_in2 <= VN_sign_in(7040) & VN_data_in(7040);
  VN1173_in3 <= VN_sign_in(7041) & VN_data_in(7041);
  VN1173_in4 <= VN_sign_in(7042) & VN_data_in(7042);
  VN1173_in5 <= VN_sign_in(7043) & VN_data_in(7043);
  VN1174_in0 <= VN_sign_in(7044) & VN_data_in(7044);
  VN1174_in1 <= VN_sign_in(7045) & VN_data_in(7045);
  VN1174_in2 <= VN_sign_in(7046) & VN_data_in(7046);
  VN1174_in3 <= VN_sign_in(7047) & VN_data_in(7047);
  VN1174_in4 <= VN_sign_in(7048) & VN_data_in(7048);
  VN1174_in5 <= VN_sign_in(7049) & VN_data_in(7049);
  VN1175_in0 <= VN_sign_in(7050) & VN_data_in(7050);
  VN1175_in1 <= VN_sign_in(7051) & VN_data_in(7051);
  VN1175_in2 <= VN_sign_in(7052) & VN_data_in(7052);
  VN1175_in3 <= VN_sign_in(7053) & VN_data_in(7053);
  VN1175_in4 <= VN_sign_in(7054) & VN_data_in(7054);
  VN1175_in5 <= VN_sign_in(7055) & VN_data_in(7055);
  VN1176_in0 <= VN_sign_in(7056) & VN_data_in(7056);
  VN1176_in1 <= VN_sign_in(7057) & VN_data_in(7057);
  VN1176_in2 <= VN_sign_in(7058) & VN_data_in(7058);
  VN1176_in3 <= VN_sign_in(7059) & VN_data_in(7059);
  VN1176_in4 <= VN_sign_in(7060) & VN_data_in(7060);
  VN1176_in5 <= VN_sign_in(7061) & VN_data_in(7061);
  VN1177_in0 <= VN_sign_in(7062) & VN_data_in(7062);
  VN1177_in1 <= VN_sign_in(7063) & VN_data_in(7063);
  VN1177_in2 <= VN_sign_in(7064) & VN_data_in(7064);
  VN1177_in3 <= VN_sign_in(7065) & VN_data_in(7065);
  VN1177_in4 <= VN_sign_in(7066) & VN_data_in(7066);
  VN1177_in5 <= VN_sign_in(7067) & VN_data_in(7067);
  VN1178_in0 <= VN_sign_in(7068) & VN_data_in(7068);
  VN1178_in1 <= VN_sign_in(7069) & VN_data_in(7069);
  VN1178_in2 <= VN_sign_in(7070) & VN_data_in(7070);
  VN1178_in3 <= VN_sign_in(7071) & VN_data_in(7071);
  VN1178_in4 <= VN_sign_in(7072) & VN_data_in(7072);
  VN1178_in5 <= VN_sign_in(7073) & VN_data_in(7073);
  VN1179_in0 <= VN_sign_in(7074) & VN_data_in(7074);
  VN1179_in1 <= VN_sign_in(7075) & VN_data_in(7075);
  VN1179_in2 <= VN_sign_in(7076) & VN_data_in(7076);
  VN1179_in3 <= VN_sign_in(7077) & VN_data_in(7077);
  VN1179_in4 <= VN_sign_in(7078) & VN_data_in(7078);
  VN1179_in5 <= VN_sign_in(7079) & VN_data_in(7079);
  VN1180_in0 <= VN_sign_in(7080) & VN_data_in(7080);
  VN1180_in1 <= VN_sign_in(7081) & VN_data_in(7081);
  VN1180_in2 <= VN_sign_in(7082) & VN_data_in(7082);
  VN1180_in3 <= VN_sign_in(7083) & VN_data_in(7083);
  VN1180_in4 <= VN_sign_in(7084) & VN_data_in(7084);
  VN1180_in5 <= VN_sign_in(7085) & VN_data_in(7085);
  VN1181_in0 <= VN_sign_in(7086) & VN_data_in(7086);
  VN1181_in1 <= VN_sign_in(7087) & VN_data_in(7087);
  VN1181_in2 <= VN_sign_in(7088) & VN_data_in(7088);
  VN1181_in3 <= VN_sign_in(7089) & VN_data_in(7089);
  VN1181_in4 <= VN_sign_in(7090) & VN_data_in(7090);
  VN1181_in5 <= VN_sign_in(7091) & VN_data_in(7091);
  VN1182_in0 <= VN_sign_in(7092) & VN_data_in(7092);
  VN1182_in1 <= VN_sign_in(7093) & VN_data_in(7093);
  VN1182_in2 <= VN_sign_in(7094) & VN_data_in(7094);
  VN1182_in3 <= VN_sign_in(7095) & VN_data_in(7095);
  VN1182_in4 <= VN_sign_in(7096) & VN_data_in(7096);
  VN1182_in5 <= VN_sign_in(7097) & VN_data_in(7097);
  VN1183_in0 <= VN_sign_in(7098) & VN_data_in(7098);
  VN1183_in1 <= VN_sign_in(7099) & VN_data_in(7099);
  VN1183_in2 <= VN_sign_in(7100) & VN_data_in(7100);
  VN1183_in3 <= VN_sign_in(7101) & VN_data_in(7101);
  VN1183_in4 <= VN_sign_in(7102) & VN_data_in(7102);
  VN1183_in5 <= VN_sign_in(7103) & VN_data_in(7103);
  VN1184_in0 <= VN_sign_in(7104) & VN_data_in(7104);
  VN1184_in1 <= VN_sign_in(7105) & VN_data_in(7105);
  VN1184_in2 <= VN_sign_in(7106) & VN_data_in(7106);
  VN1184_in3 <= VN_sign_in(7107) & VN_data_in(7107);
  VN1184_in4 <= VN_sign_in(7108) & VN_data_in(7108);
  VN1184_in5 <= VN_sign_in(7109) & VN_data_in(7109);
  VN1185_in0 <= VN_sign_in(7110) & VN_data_in(7110);
  VN1185_in1 <= VN_sign_in(7111) & VN_data_in(7111);
  VN1185_in2 <= VN_sign_in(7112) & VN_data_in(7112);
  VN1185_in3 <= VN_sign_in(7113) & VN_data_in(7113);
  VN1185_in4 <= VN_sign_in(7114) & VN_data_in(7114);
  VN1185_in5 <= VN_sign_in(7115) & VN_data_in(7115);
  VN1186_in0 <= VN_sign_in(7116) & VN_data_in(7116);
  VN1186_in1 <= VN_sign_in(7117) & VN_data_in(7117);
  VN1186_in2 <= VN_sign_in(7118) & VN_data_in(7118);
  VN1186_in3 <= VN_sign_in(7119) & VN_data_in(7119);
  VN1186_in4 <= VN_sign_in(7120) & VN_data_in(7120);
  VN1186_in5 <= VN_sign_in(7121) & VN_data_in(7121);
  VN1187_in0 <= VN_sign_in(7122) & VN_data_in(7122);
  VN1187_in1 <= VN_sign_in(7123) & VN_data_in(7123);
  VN1187_in2 <= VN_sign_in(7124) & VN_data_in(7124);
  VN1187_in3 <= VN_sign_in(7125) & VN_data_in(7125);
  VN1187_in4 <= VN_sign_in(7126) & VN_data_in(7126);
  VN1187_in5 <= VN_sign_in(7127) & VN_data_in(7127);
  VN1188_in0 <= VN_sign_in(7128) & VN_data_in(7128);
  VN1188_in1 <= VN_sign_in(7129) & VN_data_in(7129);
  VN1188_in2 <= VN_sign_in(7130) & VN_data_in(7130);
  VN1188_in3 <= VN_sign_in(7131) & VN_data_in(7131);
  VN1188_in4 <= VN_sign_in(7132) & VN_data_in(7132);
  VN1188_in5 <= VN_sign_in(7133) & VN_data_in(7133);
  VN1189_in0 <= VN_sign_in(7134) & VN_data_in(7134);
  VN1189_in1 <= VN_sign_in(7135) & VN_data_in(7135);
  VN1189_in2 <= VN_sign_in(7136) & VN_data_in(7136);
  VN1189_in3 <= VN_sign_in(7137) & VN_data_in(7137);
  VN1189_in4 <= VN_sign_in(7138) & VN_data_in(7138);
  VN1189_in5 <= VN_sign_in(7139) & VN_data_in(7139);
  VN1190_in0 <= VN_sign_in(7140) & VN_data_in(7140);
  VN1190_in1 <= VN_sign_in(7141) & VN_data_in(7141);
  VN1190_in2 <= VN_sign_in(7142) & VN_data_in(7142);
  VN1190_in3 <= VN_sign_in(7143) & VN_data_in(7143);
  VN1190_in4 <= VN_sign_in(7144) & VN_data_in(7144);
  VN1190_in5 <= VN_sign_in(7145) & VN_data_in(7145);
  VN1191_in0 <= VN_sign_in(7146) & VN_data_in(7146);
  VN1191_in1 <= VN_sign_in(7147) & VN_data_in(7147);
  VN1191_in2 <= VN_sign_in(7148) & VN_data_in(7148);
  VN1191_in3 <= VN_sign_in(7149) & VN_data_in(7149);
  VN1191_in4 <= VN_sign_in(7150) & VN_data_in(7150);
  VN1191_in5 <= VN_sign_in(7151) & VN_data_in(7151);
  VN1192_in0 <= VN_sign_in(7152) & VN_data_in(7152);
  VN1192_in1 <= VN_sign_in(7153) & VN_data_in(7153);
  VN1192_in2 <= VN_sign_in(7154) & VN_data_in(7154);
  VN1192_in3 <= VN_sign_in(7155) & VN_data_in(7155);
  VN1192_in4 <= VN_sign_in(7156) & VN_data_in(7156);
  VN1192_in5 <= VN_sign_in(7157) & VN_data_in(7157);
  VN1193_in0 <= VN_sign_in(7158) & VN_data_in(7158);
  VN1193_in1 <= VN_sign_in(7159) & VN_data_in(7159);
  VN1193_in2 <= VN_sign_in(7160) & VN_data_in(7160);
  VN1193_in3 <= VN_sign_in(7161) & VN_data_in(7161);
  VN1193_in4 <= VN_sign_in(7162) & VN_data_in(7162);
  VN1193_in5 <= VN_sign_in(7163) & VN_data_in(7163);
  VN1194_in0 <= VN_sign_in(7164) & VN_data_in(7164);
  VN1194_in1 <= VN_sign_in(7165) & VN_data_in(7165);
  VN1194_in2 <= VN_sign_in(7166) & VN_data_in(7166);
  VN1194_in3 <= VN_sign_in(7167) & VN_data_in(7167);
  VN1194_in4 <= VN_sign_in(7168) & VN_data_in(7168);
  VN1194_in5 <= VN_sign_in(7169) & VN_data_in(7169);
  VN1195_in0 <= VN_sign_in(7170) & VN_data_in(7170);
  VN1195_in1 <= VN_sign_in(7171) & VN_data_in(7171);
  VN1195_in2 <= VN_sign_in(7172) & VN_data_in(7172);
  VN1195_in3 <= VN_sign_in(7173) & VN_data_in(7173);
  VN1195_in4 <= VN_sign_in(7174) & VN_data_in(7174);
  VN1195_in5 <= VN_sign_in(7175) & VN_data_in(7175);
  VN1196_in0 <= VN_sign_in(7176) & VN_data_in(7176);
  VN1196_in1 <= VN_sign_in(7177) & VN_data_in(7177);
  VN1196_in2 <= VN_sign_in(7178) & VN_data_in(7178);
  VN1196_in3 <= VN_sign_in(7179) & VN_data_in(7179);
  VN1196_in4 <= VN_sign_in(7180) & VN_data_in(7180);
  VN1196_in5 <= VN_sign_in(7181) & VN_data_in(7181);
  VN1197_in0 <= VN_sign_in(7182) & VN_data_in(7182);
  VN1197_in1 <= VN_sign_in(7183) & VN_data_in(7183);
  VN1197_in2 <= VN_sign_in(7184) & VN_data_in(7184);
  VN1197_in3 <= VN_sign_in(7185) & VN_data_in(7185);
  VN1197_in4 <= VN_sign_in(7186) & VN_data_in(7186);
  VN1197_in5 <= VN_sign_in(7187) & VN_data_in(7187);
  VN1198_in0 <= VN_sign_in(7188) & VN_data_in(7188);
  VN1198_in1 <= VN_sign_in(7189) & VN_data_in(7189);
  VN1198_in2 <= VN_sign_in(7190) & VN_data_in(7190);
  VN1198_in3 <= VN_sign_in(7191) & VN_data_in(7191);
  VN1198_in4 <= VN_sign_in(7192) & VN_data_in(7192);
  VN1198_in5 <= VN_sign_in(7193) & VN_data_in(7193);
  VN1199_in0 <= VN_sign_in(7194) & VN_data_in(7194);
  VN1199_in1 <= VN_sign_in(7195) & VN_data_in(7195);
  VN1199_in2 <= VN_sign_in(7196) & VN_data_in(7196);
  VN1199_in3 <= VN_sign_in(7197) & VN_data_in(7197);
  VN1199_in4 <= VN_sign_in(7198) & VN_data_in(7198);
  VN1199_in5 <= VN_sign_in(7199) & VN_data_in(7199);
  VN1200_in0 <= VN_sign_in(7200) & VN_data_in(7200);
  VN1200_in1 <= VN_sign_in(7201) & VN_data_in(7201);
  VN1200_in2 <= VN_sign_in(7202) & VN_data_in(7202);
  VN1200_in3 <= VN_sign_in(7203) & VN_data_in(7203);
  VN1200_in4 <= VN_sign_in(7204) & VN_data_in(7204);
  VN1200_in5 <= VN_sign_in(7205) & VN_data_in(7205);
  VN1201_in0 <= VN_sign_in(7206) & VN_data_in(7206);
  VN1201_in1 <= VN_sign_in(7207) & VN_data_in(7207);
  VN1201_in2 <= VN_sign_in(7208) & VN_data_in(7208);
  VN1201_in3 <= VN_sign_in(7209) & VN_data_in(7209);
  VN1201_in4 <= VN_sign_in(7210) & VN_data_in(7210);
  VN1201_in5 <= VN_sign_in(7211) & VN_data_in(7211);
  VN1202_in0 <= VN_sign_in(7212) & VN_data_in(7212);
  VN1202_in1 <= VN_sign_in(7213) & VN_data_in(7213);
  VN1202_in2 <= VN_sign_in(7214) & VN_data_in(7214);
  VN1202_in3 <= VN_sign_in(7215) & VN_data_in(7215);
  VN1202_in4 <= VN_sign_in(7216) & VN_data_in(7216);
  VN1202_in5 <= VN_sign_in(7217) & VN_data_in(7217);
  VN1203_in0 <= VN_sign_in(7218) & VN_data_in(7218);
  VN1203_in1 <= VN_sign_in(7219) & VN_data_in(7219);
  VN1203_in2 <= VN_sign_in(7220) & VN_data_in(7220);
  VN1203_in3 <= VN_sign_in(7221) & VN_data_in(7221);
  VN1203_in4 <= VN_sign_in(7222) & VN_data_in(7222);
  VN1203_in5 <= VN_sign_in(7223) & VN_data_in(7223);
  VN1204_in0 <= VN_sign_in(7224) & VN_data_in(7224);
  VN1204_in1 <= VN_sign_in(7225) & VN_data_in(7225);
  VN1204_in2 <= VN_sign_in(7226) & VN_data_in(7226);
  VN1204_in3 <= VN_sign_in(7227) & VN_data_in(7227);
  VN1204_in4 <= VN_sign_in(7228) & VN_data_in(7228);
  VN1204_in5 <= VN_sign_in(7229) & VN_data_in(7229);
  VN1205_in0 <= VN_sign_in(7230) & VN_data_in(7230);
  VN1205_in1 <= VN_sign_in(7231) & VN_data_in(7231);
  VN1205_in2 <= VN_sign_in(7232) & VN_data_in(7232);
  VN1205_in3 <= VN_sign_in(7233) & VN_data_in(7233);
  VN1205_in4 <= VN_sign_in(7234) & VN_data_in(7234);
  VN1205_in5 <= VN_sign_in(7235) & VN_data_in(7235);
  VN1206_in0 <= VN_sign_in(7236) & VN_data_in(7236);
  VN1206_in1 <= VN_sign_in(7237) & VN_data_in(7237);
  VN1206_in2 <= VN_sign_in(7238) & VN_data_in(7238);
  VN1206_in3 <= VN_sign_in(7239) & VN_data_in(7239);
  VN1206_in4 <= VN_sign_in(7240) & VN_data_in(7240);
  VN1206_in5 <= VN_sign_in(7241) & VN_data_in(7241);
  VN1207_in0 <= VN_sign_in(7242) & VN_data_in(7242);
  VN1207_in1 <= VN_sign_in(7243) & VN_data_in(7243);
  VN1207_in2 <= VN_sign_in(7244) & VN_data_in(7244);
  VN1207_in3 <= VN_sign_in(7245) & VN_data_in(7245);
  VN1207_in4 <= VN_sign_in(7246) & VN_data_in(7246);
  VN1207_in5 <= VN_sign_in(7247) & VN_data_in(7247);
  VN1208_in0 <= VN_sign_in(7248) & VN_data_in(7248);
  VN1208_in1 <= VN_sign_in(7249) & VN_data_in(7249);
  VN1208_in2 <= VN_sign_in(7250) & VN_data_in(7250);
  VN1208_in3 <= VN_sign_in(7251) & VN_data_in(7251);
  VN1208_in4 <= VN_sign_in(7252) & VN_data_in(7252);
  VN1208_in5 <= VN_sign_in(7253) & VN_data_in(7253);
  VN1209_in0 <= VN_sign_in(7254) & VN_data_in(7254);
  VN1209_in1 <= VN_sign_in(7255) & VN_data_in(7255);
  VN1209_in2 <= VN_sign_in(7256) & VN_data_in(7256);
  VN1209_in3 <= VN_sign_in(7257) & VN_data_in(7257);
  VN1209_in4 <= VN_sign_in(7258) & VN_data_in(7258);
  VN1209_in5 <= VN_sign_in(7259) & VN_data_in(7259);
  VN1210_in0 <= VN_sign_in(7260) & VN_data_in(7260);
  VN1210_in1 <= VN_sign_in(7261) & VN_data_in(7261);
  VN1210_in2 <= VN_sign_in(7262) & VN_data_in(7262);
  VN1210_in3 <= VN_sign_in(7263) & VN_data_in(7263);
  VN1210_in4 <= VN_sign_in(7264) & VN_data_in(7264);
  VN1210_in5 <= VN_sign_in(7265) & VN_data_in(7265);
  VN1211_in0 <= VN_sign_in(7266) & VN_data_in(7266);
  VN1211_in1 <= VN_sign_in(7267) & VN_data_in(7267);
  VN1211_in2 <= VN_sign_in(7268) & VN_data_in(7268);
  VN1211_in3 <= VN_sign_in(7269) & VN_data_in(7269);
  VN1211_in4 <= VN_sign_in(7270) & VN_data_in(7270);
  VN1211_in5 <= VN_sign_in(7271) & VN_data_in(7271);
  VN1212_in0 <= VN_sign_in(7272) & VN_data_in(7272);
  VN1212_in1 <= VN_sign_in(7273) & VN_data_in(7273);
  VN1212_in2 <= VN_sign_in(7274) & VN_data_in(7274);
  VN1212_in3 <= VN_sign_in(7275) & VN_data_in(7275);
  VN1212_in4 <= VN_sign_in(7276) & VN_data_in(7276);
  VN1212_in5 <= VN_sign_in(7277) & VN_data_in(7277);
  VN1213_in0 <= VN_sign_in(7278) & VN_data_in(7278);
  VN1213_in1 <= VN_sign_in(7279) & VN_data_in(7279);
  VN1213_in2 <= VN_sign_in(7280) & VN_data_in(7280);
  VN1213_in3 <= VN_sign_in(7281) & VN_data_in(7281);
  VN1213_in4 <= VN_sign_in(7282) & VN_data_in(7282);
  VN1213_in5 <= VN_sign_in(7283) & VN_data_in(7283);
  VN1214_in0 <= VN_sign_in(7284) & VN_data_in(7284);
  VN1214_in1 <= VN_sign_in(7285) & VN_data_in(7285);
  VN1214_in2 <= VN_sign_in(7286) & VN_data_in(7286);
  VN1214_in3 <= VN_sign_in(7287) & VN_data_in(7287);
  VN1214_in4 <= VN_sign_in(7288) & VN_data_in(7288);
  VN1214_in5 <= VN_sign_in(7289) & VN_data_in(7289);
  VN1215_in0 <= VN_sign_in(7290) & VN_data_in(7290);
  VN1215_in1 <= VN_sign_in(7291) & VN_data_in(7291);
  VN1215_in2 <= VN_sign_in(7292) & VN_data_in(7292);
  VN1215_in3 <= VN_sign_in(7293) & VN_data_in(7293);
  VN1215_in4 <= VN_sign_in(7294) & VN_data_in(7294);
  VN1215_in5 <= VN_sign_in(7295) & VN_data_in(7295);
  VN1216_in0 <= VN_sign_in(7296) & VN_data_in(7296);
  VN1216_in1 <= VN_sign_in(7297) & VN_data_in(7297);
  VN1216_in2 <= VN_sign_in(7298) & VN_data_in(7298);
  VN1216_in3 <= VN_sign_in(7299) & VN_data_in(7299);
  VN1216_in4 <= VN_sign_in(7300) & VN_data_in(7300);
  VN1216_in5 <= VN_sign_in(7301) & VN_data_in(7301);
  VN1217_in0 <= VN_sign_in(7302) & VN_data_in(7302);
  VN1217_in1 <= VN_sign_in(7303) & VN_data_in(7303);
  VN1217_in2 <= VN_sign_in(7304) & VN_data_in(7304);
  VN1217_in3 <= VN_sign_in(7305) & VN_data_in(7305);
  VN1217_in4 <= VN_sign_in(7306) & VN_data_in(7306);
  VN1217_in5 <= VN_sign_in(7307) & VN_data_in(7307);
  VN1218_in0 <= VN_sign_in(7308) & VN_data_in(7308);
  VN1218_in1 <= VN_sign_in(7309) & VN_data_in(7309);
  VN1218_in2 <= VN_sign_in(7310) & VN_data_in(7310);
  VN1218_in3 <= VN_sign_in(7311) & VN_data_in(7311);
  VN1218_in4 <= VN_sign_in(7312) & VN_data_in(7312);
  VN1218_in5 <= VN_sign_in(7313) & VN_data_in(7313);
  VN1219_in0 <= VN_sign_in(7314) & VN_data_in(7314);
  VN1219_in1 <= VN_sign_in(7315) & VN_data_in(7315);
  VN1219_in2 <= VN_sign_in(7316) & VN_data_in(7316);
  VN1219_in3 <= VN_sign_in(7317) & VN_data_in(7317);
  VN1219_in4 <= VN_sign_in(7318) & VN_data_in(7318);
  VN1219_in5 <= VN_sign_in(7319) & VN_data_in(7319);
  VN1220_in0 <= VN_sign_in(7320) & VN_data_in(7320);
  VN1220_in1 <= VN_sign_in(7321) & VN_data_in(7321);
  VN1220_in2 <= VN_sign_in(7322) & VN_data_in(7322);
  VN1220_in3 <= VN_sign_in(7323) & VN_data_in(7323);
  VN1220_in4 <= VN_sign_in(7324) & VN_data_in(7324);
  VN1220_in5 <= VN_sign_in(7325) & VN_data_in(7325);
  VN1221_in0 <= VN_sign_in(7326) & VN_data_in(7326);
  VN1221_in1 <= VN_sign_in(7327) & VN_data_in(7327);
  VN1221_in2 <= VN_sign_in(7328) & VN_data_in(7328);
  VN1221_in3 <= VN_sign_in(7329) & VN_data_in(7329);
  VN1221_in4 <= VN_sign_in(7330) & VN_data_in(7330);
  VN1221_in5 <= VN_sign_in(7331) & VN_data_in(7331);
  VN1222_in0 <= VN_sign_in(7332) & VN_data_in(7332);
  VN1222_in1 <= VN_sign_in(7333) & VN_data_in(7333);
  VN1222_in2 <= VN_sign_in(7334) & VN_data_in(7334);
  VN1222_in3 <= VN_sign_in(7335) & VN_data_in(7335);
  VN1222_in4 <= VN_sign_in(7336) & VN_data_in(7336);
  VN1222_in5 <= VN_sign_in(7337) & VN_data_in(7337);
  VN1223_in0 <= VN_sign_in(7338) & VN_data_in(7338);
  VN1223_in1 <= VN_sign_in(7339) & VN_data_in(7339);
  VN1223_in2 <= VN_sign_in(7340) & VN_data_in(7340);
  VN1223_in3 <= VN_sign_in(7341) & VN_data_in(7341);
  VN1223_in4 <= VN_sign_in(7342) & VN_data_in(7342);
  VN1223_in5 <= VN_sign_in(7343) & VN_data_in(7343);
  VN1224_in0 <= VN_sign_in(7344) & VN_data_in(7344);
  VN1224_in1 <= VN_sign_in(7345) & VN_data_in(7345);
  VN1224_in2 <= VN_sign_in(7346) & VN_data_in(7346);
  VN1224_in3 <= VN_sign_in(7347) & VN_data_in(7347);
  VN1224_in4 <= VN_sign_in(7348) & VN_data_in(7348);
  VN1224_in5 <= VN_sign_in(7349) & VN_data_in(7349);
  VN1225_in0 <= VN_sign_in(7350) & VN_data_in(7350);
  VN1225_in1 <= VN_sign_in(7351) & VN_data_in(7351);
  VN1225_in2 <= VN_sign_in(7352) & VN_data_in(7352);
  VN1225_in3 <= VN_sign_in(7353) & VN_data_in(7353);
  VN1225_in4 <= VN_sign_in(7354) & VN_data_in(7354);
  VN1225_in5 <= VN_sign_in(7355) & VN_data_in(7355);
  VN1226_in0 <= VN_sign_in(7356) & VN_data_in(7356);
  VN1226_in1 <= VN_sign_in(7357) & VN_data_in(7357);
  VN1226_in2 <= VN_sign_in(7358) & VN_data_in(7358);
  VN1226_in3 <= VN_sign_in(7359) & VN_data_in(7359);
  VN1226_in4 <= VN_sign_in(7360) & VN_data_in(7360);
  VN1226_in5 <= VN_sign_in(7361) & VN_data_in(7361);
  VN1227_in0 <= VN_sign_in(7362) & VN_data_in(7362);
  VN1227_in1 <= VN_sign_in(7363) & VN_data_in(7363);
  VN1227_in2 <= VN_sign_in(7364) & VN_data_in(7364);
  VN1227_in3 <= VN_sign_in(7365) & VN_data_in(7365);
  VN1227_in4 <= VN_sign_in(7366) & VN_data_in(7366);
  VN1227_in5 <= VN_sign_in(7367) & VN_data_in(7367);
  VN1228_in0 <= VN_sign_in(7368) & VN_data_in(7368);
  VN1228_in1 <= VN_sign_in(7369) & VN_data_in(7369);
  VN1228_in2 <= VN_sign_in(7370) & VN_data_in(7370);
  VN1228_in3 <= VN_sign_in(7371) & VN_data_in(7371);
  VN1228_in4 <= VN_sign_in(7372) & VN_data_in(7372);
  VN1228_in5 <= VN_sign_in(7373) & VN_data_in(7373);
  VN1229_in0 <= VN_sign_in(7374) & VN_data_in(7374);
  VN1229_in1 <= VN_sign_in(7375) & VN_data_in(7375);
  VN1229_in2 <= VN_sign_in(7376) & VN_data_in(7376);
  VN1229_in3 <= VN_sign_in(7377) & VN_data_in(7377);
  VN1229_in4 <= VN_sign_in(7378) & VN_data_in(7378);
  VN1229_in5 <= VN_sign_in(7379) & VN_data_in(7379);
  VN1230_in0 <= VN_sign_in(7380) & VN_data_in(7380);
  VN1230_in1 <= VN_sign_in(7381) & VN_data_in(7381);
  VN1230_in2 <= VN_sign_in(7382) & VN_data_in(7382);
  VN1230_in3 <= VN_sign_in(7383) & VN_data_in(7383);
  VN1230_in4 <= VN_sign_in(7384) & VN_data_in(7384);
  VN1230_in5 <= VN_sign_in(7385) & VN_data_in(7385);
  VN1231_in0 <= VN_sign_in(7386) & VN_data_in(7386);
  VN1231_in1 <= VN_sign_in(7387) & VN_data_in(7387);
  VN1231_in2 <= VN_sign_in(7388) & VN_data_in(7388);
  VN1231_in3 <= VN_sign_in(7389) & VN_data_in(7389);
  VN1231_in4 <= VN_sign_in(7390) & VN_data_in(7390);
  VN1231_in5 <= VN_sign_in(7391) & VN_data_in(7391);
  VN1232_in0 <= VN_sign_in(7392) & VN_data_in(7392);
  VN1232_in1 <= VN_sign_in(7393) & VN_data_in(7393);
  VN1232_in2 <= VN_sign_in(7394) & VN_data_in(7394);
  VN1232_in3 <= VN_sign_in(7395) & VN_data_in(7395);
  VN1232_in4 <= VN_sign_in(7396) & VN_data_in(7396);
  VN1232_in5 <= VN_sign_in(7397) & VN_data_in(7397);
  VN1233_in0 <= VN_sign_in(7398) & VN_data_in(7398);
  VN1233_in1 <= VN_sign_in(7399) & VN_data_in(7399);
  VN1233_in2 <= VN_sign_in(7400) & VN_data_in(7400);
  VN1233_in3 <= VN_sign_in(7401) & VN_data_in(7401);
  VN1233_in4 <= VN_sign_in(7402) & VN_data_in(7402);
  VN1233_in5 <= VN_sign_in(7403) & VN_data_in(7403);
  VN1234_in0 <= VN_sign_in(7404) & VN_data_in(7404);
  VN1234_in1 <= VN_sign_in(7405) & VN_data_in(7405);
  VN1234_in2 <= VN_sign_in(7406) & VN_data_in(7406);
  VN1234_in3 <= VN_sign_in(7407) & VN_data_in(7407);
  VN1234_in4 <= VN_sign_in(7408) & VN_data_in(7408);
  VN1234_in5 <= VN_sign_in(7409) & VN_data_in(7409);
  VN1235_in0 <= VN_sign_in(7410) & VN_data_in(7410);
  VN1235_in1 <= VN_sign_in(7411) & VN_data_in(7411);
  VN1235_in2 <= VN_sign_in(7412) & VN_data_in(7412);
  VN1235_in3 <= VN_sign_in(7413) & VN_data_in(7413);
  VN1235_in4 <= VN_sign_in(7414) & VN_data_in(7414);
  VN1235_in5 <= VN_sign_in(7415) & VN_data_in(7415);
  VN1236_in0 <= VN_sign_in(7416) & VN_data_in(7416);
  VN1236_in1 <= VN_sign_in(7417) & VN_data_in(7417);
  VN1236_in2 <= VN_sign_in(7418) & VN_data_in(7418);
  VN1236_in3 <= VN_sign_in(7419) & VN_data_in(7419);
  VN1236_in4 <= VN_sign_in(7420) & VN_data_in(7420);
  VN1236_in5 <= VN_sign_in(7421) & VN_data_in(7421);
  VN1237_in0 <= VN_sign_in(7422) & VN_data_in(7422);
  VN1237_in1 <= VN_sign_in(7423) & VN_data_in(7423);
  VN1237_in2 <= VN_sign_in(7424) & VN_data_in(7424);
  VN1237_in3 <= VN_sign_in(7425) & VN_data_in(7425);
  VN1237_in4 <= VN_sign_in(7426) & VN_data_in(7426);
  VN1237_in5 <= VN_sign_in(7427) & VN_data_in(7427);
  VN1238_in0 <= VN_sign_in(7428) & VN_data_in(7428);
  VN1238_in1 <= VN_sign_in(7429) & VN_data_in(7429);
  VN1238_in2 <= VN_sign_in(7430) & VN_data_in(7430);
  VN1238_in3 <= VN_sign_in(7431) & VN_data_in(7431);
  VN1238_in4 <= VN_sign_in(7432) & VN_data_in(7432);
  VN1238_in5 <= VN_sign_in(7433) & VN_data_in(7433);
  VN1239_in0 <= VN_sign_in(7434) & VN_data_in(7434);
  VN1239_in1 <= VN_sign_in(7435) & VN_data_in(7435);
  VN1239_in2 <= VN_sign_in(7436) & VN_data_in(7436);
  VN1239_in3 <= VN_sign_in(7437) & VN_data_in(7437);
  VN1239_in4 <= VN_sign_in(7438) & VN_data_in(7438);
  VN1239_in5 <= VN_sign_in(7439) & VN_data_in(7439);
  VN1240_in0 <= VN_sign_in(7440) & VN_data_in(7440);
  VN1240_in1 <= VN_sign_in(7441) & VN_data_in(7441);
  VN1240_in2 <= VN_sign_in(7442) & VN_data_in(7442);
  VN1240_in3 <= VN_sign_in(7443) & VN_data_in(7443);
  VN1240_in4 <= VN_sign_in(7444) & VN_data_in(7444);
  VN1240_in5 <= VN_sign_in(7445) & VN_data_in(7445);
  VN1241_in0 <= VN_sign_in(7446) & VN_data_in(7446);
  VN1241_in1 <= VN_sign_in(7447) & VN_data_in(7447);
  VN1241_in2 <= VN_sign_in(7448) & VN_data_in(7448);
  VN1241_in3 <= VN_sign_in(7449) & VN_data_in(7449);
  VN1241_in4 <= VN_sign_in(7450) & VN_data_in(7450);
  VN1241_in5 <= VN_sign_in(7451) & VN_data_in(7451);
  VN1242_in0 <= VN_sign_in(7452) & VN_data_in(7452);
  VN1242_in1 <= VN_sign_in(7453) & VN_data_in(7453);
  VN1242_in2 <= VN_sign_in(7454) & VN_data_in(7454);
  VN1242_in3 <= VN_sign_in(7455) & VN_data_in(7455);
  VN1242_in4 <= VN_sign_in(7456) & VN_data_in(7456);
  VN1242_in5 <= VN_sign_in(7457) & VN_data_in(7457);
  VN1243_in0 <= VN_sign_in(7458) & VN_data_in(7458);
  VN1243_in1 <= VN_sign_in(7459) & VN_data_in(7459);
  VN1243_in2 <= VN_sign_in(7460) & VN_data_in(7460);
  VN1243_in3 <= VN_sign_in(7461) & VN_data_in(7461);
  VN1243_in4 <= VN_sign_in(7462) & VN_data_in(7462);
  VN1243_in5 <= VN_sign_in(7463) & VN_data_in(7463);
  VN1244_in0 <= VN_sign_in(7464) & VN_data_in(7464);
  VN1244_in1 <= VN_sign_in(7465) & VN_data_in(7465);
  VN1244_in2 <= VN_sign_in(7466) & VN_data_in(7466);
  VN1244_in3 <= VN_sign_in(7467) & VN_data_in(7467);
  VN1244_in4 <= VN_sign_in(7468) & VN_data_in(7468);
  VN1244_in5 <= VN_sign_in(7469) & VN_data_in(7469);
  VN1245_in0 <= VN_sign_in(7470) & VN_data_in(7470);
  VN1245_in1 <= VN_sign_in(7471) & VN_data_in(7471);
  VN1245_in2 <= VN_sign_in(7472) & VN_data_in(7472);
  VN1245_in3 <= VN_sign_in(7473) & VN_data_in(7473);
  VN1245_in4 <= VN_sign_in(7474) & VN_data_in(7474);
  VN1245_in5 <= VN_sign_in(7475) & VN_data_in(7475);
  VN1246_in0 <= VN_sign_in(7476) & VN_data_in(7476);
  VN1246_in1 <= VN_sign_in(7477) & VN_data_in(7477);
  VN1246_in2 <= VN_sign_in(7478) & VN_data_in(7478);
  VN1246_in3 <= VN_sign_in(7479) & VN_data_in(7479);
  VN1246_in4 <= VN_sign_in(7480) & VN_data_in(7480);
  VN1246_in5 <= VN_sign_in(7481) & VN_data_in(7481);
  VN1247_in0 <= VN_sign_in(7482) & VN_data_in(7482);
  VN1247_in1 <= VN_sign_in(7483) & VN_data_in(7483);
  VN1247_in2 <= VN_sign_in(7484) & VN_data_in(7484);
  VN1247_in3 <= VN_sign_in(7485) & VN_data_in(7485);
  VN1247_in4 <= VN_sign_in(7486) & VN_data_in(7486);
  VN1247_in5 <= VN_sign_in(7487) & VN_data_in(7487);
  VN1248_in0 <= VN_sign_in(7488) & VN_data_in(7488);
  VN1248_in1 <= VN_sign_in(7489) & VN_data_in(7489);
  VN1248_in2 <= VN_sign_in(7490) & VN_data_in(7490);
  VN1248_in3 <= VN_sign_in(7491) & VN_data_in(7491);
  VN1248_in4 <= VN_sign_in(7492) & VN_data_in(7492);
  VN1248_in5 <= VN_sign_in(7493) & VN_data_in(7493);
  VN1249_in0 <= VN_sign_in(7494) & VN_data_in(7494);
  VN1249_in1 <= VN_sign_in(7495) & VN_data_in(7495);
  VN1249_in2 <= VN_sign_in(7496) & VN_data_in(7496);
  VN1249_in3 <= VN_sign_in(7497) & VN_data_in(7497);
  VN1249_in4 <= VN_sign_in(7498) & VN_data_in(7498);
  VN1249_in5 <= VN_sign_in(7499) & VN_data_in(7499);
  VN1250_in0 <= VN_sign_in(7500) & VN_data_in(7500);
  VN1250_in1 <= VN_sign_in(7501) & VN_data_in(7501);
  VN1250_in2 <= VN_sign_in(7502) & VN_data_in(7502);
  VN1250_in3 <= VN_sign_in(7503) & VN_data_in(7503);
  VN1250_in4 <= VN_sign_in(7504) & VN_data_in(7504);
  VN1250_in5 <= VN_sign_in(7505) & VN_data_in(7505);
  VN1251_in0 <= VN_sign_in(7506) & VN_data_in(7506);
  VN1251_in1 <= VN_sign_in(7507) & VN_data_in(7507);
  VN1251_in2 <= VN_sign_in(7508) & VN_data_in(7508);
  VN1251_in3 <= VN_sign_in(7509) & VN_data_in(7509);
  VN1251_in4 <= VN_sign_in(7510) & VN_data_in(7510);
  VN1251_in5 <= VN_sign_in(7511) & VN_data_in(7511);
  VN1252_in0 <= VN_sign_in(7512) & VN_data_in(7512);
  VN1252_in1 <= VN_sign_in(7513) & VN_data_in(7513);
  VN1252_in2 <= VN_sign_in(7514) & VN_data_in(7514);
  VN1252_in3 <= VN_sign_in(7515) & VN_data_in(7515);
  VN1252_in4 <= VN_sign_in(7516) & VN_data_in(7516);
  VN1252_in5 <= VN_sign_in(7517) & VN_data_in(7517);
  VN1253_in0 <= VN_sign_in(7518) & VN_data_in(7518);
  VN1253_in1 <= VN_sign_in(7519) & VN_data_in(7519);
  VN1253_in2 <= VN_sign_in(7520) & VN_data_in(7520);
  VN1253_in3 <= VN_sign_in(7521) & VN_data_in(7521);
  VN1253_in4 <= VN_sign_in(7522) & VN_data_in(7522);
  VN1253_in5 <= VN_sign_in(7523) & VN_data_in(7523);
  VN1254_in0 <= VN_sign_in(7524) & VN_data_in(7524);
  VN1254_in1 <= VN_sign_in(7525) & VN_data_in(7525);
  VN1254_in2 <= VN_sign_in(7526) & VN_data_in(7526);
  VN1254_in3 <= VN_sign_in(7527) & VN_data_in(7527);
  VN1254_in4 <= VN_sign_in(7528) & VN_data_in(7528);
  VN1254_in5 <= VN_sign_in(7529) & VN_data_in(7529);
  VN1255_in0 <= VN_sign_in(7530) & VN_data_in(7530);
  VN1255_in1 <= VN_sign_in(7531) & VN_data_in(7531);
  VN1255_in2 <= VN_sign_in(7532) & VN_data_in(7532);
  VN1255_in3 <= VN_sign_in(7533) & VN_data_in(7533);
  VN1255_in4 <= VN_sign_in(7534) & VN_data_in(7534);
  VN1255_in5 <= VN_sign_in(7535) & VN_data_in(7535);
  VN1256_in0 <= VN_sign_in(7536) & VN_data_in(7536);
  VN1256_in1 <= VN_sign_in(7537) & VN_data_in(7537);
  VN1256_in2 <= VN_sign_in(7538) & VN_data_in(7538);
  VN1256_in3 <= VN_sign_in(7539) & VN_data_in(7539);
  VN1256_in4 <= VN_sign_in(7540) & VN_data_in(7540);
  VN1256_in5 <= VN_sign_in(7541) & VN_data_in(7541);
  VN1257_in0 <= VN_sign_in(7542) & VN_data_in(7542);
  VN1257_in1 <= VN_sign_in(7543) & VN_data_in(7543);
  VN1257_in2 <= VN_sign_in(7544) & VN_data_in(7544);
  VN1257_in3 <= VN_sign_in(7545) & VN_data_in(7545);
  VN1257_in4 <= VN_sign_in(7546) & VN_data_in(7546);
  VN1257_in5 <= VN_sign_in(7547) & VN_data_in(7547);
  VN1258_in0 <= VN_sign_in(7548) & VN_data_in(7548);
  VN1258_in1 <= VN_sign_in(7549) & VN_data_in(7549);
  VN1258_in2 <= VN_sign_in(7550) & VN_data_in(7550);
  VN1258_in3 <= VN_sign_in(7551) & VN_data_in(7551);
  VN1258_in4 <= VN_sign_in(7552) & VN_data_in(7552);
  VN1258_in5 <= VN_sign_in(7553) & VN_data_in(7553);
  VN1259_in0 <= VN_sign_in(7554) & VN_data_in(7554);
  VN1259_in1 <= VN_sign_in(7555) & VN_data_in(7555);
  VN1259_in2 <= VN_sign_in(7556) & VN_data_in(7556);
  VN1259_in3 <= VN_sign_in(7557) & VN_data_in(7557);
  VN1259_in4 <= VN_sign_in(7558) & VN_data_in(7558);
  VN1259_in5 <= VN_sign_in(7559) & VN_data_in(7559);
  VN1260_in0 <= VN_sign_in(7560) & VN_data_in(7560);
  VN1260_in1 <= VN_sign_in(7561) & VN_data_in(7561);
  VN1260_in2 <= VN_sign_in(7562) & VN_data_in(7562);
  VN1260_in3 <= VN_sign_in(7563) & VN_data_in(7563);
  VN1260_in4 <= VN_sign_in(7564) & VN_data_in(7564);
  VN1260_in5 <= VN_sign_in(7565) & VN_data_in(7565);
  VN1261_in0 <= VN_sign_in(7566) & VN_data_in(7566);
  VN1261_in1 <= VN_sign_in(7567) & VN_data_in(7567);
  VN1261_in2 <= VN_sign_in(7568) & VN_data_in(7568);
  VN1261_in3 <= VN_sign_in(7569) & VN_data_in(7569);
  VN1261_in4 <= VN_sign_in(7570) & VN_data_in(7570);
  VN1261_in5 <= VN_sign_in(7571) & VN_data_in(7571);
  VN1262_in0 <= VN_sign_in(7572) & VN_data_in(7572);
  VN1262_in1 <= VN_sign_in(7573) & VN_data_in(7573);
  VN1262_in2 <= VN_sign_in(7574) & VN_data_in(7574);
  VN1262_in3 <= VN_sign_in(7575) & VN_data_in(7575);
  VN1262_in4 <= VN_sign_in(7576) & VN_data_in(7576);
  VN1262_in5 <= VN_sign_in(7577) & VN_data_in(7577);
  VN1263_in0 <= VN_sign_in(7578) & VN_data_in(7578);
  VN1263_in1 <= VN_sign_in(7579) & VN_data_in(7579);
  VN1263_in2 <= VN_sign_in(7580) & VN_data_in(7580);
  VN1263_in3 <= VN_sign_in(7581) & VN_data_in(7581);
  VN1263_in4 <= VN_sign_in(7582) & VN_data_in(7582);
  VN1263_in5 <= VN_sign_in(7583) & VN_data_in(7583);
  VN1264_in0 <= VN_sign_in(7584) & VN_data_in(7584);
  VN1264_in1 <= VN_sign_in(7585) & VN_data_in(7585);
  VN1264_in2 <= VN_sign_in(7586) & VN_data_in(7586);
  VN1264_in3 <= VN_sign_in(7587) & VN_data_in(7587);
  VN1264_in4 <= VN_sign_in(7588) & VN_data_in(7588);
  VN1264_in5 <= VN_sign_in(7589) & VN_data_in(7589);
  VN1265_in0 <= VN_sign_in(7590) & VN_data_in(7590);
  VN1265_in1 <= VN_sign_in(7591) & VN_data_in(7591);
  VN1265_in2 <= VN_sign_in(7592) & VN_data_in(7592);
  VN1265_in3 <= VN_sign_in(7593) & VN_data_in(7593);
  VN1265_in4 <= VN_sign_in(7594) & VN_data_in(7594);
  VN1265_in5 <= VN_sign_in(7595) & VN_data_in(7595);
  VN1266_in0 <= VN_sign_in(7596) & VN_data_in(7596);
  VN1266_in1 <= VN_sign_in(7597) & VN_data_in(7597);
  VN1266_in2 <= VN_sign_in(7598) & VN_data_in(7598);
  VN1266_in3 <= VN_sign_in(7599) & VN_data_in(7599);
  VN1266_in4 <= VN_sign_in(7600) & VN_data_in(7600);
  VN1266_in5 <= VN_sign_in(7601) & VN_data_in(7601);
  VN1267_in0 <= VN_sign_in(7602) & VN_data_in(7602);
  VN1267_in1 <= VN_sign_in(7603) & VN_data_in(7603);
  VN1267_in2 <= VN_sign_in(7604) & VN_data_in(7604);
  VN1267_in3 <= VN_sign_in(7605) & VN_data_in(7605);
  VN1267_in4 <= VN_sign_in(7606) & VN_data_in(7606);
  VN1267_in5 <= VN_sign_in(7607) & VN_data_in(7607);
  VN1268_in0 <= VN_sign_in(7608) & VN_data_in(7608);
  VN1268_in1 <= VN_sign_in(7609) & VN_data_in(7609);
  VN1268_in2 <= VN_sign_in(7610) & VN_data_in(7610);
  VN1268_in3 <= VN_sign_in(7611) & VN_data_in(7611);
  VN1268_in4 <= VN_sign_in(7612) & VN_data_in(7612);
  VN1268_in5 <= VN_sign_in(7613) & VN_data_in(7613);
  VN1269_in0 <= VN_sign_in(7614) & VN_data_in(7614);
  VN1269_in1 <= VN_sign_in(7615) & VN_data_in(7615);
  VN1269_in2 <= VN_sign_in(7616) & VN_data_in(7616);
  VN1269_in3 <= VN_sign_in(7617) & VN_data_in(7617);
  VN1269_in4 <= VN_sign_in(7618) & VN_data_in(7618);
  VN1269_in5 <= VN_sign_in(7619) & VN_data_in(7619);
  VN1270_in0 <= VN_sign_in(7620) & VN_data_in(7620);
  VN1270_in1 <= VN_sign_in(7621) & VN_data_in(7621);
  VN1270_in2 <= VN_sign_in(7622) & VN_data_in(7622);
  VN1270_in3 <= VN_sign_in(7623) & VN_data_in(7623);
  VN1270_in4 <= VN_sign_in(7624) & VN_data_in(7624);
  VN1270_in5 <= VN_sign_in(7625) & VN_data_in(7625);
  VN1271_in0 <= VN_sign_in(7626) & VN_data_in(7626);
  VN1271_in1 <= VN_sign_in(7627) & VN_data_in(7627);
  VN1271_in2 <= VN_sign_in(7628) & VN_data_in(7628);
  VN1271_in3 <= VN_sign_in(7629) & VN_data_in(7629);
  VN1271_in4 <= VN_sign_in(7630) & VN_data_in(7630);
  VN1271_in5 <= VN_sign_in(7631) & VN_data_in(7631);
  VN1272_in0 <= VN_sign_in(7632) & VN_data_in(7632);
  VN1272_in1 <= VN_sign_in(7633) & VN_data_in(7633);
  VN1272_in2 <= VN_sign_in(7634) & VN_data_in(7634);
  VN1272_in3 <= VN_sign_in(7635) & VN_data_in(7635);
  VN1272_in4 <= VN_sign_in(7636) & VN_data_in(7636);
  VN1272_in5 <= VN_sign_in(7637) & VN_data_in(7637);
  VN1273_in0 <= VN_sign_in(7638) & VN_data_in(7638);
  VN1273_in1 <= VN_sign_in(7639) & VN_data_in(7639);
  VN1273_in2 <= VN_sign_in(7640) & VN_data_in(7640);
  VN1273_in3 <= VN_sign_in(7641) & VN_data_in(7641);
  VN1273_in4 <= VN_sign_in(7642) & VN_data_in(7642);
  VN1273_in5 <= VN_sign_in(7643) & VN_data_in(7643);
  VN1274_in0 <= VN_sign_in(7644) & VN_data_in(7644);
  VN1274_in1 <= VN_sign_in(7645) & VN_data_in(7645);
  VN1274_in2 <= VN_sign_in(7646) & VN_data_in(7646);
  VN1274_in3 <= VN_sign_in(7647) & VN_data_in(7647);
  VN1274_in4 <= VN_sign_in(7648) & VN_data_in(7648);
  VN1274_in5 <= VN_sign_in(7649) & VN_data_in(7649);
  VN1275_in0 <= VN_sign_in(7650) & VN_data_in(7650);
  VN1275_in1 <= VN_sign_in(7651) & VN_data_in(7651);
  VN1275_in2 <= VN_sign_in(7652) & VN_data_in(7652);
  VN1275_in3 <= VN_sign_in(7653) & VN_data_in(7653);
  VN1275_in4 <= VN_sign_in(7654) & VN_data_in(7654);
  VN1275_in5 <= VN_sign_in(7655) & VN_data_in(7655);
  VN1276_in0 <= VN_sign_in(7656) & VN_data_in(7656);
  VN1276_in1 <= VN_sign_in(7657) & VN_data_in(7657);
  VN1276_in2 <= VN_sign_in(7658) & VN_data_in(7658);
  VN1276_in3 <= VN_sign_in(7659) & VN_data_in(7659);
  VN1276_in4 <= VN_sign_in(7660) & VN_data_in(7660);
  VN1276_in5 <= VN_sign_in(7661) & VN_data_in(7661);
  VN1277_in0 <= VN_sign_in(7662) & VN_data_in(7662);
  VN1277_in1 <= VN_sign_in(7663) & VN_data_in(7663);
  VN1277_in2 <= VN_sign_in(7664) & VN_data_in(7664);
  VN1277_in3 <= VN_sign_in(7665) & VN_data_in(7665);
  VN1277_in4 <= VN_sign_in(7666) & VN_data_in(7666);
  VN1277_in5 <= VN_sign_in(7667) & VN_data_in(7667);
  VN1278_in0 <= VN_sign_in(7668) & VN_data_in(7668);
  VN1278_in1 <= VN_sign_in(7669) & VN_data_in(7669);
  VN1278_in2 <= VN_sign_in(7670) & VN_data_in(7670);
  VN1278_in3 <= VN_sign_in(7671) & VN_data_in(7671);
  VN1278_in4 <= VN_sign_in(7672) & VN_data_in(7672);
  VN1278_in5 <= VN_sign_in(7673) & VN_data_in(7673);
  VN1279_in0 <= VN_sign_in(7674) & VN_data_in(7674);
  VN1279_in1 <= VN_sign_in(7675) & VN_data_in(7675);
  VN1279_in2 <= VN_sign_in(7676) & VN_data_in(7676);
  VN1279_in3 <= VN_sign_in(7677) & VN_data_in(7677);
  VN1279_in4 <= VN_sign_in(7678) & VN_data_in(7678);
  VN1279_in5 <= VN_sign_in(7679) & VN_data_in(7679);
  VN1280_in0 <= VN_sign_in(7680) & VN_data_in(7680);
  VN1280_in1 <= VN_sign_in(7681) & VN_data_in(7681);
  VN1280_in2 <= VN_sign_in(7682) & VN_data_in(7682);
  VN1280_in3 <= VN_sign_in(7683) & VN_data_in(7683);
  VN1280_in4 <= VN_sign_in(7684) & VN_data_in(7684);
  VN1280_in5 <= VN_sign_in(7685) & VN_data_in(7685);
  VN1281_in0 <= VN_sign_in(7686) & VN_data_in(7686);
  VN1281_in1 <= VN_sign_in(7687) & VN_data_in(7687);
  VN1281_in2 <= VN_sign_in(7688) & VN_data_in(7688);
  VN1281_in3 <= VN_sign_in(7689) & VN_data_in(7689);
  VN1281_in4 <= VN_sign_in(7690) & VN_data_in(7690);
  VN1281_in5 <= VN_sign_in(7691) & VN_data_in(7691);
  VN1282_in0 <= VN_sign_in(7692) & VN_data_in(7692);
  VN1282_in1 <= VN_sign_in(7693) & VN_data_in(7693);
  VN1282_in2 <= VN_sign_in(7694) & VN_data_in(7694);
  VN1282_in3 <= VN_sign_in(7695) & VN_data_in(7695);
  VN1282_in4 <= VN_sign_in(7696) & VN_data_in(7696);
  VN1282_in5 <= VN_sign_in(7697) & VN_data_in(7697);
  VN1283_in0 <= VN_sign_in(7698) & VN_data_in(7698);
  VN1283_in1 <= VN_sign_in(7699) & VN_data_in(7699);
  VN1283_in2 <= VN_sign_in(7700) & VN_data_in(7700);
  VN1283_in3 <= VN_sign_in(7701) & VN_data_in(7701);
  VN1283_in4 <= VN_sign_in(7702) & VN_data_in(7702);
  VN1283_in5 <= VN_sign_in(7703) & VN_data_in(7703);
  VN1284_in0 <= VN_sign_in(7704) & VN_data_in(7704);
  VN1284_in1 <= VN_sign_in(7705) & VN_data_in(7705);
  VN1284_in2 <= VN_sign_in(7706) & VN_data_in(7706);
  VN1284_in3 <= VN_sign_in(7707) & VN_data_in(7707);
  VN1284_in4 <= VN_sign_in(7708) & VN_data_in(7708);
  VN1284_in5 <= VN_sign_in(7709) & VN_data_in(7709);
  VN1285_in0 <= VN_sign_in(7710) & VN_data_in(7710);
  VN1285_in1 <= VN_sign_in(7711) & VN_data_in(7711);
  VN1285_in2 <= VN_sign_in(7712) & VN_data_in(7712);
  VN1285_in3 <= VN_sign_in(7713) & VN_data_in(7713);
  VN1285_in4 <= VN_sign_in(7714) & VN_data_in(7714);
  VN1285_in5 <= VN_sign_in(7715) & VN_data_in(7715);
  VN1286_in0 <= VN_sign_in(7716) & VN_data_in(7716);
  VN1286_in1 <= VN_sign_in(7717) & VN_data_in(7717);
  VN1286_in2 <= VN_sign_in(7718) & VN_data_in(7718);
  VN1286_in3 <= VN_sign_in(7719) & VN_data_in(7719);
  VN1286_in4 <= VN_sign_in(7720) & VN_data_in(7720);
  VN1286_in5 <= VN_sign_in(7721) & VN_data_in(7721);
  VN1287_in0 <= VN_sign_in(7722) & VN_data_in(7722);
  VN1287_in1 <= VN_sign_in(7723) & VN_data_in(7723);
  VN1287_in2 <= VN_sign_in(7724) & VN_data_in(7724);
  VN1287_in3 <= VN_sign_in(7725) & VN_data_in(7725);
  VN1287_in4 <= VN_sign_in(7726) & VN_data_in(7726);
  VN1287_in5 <= VN_sign_in(7727) & VN_data_in(7727);
  VN1288_in0 <= VN_sign_in(7728) & VN_data_in(7728);
  VN1288_in1 <= VN_sign_in(7729) & VN_data_in(7729);
  VN1288_in2 <= VN_sign_in(7730) & VN_data_in(7730);
  VN1288_in3 <= VN_sign_in(7731) & VN_data_in(7731);
  VN1288_in4 <= VN_sign_in(7732) & VN_data_in(7732);
  VN1288_in5 <= VN_sign_in(7733) & VN_data_in(7733);
  VN1289_in0 <= VN_sign_in(7734) & VN_data_in(7734);
  VN1289_in1 <= VN_sign_in(7735) & VN_data_in(7735);
  VN1289_in2 <= VN_sign_in(7736) & VN_data_in(7736);
  VN1289_in3 <= VN_sign_in(7737) & VN_data_in(7737);
  VN1289_in4 <= VN_sign_in(7738) & VN_data_in(7738);
  VN1289_in5 <= VN_sign_in(7739) & VN_data_in(7739);
  VN1290_in0 <= VN_sign_in(7740) & VN_data_in(7740);
  VN1290_in1 <= VN_sign_in(7741) & VN_data_in(7741);
  VN1290_in2 <= VN_sign_in(7742) & VN_data_in(7742);
  VN1290_in3 <= VN_sign_in(7743) & VN_data_in(7743);
  VN1290_in4 <= VN_sign_in(7744) & VN_data_in(7744);
  VN1290_in5 <= VN_sign_in(7745) & VN_data_in(7745);
  VN1291_in0 <= VN_sign_in(7746) & VN_data_in(7746);
  VN1291_in1 <= VN_sign_in(7747) & VN_data_in(7747);
  VN1291_in2 <= VN_sign_in(7748) & VN_data_in(7748);
  VN1291_in3 <= VN_sign_in(7749) & VN_data_in(7749);
  VN1291_in4 <= VN_sign_in(7750) & VN_data_in(7750);
  VN1291_in5 <= VN_sign_in(7751) & VN_data_in(7751);
  VN1292_in0 <= VN_sign_in(7752) & VN_data_in(7752);
  VN1292_in1 <= VN_sign_in(7753) & VN_data_in(7753);
  VN1292_in2 <= VN_sign_in(7754) & VN_data_in(7754);
  VN1292_in3 <= VN_sign_in(7755) & VN_data_in(7755);
  VN1292_in4 <= VN_sign_in(7756) & VN_data_in(7756);
  VN1292_in5 <= VN_sign_in(7757) & VN_data_in(7757);
  VN1293_in0 <= VN_sign_in(7758) & VN_data_in(7758);
  VN1293_in1 <= VN_sign_in(7759) & VN_data_in(7759);
  VN1293_in2 <= VN_sign_in(7760) & VN_data_in(7760);
  VN1293_in3 <= VN_sign_in(7761) & VN_data_in(7761);
  VN1293_in4 <= VN_sign_in(7762) & VN_data_in(7762);
  VN1293_in5 <= VN_sign_in(7763) & VN_data_in(7763);
  VN1294_in0 <= VN_sign_in(7764) & VN_data_in(7764);
  VN1294_in1 <= VN_sign_in(7765) & VN_data_in(7765);
  VN1294_in2 <= VN_sign_in(7766) & VN_data_in(7766);
  VN1294_in3 <= VN_sign_in(7767) & VN_data_in(7767);
  VN1294_in4 <= VN_sign_in(7768) & VN_data_in(7768);
  VN1294_in5 <= VN_sign_in(7769) & VN_data_in(7769);
  VN1295_in0 <= VN_sign_in(7770) & VN_data_in(7770);
  VN1295_in1 <= VN_sign_in(7771) & VN_data_in(7771);
  VN1295_in2 <= VN_sign_in(7772) & VN_data_in(7772);
  VN1295_in3 <= VN_sign_in(7773) & VN_data_in(7773);
  VN1295_in4 <= VN_sign_in(7774) & VN_data_in(7774);
  VN1295_in5 <= VN_sign_in(7775) & VN_data_in(7775);
  VN1296_in0 <= VN_sign_in(7776) & VN_data_in(7776);
  VN1296_in1 <= VN_sign_in(7777) & VN_data_in(7777);
  VN1296_in2 <= VN_sign_in(7778) & VN_data_in(7778);
  VN1296_in3 <= VN_sign_in(7779) & VN_data_in(7779);
  VN1296_in4 <= VN_sign_in(7780) & VN_data_in(7780);
  VN1296_in5 <= VN_sign_in(7781) & VN_data_in(7781);
  VN1297_in0 <= VN_sign_in(7782) & VN_data_in(7782);
  VN1297_in1 <= VN_sign_in(7783) & VN_data_in(7783);
  VN1297_in2 <= VN_sign_in(7784) & VN_data_in(7784);
  VN1297_in3 <= VN_sign_in(7785) & VN_data_in(7785);
  VN1297_in4 <= VN_sign_in(7786) & VN_data_in(7786);
  VN1297_in5 <= VN_sign_in(7787) & VN_data_in(7787);
  VN1298_in0 <= VN_sign_in(7788) & VN_data_in(7788);
  VN1298_in1 <= VN_sign_in(7789) & VN_data_in(7789);
  VN1298_in2 <= VN_sign_in(7790) & VN_data_in(7790);
  VN1298_in3 <= VN_sign_in(7791) & VN_data_in(7791);
  VN1298_in4 <= VN_sign_in(7792) & VN_data_in(7792);
  VN1298_in5 <= VN_sign_in(7793) & VN_data_in(7793);
  VN1299_in0 <= VN_sign_in(7794) & VN_data_in(7794);
  VN1299_in1 <= VN_sign_in(7795) & VN_data_in(7795);
  VN1299_in2 <= VN_sign_in(7796) & VN_data_in(7796);
  VN1299_in3 <= VN_sign_in(7797) & VN_data_in(7797);
  VN1299_in4 <= VN_sign_in(7798) & VN_data_in(7798);
  VN1299_in5 <= VN_sign_in(7799) & VN_data_in(7799);
  VN1300_in0 <= VN_sign_in(7800) & VN_data_in(7800);
  VN1300_in1 <= VN_sign_in(7801) & VN_data_in(7801);
  VN1300_in2 <= VN_sign_in(7802) & VN_data_in(7802);
  VN1300_in3 <= VN_sign_in(7803) & VN_data_in(7803);
  VN1300_in4 <= VN_sign_in(7804) & VN_data_in(7804);
  VN1300_in5 <= VN_sign_in(7805) & VN_data_in(7805);
  VN1301_in0 <= VN_sign_in(7806) & VN_data_in(7806);
  VN1301_in1 <= VN_sign_in(7807) & VN_data_in(7807);
  VN1301_in2 <= VN_sign_in(7808) & VN_data_in(7808);
  VN1301_in3 <= VN_sign_in(7809) & VN_data_in(7809);
  VN1301_in4 <= VN_sign_in(7810) & VN_data_in(7810);
  VN1301_in5 <= VN_sign_in(7811) & VN_data_in(7811);
  VN1302_in0 <= VN_sign_in(7812) & VN_data_in(7812);
  VN1302_in1 <= VN_sign_in(7813) & VN_data_in(7813);
  VN1302_in2 <= VN_sign_in(7814) & VN_data_in(7814);
  VN1302_in3 <= VN_sign_in(7815) & VN_data_in(7815);
  VN1302_in4 <= VN_sign_in(7816) & VN_data_in(7816);
  VN1302_in5 <= VN_sign_in(7817) & VN_data_in(7817);
  VN1303_in0 <= VN_sign_in(7818) & VN_data_in(7818);
  VN1303_in1 <= VN_sign_in(7819) & VN_data_in(7819);
  VN1303_in2 <= VN_sign_in(7820) & VN_data_in(7820);
  VN1303_in3 <= VN_sign_in(7821) & VN_data_in(7821);
  VN1303_in4 <= VN_sign_in(7822) & VN_data_in(7822);
  VN1303_in5 <= VN_sign_in(7823) & VN_data_in(7823);
  VN1304_in0 <= VN_sign_in(7824) & VN_data_in(7824);
  VN1304_in1 <= VN_sign_in(7825) & VN_data_in(7825);
  VN1304_in2 <= VN_sign_in(7826) & VN_data_in(7826);
  VN1304_in3 <= VN_sign_in(7827) & VN_data_in(7827);
  VN1304_in4 <= VN_sign_in(7828) & VN_data_in(7828);
  VN1304_in5 <= VN_sign_in(7829) & VN_data_in(7829);
  VN1305_in0 <= VN_sign_in(7830) & VN_data_in(7830);
  VN1305_in1 <= VN_sign_in(7831) & VN_data_in(7831);
  VN1305_in2 <= VN_sign_in(7832) & VN_data_in(7832);
  VN1305_in3 <= VN_sign_in(7833) & VN_data_in(7833);
  VN1305_in4 <= VN_sign_in(7834) & VN_data_in(7834);
  VN1305_in5 <= VN_sign_in(7835) & VN_data_in(7835);
  VN1306_in0 <= VN_sign_in(7836) & VN_data_in(7836);
  VN1306_in1 <= VN_sign_in(7837) & VN_data_in(7837);
  VN1306_in2 <= VN_sign_in(7838) & VN_data_in(7838);
  VN1306_in3 <= VN_sign_in(7839) & VN_data_in(7839);
  VN1306_in4 <= VN_sign_in(7840) & VN_data_in(7840);
  VN1306_in5 <= VN_sign_in(7841) & VN_data_in(7841);
  VN1307_in0 <= VN_sign_in(7842) & VN_data_in(7842);
  VN1307_in1 <= VN_sign_in(7843) & VN_data_in(7843);
  VN1307_in2 <= VN_sign_in(7844) & VN_data_in(7844);
  VN1307_in3 <= VN_sign_in(7845) & VN_data_in(7845);
  VN1307_in4 <= VN_sign_in(7846) & VN_data_in(7846);
  VN1307_in5 <= VN_sign_in(7847) & VN_data_in(7847);
  VN1308_in0 <= VN_sign_in(7848) & VN_data_in(7848);
  VN1308_in1 <= VN_sign_in(7849) & VN_data_in(7849);
  VN1308_in2 <= VN_sign_in(7850) & VN_data_in(7850);
  VN1308_in3 <= VN_sign_in(7851) & VN_data_in(7851);
  VN1308_in4 <= VN_sign_in(7852) & VN_data_in(7852);
  VN1308_in5 <= VN_sign_in(7853) & VN_data_in(7853);
  VN1309_in0 <= VN_sign_in(7854) & VN_data_in(7854);
  VN1309_in1 <= VN_sign_in(7855) & VN_data_in(7855);
  VN1309_in2 <= VN_sign_in(7856) & VN_data_in(7856);
  VN1309_in3 <= VN_sign_in(7857) & VN_data_in(7857);
  VN1309_in4 <= VN_sign_in(7858) & VN_data_in(7858);
  VN1309_in5 <= VN_sign_in(7859) & VN_data_in(7859);
  VN1310_in0 <= VN_sign_in(7860) & VN_data_in(7860);
  VN1310_in1 <= VN_sign_in(7861) & VN_data_in(7861);
  VN1310_in2 <= VN_sign_in(7862) & VN_data_in(7862);
  VN1310_in3 <= VN_sign_in(7863) & VN_data_in(7863);
  VN1310_in4 <= VN_sign_in(7864) & VN_data_in(7864);
  VN1310_in5 <= VN_sign_in(7865) & VN_data_in(7865);
  VN1311_in0 <= VN_sign_in(7866) & VN_data_in(7866);
  VN1311_in1 <= VN_sign_in(7867) & VN_data_in(7867);
  VN1311_in2 <= VN_sign_in(7868) & VN_data_in(7868);
  VN1311_in3 <= VN_sign_in(7869) & VN_data_in(7869);
  VN1311_in4 <= VN_sign_in(7870) & VN_data_in(7870);
  VN1311_in5 <= VN_sign_in(7871) & VN_data_in(7871);
  VN1312_in0 <= VN_sign_in(7872) & VN_data_in(7872);
  VN1312_in1 <= VN_sign_in(7873) & VN_data_in(7873);
  VN1312_in2 <= VN_sign_in(7874) & VN_data_in(7874);
  VN1312_in3 <= VN_sign_in(7875) & VN_data_in(7875);
  VN1312_in4 <= VN_sign_in(7876) & VN_data_in(7876);
  VN1312_in5 <= VN_sign_in(7877) & VN_data_in(7877);
  VN1313_in0 <= VN_sign_in(7878) & VN_data_in(7878);
  VN1313_in1 <= VN_sign_in(7879) & VN_data_in(7879);
  VN1313_in2 <= VN_sign_in(7880) & VN_data_in(7880);
  VN1313_in3 <= VN_sign_in(7881) & VN_data_in(7881);
  VN1313_in4 <= VN_sign_in(7882) & VN_data_in(7882);
  VN1313_in5 <= VN_sign_in(7883) & VN_data_in(7883);
  VN1314_in0 <= VN_sign_in(7884) & VN_data_in(7884);
  VN1314_in1 <= VN_sign_in(7885) & VN_data_in(7885);
  VN1314_in2 <= VN_sign_in(7886) & VN_data_in(7886);
  VN1314_in3 <= VN_sign_in(7887) & VN_data_in(7887);
  VN1314_in4 <= VN_sign_in(7888) & VN_data_in(7888);
  VN1314_in5 <= VN_sign_in(7889) & VN_data_in(7889);
  VN1315_in0 <= VN_sign_in(7890) & VN_data_in(7890);
  VN1315_in1 <= VN_sign_in(7891) & VN_data_in(7891);
  VN1315_in2 <= VN_sign_in(7892) & VN_data_in(7892);
  VN1315_in3 <= VN_sign_in(7893) & VN_data_in(7893);
  VN1315_in4 <= VN_sign_in(7894) & VN_data_in(7894);
  VN1315_in5 <= VN_sign_in(7895) & VN_data_in(7895);
  VN1316_in0 <= VN_sign_in(7896) & VN_data_in(7896);
  VN1316_in1 <= VN_sign_in(7897) & VN_data_in(7897);
  VN1316_in2 <= VN_sign_in(7898) & VN_data_in(7898);
  VN1316_in3 <= VN_sign_in(7899) & VN_data_in(7899);
  VN1316_in4 <= VN_sign_in(7900) & VN_data_in(7900);
  VN1316_in5 <= VN_sign_in(7901) & VN_data_in(7901);
  VN1317_in0 <= VN_sign_in(7902) & VN_data_in(7902);
  VN1317_in1 <= VN_sign_in(7903) & VN_data_in(7903);
  VN1317_in2 <= VN_sign_in(7904) & VN_data_in(7904);
  VN1317_in3 <= VN_sign_in(7905) & VN_data_in(7905);
  VN1317_in4 <= VN_sign_in(7906) & VN_data_in(7906);
  VN1317_in5 <= VN_sign_in(7907) & VN_data_in(7907);
  VN1318_in0 <= VN_sign_in(7908) & VN_data_in(7908);
  VN1318_in1 <= VN_sign_in(7909) & VN_data_in(7909);
  VN1318_in2 <= VN_sign_in(7910) & VN_data_in(7910);
  VN1318_in3 <= VN_sign_in(7911) & VN_data_in(7911);
  VN1318_in4 <= VN_sign_in(7912) & VN_data_in(7912);
  VN1318_in5 <= VN_sign_in(7913) & VN_data_in(7913);
  VN1319_in0 <= VN_sign_in(7914) & VN_data_in(7914);
  VN1319_in1 <= VN_sign_in(7915) & VN_data_in(7915);
  VN1319_in2 <= VN_sign_in(7916) & VN_data_in(7916);
  VN1319_in3 <= VN_sign_in(7917) & VN_data_in(7917);
  VN1319_in4 <= VN_sign_in(7918) & VN_data_in(7918);
  VN1319_in5 <= VN_sign_in(7919) & VN_data_in(7919);
  VN1320_in0 <= VN_sign_in(7920) & VN_data_in(7920);
  VN1320_in1 <= VN_sign_in(7921) & VN_data_in(7921);
  VN1320_in2 <= VN_sign_in(7922) & VN_data_in(7922);
  VN1320_in3 <= VN_sign_in(7923) & VN_data_in(7923);
  VN1320_in4 <= VN_sign_in(7924) & VN_data_in(7924);
  VN1320_in5 <= VN_sign_in(7925) & VN_data_in(7925);
  VN1321_in0 <= VN_sign_in(7926) & VN_data_in(7926);
  VN1321_in1 <= VN_sign_in(7927) & VN_data_in(7927);
  VN1321_in2 <= VN_sign_in(7928) & VN_data_in(7928);
  VN1321_in3 <= VN_sign_in(7929) & VN_data_in(7929);
  VN1321_in4 <= VN_sign_in(7930) & VN_data_in(7930);
  VN1321_in5 <= VN_sign_in(7931) & VN_data_in(7931);
  VN1322_in0 <= VN_sign_in(7932) & VN_data_in(7932);
  VN1322_in1 <= VN_sign_in(7933) & VN_data_in(7933);
  VN1322_in2 <= VN_sign_in(7934) & VN_data_in(7934);
  VN1322_in3 <= VN_sign_in(7935) & VN_data_in(7935);
  VN1322_in4 <= VN_sign_in(7936) & VN_data_in(7936);
  VN1322_in5 <= VN_sign_in(7937) & VN_data_in(7937);
  VN1323_in0 <= VN_sign_in(7938) & VN_data_in(7938);
  VN1323_in1 <= VN_sign_in(7939) & VN_data_in(7939);
  VN1323_in2 <= VN_sign_in(7940) & VN_data_in(7940);
  VN1323_in3 <= VN_sign_in(7941) & VN_data_in(7941);
  VN1323_in4 <= VN_sign_in(7942) & VN_data_in(7942);
  VN1323_in5 <= VN_sign_in(7943) & VN_data_in(7943);
  VN1324_in0 <= VN_sign_in(7944) & VN_data_in(7944);
  VN1324_in1 <= VN_sign_in(7945) & VN_data_in(7945);
  VN1324_in2 <= VN_sign_in(7946) & VN_data_in(7946);
  VN1324_in3 <= VN_sign_in(7947) & VN_data_in(7947);
  VN1324_in4 <= VN_sign_in(7948) & VN_data_in(7948);
  VN1324_in5 <= VN_sign_in(7949) & VN_data_in(7949);
  VN1325_in0 <= VN_sign_in(7950) & VN_data_in(7950);
  VN1325_in1 <= VN_sign_in(7951) & VN_data_in(7951);
  VN1325_in2 <= VN_sign_in(7952) & VN_data_in(7952);
  VN1325_in3 <= VN_sign_in(7953) & VN_data_in(7953);
  VN1325_in4 <= VN_sign_in(7954) & VN_data_in(7954);
  VN1325_in5 <= VN_sign_in(7955) & VN_data_in(7955);
  VN1326_in0 <= VN_sign_in(7956) & VN_data_in(7956);
  VN1326_in1 <= VN_sign_in(7957) & VN_data_in(7957);
  VN1326_in2 <= VN_sign_in(7958) & VN_data_in(7958);
  VN1326_in3 <= VN_sign_in(7959) & VN_data_in(7959);
  VN1326_in4 <= VN_sign_in(7960) & VN_data_in(7960);
  VN1326_in5 <= VN_sign_in(7961) & VN_data_in(7961);
  VN1327_in0 <= VN_sign_in(7962) & VN_data_in(7962);
  VN1327_in1 <= VN_sign_in(7963) & VN_data_in(7963);
  VN1327_in2 <= VN_sign_in(7964) & VN_data_in(7964);
  VN1327_in3 <= VN_sign_in(7965) & VN_data_in(7965);
  VN1327_in4 <= VN_sign_in(7966) & VN_data_in(7966);
  VN1327_in5 <= VN_sign_in(7967) & VN_data_in(7967);
  VN1328_in0 <= VN_sign_in(7968) & VN_data_in(7968);
  VN1328_in1 <= VN_sign_in(7969) & VN_data_in(7969);
  VN1328_in2 <= VN_sign_in(7970) & VN_data_in(7970);
  VN1328_in3 <= VN_sign_in(7971) & VN_data_in(7971);
  VN1328_in4 <= VN_sign_in(7972) & VN_data_in(7972);
  VN1328_in5 <= VN_sign_in(7973) & VN_data_in(7973);
  VN1329_in0 <= VN_sign_in(7974) & VN_data_in(7974);
  VN1329_in1 <= VN_sign_in(7975) & VN_data_in(7975);
  VN1329_in2 <= VN_sign_in(7976) & VN_data_in(7976);
  VN1329_in3 <= VN_sign_in(7977) & VN_data_in(7977);
  VN1329_in4 <= VN_sign_in(7978) & VN_data_in(7978);
  VN1329_in5 <= VN_sign_in(7979) & VN_data_in(7979);
  VN1330_in0 <= VN_sign_in(7980) & VN_data_in(7980);
  VN1330_in1 <= VN_sign_in(7981) & VN_data_in(7981);
  VN1330_in2 <= VN_sign_in(7982) & VN_data_in(7982);
  VN1330_in3 <= VN_sign_in(7983) & VN_data_in(7983);
  VN1330_in4 <= VN_sign_in(7984) & VN_data_in(7984);
  VN1330_in5 <= VN_sign_in(7985) & VN_data_in(7985);
  VN1331_in0 <= VN_sign_in(7986) & VN_data_in(7986);
  VN1331_in1 <= VN_sign_in(7987) & VN_data_in(7987);
  VN1331_in2 <= VN_sign_in(7988) & VN_data_in(7988);
  VN1331_in3 <= VN_sign_in(7989) & VN_data_in(7989);
  VN1331_in4 <= VN_sign_in(7990) & VN_data_in(7990);
  VN1331_in5 <= VN_sign_in(7991) & VN_data_in(7991);
  VN1332_in0 <= VN_sign_in(7992) & VN_data_in(7992);
  VN1332_in1 <= VN_sign_in(7993) & VN_data_in(7993);
  VN1332_in2 <= VN_sign_in(7994) & VN_data_in(7994);
  VN1332_in3 <= VN_sign_in(7995) & VN_data_in(7995);
  VN1332_in4 <= VN_sign_in(7996) & VN_data_in(7996);
  VN1332_in5 <= VN_sign_in(7997) & VN_data_in(7997);
  VN1333_in0 <= VN_sign_in(7998) & VN_data_in(7998);
  VN1333_in1 <= VN_sign_in(7999) & VN_data_in(7999);
  VN1333_in2 <= VN_sign_in(8000) & VN_data_in(8000);
  VN1333_in3 <= VN_sign_in(8001) & VN_data_in(8001);
  VN1333_in4 <= VN_sign_in(8002) & VN_data_in(8002);
  VN1333_in5 <= VN_sign_in(8003) & VN_data_in(8003);
  VN1334_in0 <= VN_sign_in(8004) & VN_data_in(8004);
  VN1334_in1 <= VN_sign_in(8005) & VN_data_in(8005);
  VN1334_in2 <= VN_sign_in(8006) & VN_data_in(8006);
  VN1334_in3 <= VN_sign_in(8007) & VN_data_in(8007);
  VN1334_in4 <= VN_sign_in(8008) & VN_data_in(8008);
  VN1334_in5 <= VN_sign_in(8009) & VN_data_in(8009);
  VN1335_in0 <= VN_sign_in(8010) & VN_data_in(8010);
  VN1335_in1 <= VN_sign_in(8011) & VN_data_in(8011);
  VN1335_in2 <= VN_sign_in(8012) & VN_data_in(8012);
  VN1335_in3 <= VN_sign_in(8013) & VN_data_in(8013);
  VN1335_in4 <= VN_sign_in(8014) & VN_data_in(8014);
  VN1335_in5 <= VN_sign_in(8015) & VN_data_in(8015);
  VN1336_in0 <= VN_sign_in(8016) & VN_data_in(8016);
  VN1336_in1 <= VN_sign_in(8017) & VN_data_in(8017);
  VN1336_in2 <= VN_sign_in(8018) & VN_data_in(8018);
  VN1336_in3 <= VN_sign_in(8019) & VN_data_in(8019);
  VN1336_in4 <= VN_sign_in(8020) & VN_data_in(8020);
  VN1336_in5 <= VN_sign_in(8021) & VN_data_in(8021);
  VN1337_in0 <= VN_sign_in(8022) & VN_data_in(8022);
  VN1337_in1 <= VN_sign_in(8023) & VN_data_in(8023);
  VN1337_in2 <= VN_sign_in(8024) & VN_data_in(8024);
  VN1337_in3 <= VN_sign_in(8025) & VN_data_in(8025);
  VN1337_in4 <= VN_sign_in(8026) & VN_data_in(8026);
  VN1337_in5 <= VN_sign_in(8027) & VN_data_in(8027);
  VN1338_in0 <= VN_sign_in(8028) & VN_data_in(8028);
  VN1338_in1 <= VN_sign_in(8029) & VN_data_in(8029);
  VN1338_in2 <= VN_sign_in(8030) & VN_data_in(8030);
  VN1338_in3 <= VN_sign_in(8031) & VN_data_in(8031);
  VN1338_in4 <= VN_sign_in(8032) & VN_data_in(8032);
  VN1338_in5 <= VN_sign_in(8033) & VN_data_in(8033);
  VN1339_in0 <= VN_sign_in(8034) & VN_data_in(8034);
  VN1339_in1 <= VN_sign_in(8035) & VN_data_in(8035);
  VN1339_in2 <= VN_sign_in(8036) & VN_data_in(8036);
  VN1339_in3 <= VN_sign_in(8037) & VN_data_in(8037);
  VN1339_in4 <= VN_sign_in(8038) & VN_data_in(8038);
  VN1339_in5 <= VN_sign_in(8039) & VN_data_in(8039);
  VN1340_in0 <= VN_sign_in(8040) & VN_data_in(8040);
  VN1340_in1 <= VN_sign_in(8041) & VN_data_in(8041);
  VN1340_in2 <= VN_sign_in(8042) & VN_data_in(8042);
  VN1340_in3 <= VN_sign_in(8043) & VN_data_in(8043);
  VN1340_in4 <= VN_sign_in(8044) & VN_data_in(8044);
  VN1340_in5 <= VN_sign_in(8045) & VN_data_in(8045);
  VN1341_in0 <= VN_sign_in(8046) & VN_data_in(8046);
  VN1341_in1 <= VN_sign_in(8047) & VN_data_in(8047);
  VN1341_in2 <= VN_sign_in(8048) & VN_data_in(8048);
  VN1341_in3 <= VN_sign_in(8049) & VN_data_in(8049);
  VN1341_in4 <= VN_sign_in(8050) & VN_data_in(8050);
  VN1341_in5 <= VN_sign_in(8051) & VN_data_in(8051);
  VN1342_in0 <= VN_sign_in(8052) & VN_data_in(8052);
  VN1342_in1 <= VN_sign_in(8053) & VN_data_in(8053);
  VN1342_in2 <= VN_sign_in(8054) & VN_data_in(8054);
  VN1342_in3 <= VN_sign_in(8055) & VN_data_in(8055);
  VN1342_in4 <= VN_sign_in(8056) & VN_data_in(8056);
  VN1342_in5 <= VN_sign_in(8057) & VN_data_in(8057);
  VN1343_in0 <= VN_sign_in(8058) & VN_data_in(8058);
  VN1343_in1 <= VN_sign_in(8059) & VN_data_in(8059);
  VN1343_in2 <= VN_sign_in(8060) & VN_data_in(8060);
  VN1343_in3 <= VN_sign_in(8061) & VN_data_in(8061);
  VN1343_in4 <= VN_sign_in(8062) & VN_data_in(8062);
  VN1343_in5 <= VN_sign_in(8063) & VN_data_in(8063);
  VN1344_in0 <= VN_sign_in(8064) & VN_data_in(8064);
  VN1344_in1 <= VN_sign_in(8065) & VN_data_in(8065);
  VN1344_in2 <= VN_sign_in(8066) & VN_data_in(8066);
  VN1344_in3 <= VN_sign_in(8067) & VN_data_in(8067);
  VN1344_in4 <= VN_sign_in(8068) & VN_data_in(8068);
  VN1344_in5 <= VN_sign_in(8069) & VN_data_in(8069);
  VN1345_in0 <= VN_sign_in(8070) & VN_data_in(8070);
  VN1345_in1 <= VN_sign_in(8071) & VN_data_in(8071);
  VN1345_in2 <= VN_sign_in(8072) & VN_data_in(8072);
  VN1345_in3 <= VN_sign_in(8073) & VN_data_in(8073);
  VN1345_in4 <= VN_sign_in(8074) & VN_data_in(8074);
  VN1345_in5 <= VN_sign_in(8075) & VN_data_in(8075);
  VN1346_in0 <= VN_sign_in(8076) & VN_data_in(8076);
  VN1346_in1 <= VN_sign_in(8077) & VN_data_in(8077);
  VN1346_in2 <= VN_sign_in(8078) & VN_data_in(8078);
  VN1346_in3 <= VN_sign_in(8079) & VN_data_in(8079);
  VN1346_in4 <= VN_sign_in(8080) & VN_data_in(8080);
  VN1346_in5 <= VN_sign_in(8081) & VN_data_in(8081);
  VN1347_in0 <= VN_sign_in(8082) & VN_data_in(8082);
  VN1347_in1 <= VN_sign_in(8083) & VN_data_in(8083);
  VN1347_in2 <= VN_sign_in(8084) & VN_data_in(8084);
  VN1347_in3 <= VN_sign_in(8085) & VN_data_in(8085);
  VN1347_in4 <= VN_sign_in(8086) & VN_data_in(8086);
  VN1347_in5 <= VN_sign_in(8087) & VN_data_in(8087);
  VN1348_in0 <= VN_sign_in(8088) & VN_data_in(8088);
  VN1348_in1 <= VN_sign_in(8089) & VN_data_in(8089);
  VN1348_in2 <= VN_sign_in(8090) & VN_data_in(8090);
  VN1348_in3 <= VN_sign_in(8091) & VN_data_in(8091);
  VN1348_in4 <= VN_sign_in(8092) & VN_data_in(8092);
  VN1348_in5 <= VN_sign_in(8093) & VN_data_in(8093);
  VN1349_in0 <= VN_sign_in(8094) & VN_data_in(8094);
  VN1349_in1 <= VN_sign_in(8095) & VN_data_in(8095);
  VN1349_in2 <= VN_sign_in(8096) & VN_data_in(8096);
  VN1349_in3 <= VN_sign_in(8097) & VN_data_in(8097);
  VN1349_in4 <= VN_sign_in(8098) & VN_data_in(8098);
  VN1349_in5 <= VN_sign_in(8099) & VN_data_in(8099);
  VN1350_in0 <= VN_sign_in(8100) & VN_data_in(8100);
  VN1350_in1 <= VN_sign_in(8101) & VN_data_in(8101);
  VN1350_in2 <= VN_sign_in(8102) & VN_data_in(8102);
  VN1350_in3 <= VN_sign_in(8103) & VN_data_in(8103);
  VN1350_in4 <= VN_sign_in(8104) & VN_data_in(8104);
  VN1350_in5 <= VN_sign_in(8105) & VN_data_in(8105);
  VN1351_in0 <= VN_sign_in(8106) & VN_data_in(8106);
  VN1351_in1 <= VN_sign_in(8107) & VN_data_in(8107);
  VN1351_in2 <= VN_sign_in(8108) & VN_data_in(8108);
  VN1351_in3 <= VN_sign_in(8109) & VN_data_in(8109);
  VN1351_in4 <= VN_sign_in(8110) & VN_data_in(8110);
  VN1351_in5 <= VN_sign_in(8111) & VN_data_in(8111);
  VN1352_in0 <= VN_sign_in(8112) & VN_data_in(8112);
  VN1352_in1 <= VN_sign_in(8113) & VN_data_in(8113);
  VN1352_in2 <= VN_sign_in(8114) & VN_data_in(8114);
  VN1352_in3 <= VN_sign_in(8115) & VN_data_in(8115);
  VN1352_in4 <= VN_sign_in(8116) & VN_data_in(8116);
  VN1352_in5 <= VN_sign_in(8117) & VN_data_in(8117);
  VN1353_in0 <= VN_sign_in(8118) & VN_data_in(8118);
  VN1353_in1 <= VN_sign_in(8119) & VN_data_in(8119);
  VN1353_in2 <= VN_sign_in(8120) & VN_data_in(8120);
  VN1353_in3 <= VN_sign_in(8121) & VN_data_in(8121);
  VN1353_in4 <= VN_sign_in(8122) & VN_data_in(8122);
  VN1353_in5 <= VN_sign_in(8123) & VN_data_in(8123);
  VN1354_in0 <= VN_sign_in(8124) & VN_data_in(8124);
  VN1354_in1 <= VN_sign_in(8125) & VN_data_in(8125);
  VN1354_in2 <= VN_sign_in(8126) & VN_data_in(8126);
  VN1354_in3 <= VN_sign_in(8127) & VN_data_in(8127);
  VN1354_in4 <= VN_sign_in(8128) & VN_data_in(8128);
  VN1354_in5 <= VN_sign_in(8129) & VN_data_in(8129);
  VN1355_in0 <= VN_sign_in(8130) & VN_data_in(8130);
  VN1355_in1 <= VN_sign_in(8131) & VN_data_in(8131);
  VN1355_in2 <= VN_sign_in(8132) & VN_data_in(8132);
  VN1355_in3 <= VN_sign_in(8133) & VN_data_in(8133);
  VN1355_in4 <= VN_sign_in(8134) & VN_data_in(8134);
  VN1355_in5 <= VN_sign_in(8135) & VN_data_in(8135);
  VN1356_in0 <= VN_sign_in(8136) & VN_data_in(8136);
  VN1356_in1 <= VN_sign_in(8137) & VN_data_in(8137);
  VN1356_in2 <= VN_sign_in(8138) & VN_data_in(8138);
  VN1356_in3 <= VN_sign_in(8139) & VN_data_in(8139);
  VN1356_in4 <= VN_sign_in(8140) & VN_data_in(8140);
  VN1356_in5 <= VN_sign_in(8141) & VN_data_in(8141);
  VN1357_in0 <= VN_sign_in(8142) & VN_data_in(8142);
  VN1357_in1 <= VN_sign_in(8143) & VN_data_in(8143);
  VN1357_in2 <= VN_sign_in(8144) & VN_data_in(8144);
  VN1357_in3 <= VN_sign_in(8145) & VN_data_in(8145);
  VN1357_in4 <= VN_sign_in(8146) & VN_data_in(8146);
  VN1357_in5 <= VN_sign_in(8147) & VN_data_in(8147);
  VN1358_in0 <= VN_sign_in(8148) & VN_data_in(8148);
  VN1358_in1 <= VN_sign_in(8149) & VN_data_in(8149);
  VN1358_in2 <= VN_sign_in(8150) & VN_data_in(8150);
  VN1358_in3 <= VN_sign_in(8151) & VN_data_in(8151);
  VN1358_in4 <= VN_sign_in(8152) & VN_data_in(8152);
  VN1358_in5 <= VN_sign_in(8153) & VN_data_in(8153);
  VN1359_in0 <= VN_sign_in(8154) & VN_data_in(8154);
  VN1359_in1 <= VN_sign_in(8155) & VN_data_in(8155);
  VN1359_in2 <= VN_sign_in(8156) & VN_data_in(8156);
  VN1359_in3 <= VN_sign_in(8157) & VN_data_in(8157);
  VN1359_in4 <= VN_sign_in(8158) & VN_data_in(8158);
  VN1359_in5 <= VN_sign_in(8159) & VN_data_in(8159);
  VN1360_in0 <= VN_sign_in(8160) & VN_data_in(8160);
  VN1360_in1 <= VN_sign_in(8161) & VN_data_in(8161);
  VN1360_in2 <= VN_sign_in(8162) & VN_data_in(8162);
  VN1360_in3 <= VN_sign_in(8163) & VN_data_in(8163);
  VN1360_in4 <= VN_sign_in(8164) & VN_data_in(8164);
  VN1360_in5 <= VN_sign_in(8165) & VN_data_in(8165);
  VN1361_in0 <= VN_sign_in(8166) & VN_data_in(8166);
  VN1361_in1 <= VN_sign_in(8167) & VN_data_in(8167);
  VN1361_in2 <= VN_sign_in(8168) & VN_data_in(8168);
  VN1361_in3 <= VN_sign_in(8169) & VN_data_in(8169);
  VN1361_in4 <= VN_sign_in(8170) & VN_data_in(8170);
  VN1361_in5 <= VN_sign_in(8171) & VN_data_in(8171);
  VN1362_in0 <= VN_sign_in(8172) & VN_data_in(8172);
  VN1362_in1 <= VN_sign_in(8173) & VN_data_in(8173);
  VN1362_in2 <= VN_sign_in(8174) & VN_data_in(8174);
  VN1362_in3 <= VN_sign_in(8175) & VN_data_in(8175);
  VN1362_in4 <= VN_sign_in(8176) & VN_data_in(8176);
  VN1362_in5 <= VN_sign_in(8177) & VN_data_in(8177);
  VN1363_in0 <= VN_sign_in(8178) & VN_data_in(8178);
  VN1363_in1 <= VN_sign_in(8179) & VN_data_in(8179);
  VN1363_in2 <= VN_sign_in(8180) & VN_data_in(8180);
  VN1363_in3 <= VN_sign_in(8181) & VN_data_in(8181);
  VN1363_in4 <= VN_sign_in(8182) & VN_data_in(8182);
  VN1363_in5 <= VN_sign_in(8183) & VN_data_in(8183);
  VN1364_in0 <= VN_sign_in(8184) & VN_data_in(8184);
  VN1364_in1 <= VN_sign_in(8185) & VN_data_in(8185);
  VN1364_in2 <= VN_sign_in(8186) & VN_data_in(8186);
  VN1364_in3 <= VN_sign_in(8187) & VN_data_in(8187);
  VN1364_in4 <= VN_sign_in(8188) & VN_data_in(8188);
  VN1364_in5 <= VN_sign_in(8189) & VN_data_in(8189);
  VN1365_in0 <= VN_sign_in(8190) & VN_data_in(8190);
  VN1365_in1 <= VN_sign_in(8191) & VN_data_in(8191);
  VN1365_in2 <= VN_sign_in(8192) & VN_data_in(8192);
  VN1365_in3 <= VN_sign_in(8193) & VN_data_in(8193);
  VN1365_in4 <= VN_sign_in(8194) & VN_data_in(8194);
  VN1365_in5 <= VN_sign_in(8195) & VN_data_in(8195);
  VN1366_in0 <= VN_sign_in(8196) & VN_data_in(8196);
  VN1366_in1 <= VN_sign_in(8197) & VN_data_in(8197);
  VN1366_in2 <= VN_sign_in(8198) & VN_data_in(8198);
  VN1366_in3 <= VN_sign_in(8199) & VN_data_in(8199);
  VN1366_in4 <= VN_sign_in(8200) & VN_data_in(8200);
  VN1366_in5 <= VN_sign_in(8201) & VN_data_in(8201);
  VN1367_in0 <= VN_sign_in(8202) & VN_data_in(8202);
  VN1367_in1 <= VN_sign_in(8203) & VN_data_in(8203);
  VN1367_in2 <= VN_sign_in(8204) & VN_data_in(8204);
  VN1367_in3 <= VN_sign_in(8205) & VN_data_in(8205);
  VN1367_in4 <= VN_sign_in(8206) & VN_data_in(8206);
  VN1367_in5 <= VN_sign_in(8207) & VN_data_in(8207);
  VN1368_in0 <= VN_sign_in(8208) & VN_data_in(8208);
  VN1368_in1 <= VN_sign_in(8209) & VN_data_in(8209);
  VN1368_in2 <= VN_sign_in(8210) & VN_data_in(8210);
  VN1368_in3 <= VN_sign_in(8211) & VN_data_in(8211);
  VN1368_in4 <= VN_sign_in(8212) & VN_data_in(8212);
  VN1368_in5 <= VN_sign_in(8213) & VN_data_in(8213);
  VN1369_in0 <= VN_sign_in(8214) & VN_data_in(8214);
  VN1369_in1 <= VN_sign_in(8215) & VN_data_in(8215);
  VN1369_in2 <= VN_sign_in(8216) & VN_data_in(8216);
  VN1369_in3 <= VN_sign_in(8217) & VN_data_in(8217);
  VN1369_in4 <= VN_sign_in(8218) & VN_data_in(8218);
  VN1369_in5 <= VN_sign_in(8219) & VN_data_in(8219);
  VN1370_in0 <= VN_sign_in(8220) & VN_data_in(8220);
  VN1370_in1 <= VN_sign_in(8221) & VN_data_in(8221);
  VN1370_in2 <= VN_sign_in(8222) & VN_data_in(8222);
  VN1370_in3 <= VN_sign_in(8223) & VN_data_in(8223);
  VN1370_in4 <= VN_sign_in(8224) & VN_data_in(8224);
  VN1370_in5 <= VN_sign_in(8225) & VN_data_in(8225);
  VN1371_in0 <= VN_sign_in(8226) & VN_data_in(8226);
  VN1371_in1 <= VN_sign_in(8227) & VN_data_in(8227);
  VN1371_in2 <= VN_sign_in(8228) & VN_data_in(8228);
  VN1371_in3 <= VN_sign_in(8229) & VN_data_in(8229);
  VN1371_in4 <= VN_sign_in(8230) & VN_data_in(8230);
  VN1371_in5 <= VN_sign_in(8231) & VN_data_in(8231);
  VN1372_in0 <= VN_sign_in(8232) & VN_data_in(8232);
  VN1372_in1 <= VN_sign_in(8233) & VN_data_in(8233);
  VN1372_in2 <= VN_sign_in(8234) & VN_data_in(8234);
  VN1372_in3 <= VN_sign_in(8235) & VN_data_in(8235);
  VN1372_in4 <= VN_sign_in(8236) & VN_data_in(8236);
  VN1372_in5 <= VN_sign_in(8237) & VN_data_in(8237);
  VN1373_in0 <= VN_sign_in(8238) & VN_data_in(8238);
  VN1373_in1 <= VN_sign_in(8239) & VN_data_in(8239);
  VN1373_in2 <= VN_sign_in(8240) & VN_data_in(8240);
  VN1373_in3 <= VN_sign_in(8241) & VN_data_in(8241);
  VN1373_in4 <= VN_sign_in(8242) & VN_data_in(8242);
  VN1373_in5 <= VN_sign_in(8243) & VN_data_in(8243);
  VN1374_in0 <= VN_sign_in(8244) & VN_data_in(8244);
  VN1374_in1 <= VN_sign_in(8245) & VN_data_in(8245);
  VN1374_in2 <= VN_sign_in(8246) & VN_data_in(8246);
  VN1374_in3 <= VN_sign_in(8247) & VN_data_in(8247);
  VN1374_in4 <= VN_sign_in(8248) & VN_data_in(8248);
  VN1374_in5 <= VN_sign_in(8249) & VN_data_in(8249);
  VN1375_in0 <= VN_sign_in(8250) & VN_data_in(8250);
  VN1375_in1 <= VN_sign_in(8251) & VN_data_in(8251);
  VN1375_in2 <= VN_sign_in(8252) & VN_data_in(8252);
  VN1375_in3 <= VN_sign_in(8253) & VN_data_in(8253);
  VN1375_in4 <= VN_sign_in(8254) & VN_data_in(8254);
  VN1375_in5 <= VN_sign_in(8255) & VN_data_in(8255);
  VN1376_in0 <= VN_sign_in(8256) & VN_data_in(8256);
  VN1376_in1 <= VN_sign_in(8257) & VN_data_in(8257);
  VN1376_in2 <= VN_sign_in(8258) & VN_data_in(8258);
  VN1376_in3 <= VN_sign_in(8259) & VN_data_in(8259);
  VN1376_in4 <= VN_sign_in(8260) & VN_data_in(8260);
  VN1376_in5 <= VN_sign_in(8261) & VN_data_in(8261);
  VN1377_in0 <= VN_sign_in(8262) & VN_data_in(8262);
  VN1377_in1 <= VN_sign_in(8263) & VN_data_in(8263);
  VN1377_in2 <= VN_sign_in(8264) & VN_data_in(8264);
  VN1377_in3 <= VN_sign_in(8265) & VN_data_in(8265);
  VN1377_in4 <= VN_sign_in(8266) & VN_data_in(8266);
  VN1377_in5 <= VN_sign_in(8267) & VN_data_in(8267);
  VN1378_in0 <= VN_sign_in(8268) & VN_data_in(8268);
  VN1378_in1 <= VN_sign_in(8269) & VN_data_in(8269);
  VN1378_in2 <= VN_sign_in(8270) & VN_data_in(8270);
  VN1378_in3 <= VN_sign_in(8271) & VN_data_in(8271);
  VN1378_in4 <= VN_sign_in(8272) & VN_data_in(8272);
  VN1378_in5 <= VN_sign_in(8273) & VN_data_in(8273);
  VN1379_in0 <= VN_sign_in(8274) & VN_data_in(8274);
  VN1379_in1 <= VN_sign_in(8275) & VN_data_in(8275);
  VN1379_in2 <= VN_sign_in(8276) & VN_data_in(8276);
  VN1379_in3 <= VN_sign_in(8277) & VN_data_in(8277);
  VN1379_in4 <= VN_sign_in(8278) & VN_data_in(8278);
  VN1379_in5 <= VN_sign_in(8279) & VN_data_in(8279);
  VN1380_in0 <= VN_sign_in(8280) & VN_data_in(8280);
  VN1380_in1 <= VN_sign_in(8281) & VN_data_in(8281);
  VN1380_in2 <= VN_sign_in(8282) & VN_data_in(8282);
  VN1380_in3 <= VN_sign_in(8283) & VN_data_in(8283);
  VN1380_in4 <= VN_sign_in(8284) & VN_data_in(8284);
  VN1380_in5 <= VN_sign_in(8285) & VN_data_in(8285);
  VN1381_in0 <= VN_sign_in(8286) & VN_data_in(8286);
  VN1381_in1 <= VN_sign_in(8287) & VN_data_in(8287);
  VN1381_in2 <= VN_sign_in(8288) & VN_data_in(8288);
  VN1381_in3 <= VN_sign_in(8289) & VN_data_in(8289);
  VN1381_in4 <= VN_sign_in(8290) & VN_data_in(8290);
  VN1381_in5 <= VN_sign_in(8291) & VN_data_in(8291);
  VN1382_in0 <= VN_sign_in(8292) & VN_data_in(8292);
  VN1382_in1 <= VN_sign_in(8293) & VN_data_in(8293);
  VN1382_in2 <= VN_sign_in(8294) & VN_data_in(8294);
  VN1382_in3 <= VN_sign_in(8295) & VN_data_in(8295);
  VN1382_in4 <= VN_sign_in(8296) & VN_data_in(8296);
  VN1382_in5 <= VN_sign_in(8297) & VN_data_in(8297);
  VN1383_in0 <= VN_sign_in(8298) & VN_data_in(8298);
  VN1383_in1 <= VN_sign_in(8299) & VN_data_in(8299);
  VN1383_in2 <= VN_sign_in(8300) & VN_data_in(8300);
  VN1383_in3 <= VN_sign_in(8301) & VN_data_in(8301);
  VN1383_in4 <= VN_sign_in(8302) & VN_data_in(8302);
  VN1383_in5 <= VN_sign_in(8303) & VN_data_in(8303);
  VN1384_in0 <= VN_sign_in(8304) & VN_data_in(8304);
  VN1384_in1 <= VN_sign_in(8305) & VN_data_in(8305);
  VN1384_in2 <= VN_sign_in(8306) & VN_data_in(8306);
  VN1384_in3 <= VN_sign_in(8307) & VN_data_in(8307);
  VN1384_in4 <= VN_sign_in(8308) & VN_data_in(8308);
  VN1384_in5 <= VN_sign_in(8309) & VN_data_in(8309);
  VN1385_in0 <= VN_sign_in(8310) & VN_data_in(8310);
  VN1385_in1 <= VN_sign_in(8311) & VN_data_in(8311);
  VN1385_in2 <= VN_sign_in(8312) & VN_data_in(8312);
  VN1385_in3 <= VN_sign_in(8313) & VN_data_in(8313);
  VN1385_in4 <= VN_sign_in(8314) & VN_data_in(8314);
  VN1385_in5 <= VN_sign_in(8315) & VN_data_in(8315);
  VN1386_in0 <= VN_sign_in(8316) & VN_data_in(8316);
  VN1386_in1 <= VN_sign_in(8317) & VN_data_in(8317);
  VN1386_in2 <= VN_sign_in(8318) & VN_data_in(8318);
  VN1386_in3 <= VN_sign_in(8319) & VN_data_in(8319);
  VN1386_in4 <= VN_sign_in(8320) & VN_data_in(8320);
  VN1386_in5 <= VN_sign_in(8321) & VN_data_in(8321);
  VN1387_in0 <= VN_sign_in(8322) & VN_data_in(8322);
  VN1387_in1 <= VN_sign_in(8323) & VN_data_in(8323);
  VN1387_in2 <= VN_sign_in(8324) & VN_data_in(8324);
  VN1387_in3 <= VN_sign_in(8325) & VN_data_in(8325);
  VN1387_in4 <= VN_sign_in(8326) & VN_data_in(8326);
  VN1387_in5 <= VN_sign_in(8327) & VN_data_in(8327);
  VN1388_in0 <= VN_sign_in(8328) & VN_data_in(8328);
  VN1388_in1 <= VN_sign_in(8329) & VN_data_in(8329);
  VN1388_in2 <= VN_sign_in(8330) & VN_data_in(8330);
  VN1388_in3 <= VN_sign_in(8331) & VN_data_in(8331);
  VN1388_in4 <= VN_sign_in(8332) & VN_data_in(8332);
  VN1388_in5 <= VN_sign_in(8333) & VN_data_in(8333);
  VN1389_in0 <= VN_sign_in(8334) & VN_data_in(8334);
  VN1389_in1 <= VN_sign_in(8335) & VN_data_in(8335);
  VN1389_in2 <= VN_sign_in(8336) & VN_data_in(8336);
  VN1389_in3 <= VN_sign_in(8337) & VN_data_in(8337);
  VN1389_in4 <= VN_sign_in(8338) & VN_data_in(8338);
  VN1389_in5 <= VN_sign_in(8339) & VN_data_in(8339);
  VN1390_in0 <= VN_sign_in(8340) & VN_data_in(8340);
  VN1390_in1 <= VN_sign_in(8341) & VN_data_in(8341);
  VN1390_in2 <= VN_sign_in(8342) & VN_data_in(8342);
  VN1390_in3 <= VN_sign_in(8343) & VN_data_in(8343);
  VN1390_in4 <= VN_sign_in(8344) & VN_data_in(8344);
  VN1390_in5 <= VN_sign_in(8345) & VN_data_in(8345);
  VN1391_in0 <= VN_sign_in(8346) & VN_data_in(8346);
  VN1391_in1 <= VN_sign_in(8347) & VN_data_in(8347);
  VN1391_in2 <= VN_sign_in(8348) & VN_data_in(8348);
  VN1391_in3 <= VN_sign_in(8349) & VN_data_in(8349);
  VN1391_in4 <= VN_sign_in(8350) & VN_data_in(8350);
  VN1391_in5 <= VN_sign_in(8351) & VN_data_in(8351);
  VN1392_in0 <= VN_sign_in(8352) & VN_data_in(8352);
  VN1392_in1 <= VN_sign_in(8353) & VN_data_in(8353);
  VN1392_in2 <= VN_sign_in(8354) & VN_data_in(8354);
  VN1392_in3 <= VN_sign_in(8355) & VN_data_in(8355);
  VN1392_in4 <= VN_sign_in(8356) & VN_data_in(8356);
  VN1392_in5 <= VN_sign_in(8357) & VN_data_in(8357);
  VN1393_in0 <= VN_sign_in(8358) & VN_data_in(8358);
  VN1393_in1 <= VN_sign_in(8359) & VN_data_in(8359);
  VN1393_in2 <= VN_sign_in(8360) & VN_data_in(8360);
  VN1393_in3 <= VN_sign_in(8361) & VN_data_in(8361);
  VN1393_in4 <= VN_sign_in(8362) & VN_data_in(8362);
  VN1393_in5 <= VN_sign_in(8363) & VN_data_in(8363);
  VN1394_in0 <= VN_sign_in(8364) & VN_data_in(8364);
  VN1394_in1 <= VN_sign_in(8365) & VN_data_in(8365);
  VN1394_in2 <= VN_sign_in(8366) & VN_data_in(8366);
  VN1394_in3 <= VN_sign_in(8367) & VN_data_in(8367);
  VN1394_in4 <= VN_sign_in(8368) & VN_data_in(8368);
  VN1394_in5 <= VN_sign_in(8369) & VN_data_in(8369);
  VN1395_in0 <= VN_sign_in(8370) & VN_data_in(8370);
  VN1395_in1 <= VN_sign_in(8371) & VN_data_in(8371);
  VN1395_in2 <= VN_sign_in(8372) & VN_data_in(8372);
  VN1395_in3 <= VN_sign_in(8373) & VN_data_in(8373);
  VN1395_in4 <= VN_sign_in(8374) & VN_data_in(8374);
  VN1395_in5 <= VN_sign_in(8375) & VN_data_in(8375);
  VN1396_in0 <= VN_sign_in(8376) & VN_data_in(8376);
  VN1396_in1 <= VN_sign_in(8377) & VN_data_in(8377);
  VN1396_in2 <= VN_sign_in(8378) & VN_data_in(8378);
  VN1396_in3 <= VN_sign_in(8379) & VN_data_in(8379);
  VN1396_in4 <= VN_sign_in(8380) & VN_data_in(8380);
  VN1396_in5 <= VN_sign_in(8381) & VN_data_in(8381);
  VN1397_in0 <= VN_sign_in(8382) & VN_data_in(8382);
  VN1397_in1 <= VN_sign_in(8383) & VN_data_in(8383);
  VN1397_in2 <= VN_sign_in(8384) & VN_data_in(8384);
  VN1397_in3 <= VN_sign_in(8385) & VN_data_in(8385);
  VN1397_in4 <= VN_sign_in(8386) & VN_data_in(8386);
  VN1397_in5 <= VN_sign_in(8387) & VN_data_in(8387);
  VN1398_in0 <= VN_sign_in(8388) & VN_data_in(8388);
  VN1398_in1 <= VN_sign_in(8389) & VN_data_in(8389);
  VN1398_in2 <= VN_sign_in(8390) & VN_data_in(8390);
  VN1398_in3 <= VN_sign_in(8391) & VN_data_in(8391);
  VN1398_in4 <= VN_sign_in(8392) & VN_data_in(8392);
  VN1398_in5 <= VN_sign_in(8393) & VN_data_in(8393);
  VN1399_in0 <= VN_sign_in(8394) & VN_data_in(8394);
  VN1399_in1 <= VN_sign_in(8395) & VN_data_in(8395);
  VN1399_in2 <= VN_sign_in(8396) & VN_data_in(8396);
  VN1399_in3 <= VN_sign_in(8397) & VN_data_in(8397);
  VN1399_in4 <= VN_sign_in(8398) & VN_data_in(8398);
  VN1399_in5 <= VN_sign_in(8399) & VN_data_in(8399);
  VN1400_in0 <= VN_sign_in(8400) & VN_data_in(8400);
  VN1400_in1 <= VN_sign_in(8401) & VN_data_in(8401);
  VN1400_in2 <= VN_sign_in(8402) & VN_data_in(8402);
  VN1400_in3 <= VN_sign_in(8403) & VN_data_in(8403);
  VN1400_in4 <= VN_sign_in(8404) & VN_data_in(8404);
  VN1400_in5 <= VN_sign_in(8405) & VN_data_in(8405);
  VN1401_in0 <= VN_sign_in(8406) & VN_data_in(8406);
  VN1401_in1 <= VN_sign_in(8407) & VN_data_in(8407);
  VN1401_in2 <= VN_sign_in(8408) & VN_data_in(8408);
  VN1401_in3 <= VN_sign_in(8409) & VN_data_in(8409);
  VN1401_in4 <= VN_sign_in(8410) & VN_data_in(8410);
  VN1401_in5 <= VN_sign_in(8411) & VN_data_in(8411);
  VN1402_in0 <= VN_sign_in(8412) & VN_data_in(8412);
  VN1402_in1 <= VN_sign_in(8413) & VN_data_in(8413);
  VN1402_in2 <= VN_sign_in(8414) & VN_data_in(8414);
  VN1402_in3 <= VN_sign_in(8415) & VN_data_in(8415);
  VN1402_in4 <= VN_sign_in(8416) & VN_data_in(8416);
  VN1402_in5 <= VN_sign_in(8417) & VN_data_in(8417);
  VN1403_in0 <= VN_sign_in(8418) & VN_data_in(8418);
  VN1403_in1 <= VN_sign_in(8419) & VN_data_in(8419);
  VN1403_in2 <= VN_sign_in(8420) & VN_data_in(8420);
  VN1403_in3 <= VN_sign_in(8421) & VN_data_in(8421);
  VN1403_in4 <= VN_sign_in(8422) & VN_data_in(8422);
  VN1403_in5 <= VN_sign_in(8423) & VN_data_in(8423);
  VN1404_in0 <= VN_sign_in(8424) & VN_data_in(8424);
  VN1404_in1 <= VN_sign_in(8425) & VN_data_in(8425);
  VN1404_in2 <= VN_sign_in(8426) & VN_data_in(8426);
  VN1404_in3 <= VN_sign_in(8427) & VN_data_in(8427);
  VN1404_in4 <= VN_sign_in(8428) & VN_data_in(8428);
  VN1404_in5 <= VN_sign_in(8429) & VN_data_in(8429);
  VN1405_in0 <= VN_sign_in(8430) & VN_data_in(8430);
  VN1405_in1 <= VN_sign_in(8431) & VN_data_in(8431);
  VN1405_in2 <= VN_sign_in(8432) & VN_data_in(8432);
  VN1405_in3 <= VN_sign_in(8433) & VN_data_in(8433);
  VN1405_in4 <= VN_sign_in(8434) & VN_data_in(8434);
  VN1405_in5 <= VN_sign_in(8435) & VN_data_in(8435);
  VN1406_in0 <= VN_sign_in(8436) & VN_data_in(8436);
  VN1406_in1 <= VN_sign_in(8437) & VN_data_in(8437);
  VN1406_in2 <= VN_sign_in(8438) & VN_data_in(8438);
  VN1406_in3 <= VN_sign_in(8439) & VN_data_in(8439);
  VN1406_in4 <= VN_sign_in(8440) & VN_data_in(8440);
  VN1406_in5 <= VN_sign_in(8441) & VN_data_in(8441);
  VN1407_in0 <= VN_sign_in(8442) & VN_data_in(8442);
  VN1407_in1 <= VN_sign_in(8443) & VN_data_in(8443);
  VN1407_in2 <= VN_sign_in(8444) & VN_data_in(8444);
  VN1407_in3 <= VN_sign_in(8445) & VN_data_in(8445);
  VN1407_in4 <= VN_sign_in(8446) & VN_data_in(8446);
  VN1407_in5 <= VN_sign_in(8447) & VN_data_in(8447);
  VN1408_in0 <= VN_sign_in(8448) & VN_data_in(8448);
  VN1408_in1 <= VN_sign_in(8449) & VN_data_in(8449);
  VN1408_in2 <= VN_sign_in(8450) & VN_data_in(8450);
  VN1408_in3 <= VN_sign_in(8451) & VN_data_in(8451);
  VN1408_in4 <= VN_sign_in(8452) & VN_data_in(8452);
  VN1408_in5 <= VN_sign_in(8453) & VN_data_in(8453);
  VN1409_in0 <= VN_sign_in(8454) & VN_data_in(8454);
  VN1409_in1 <= VN_sign_in(8455) & VN_data_in(8455);
  VN1409_in2 <= VN_sign_in(8456) & VN_data_in(8456);
  VN1409_in3 <= VN_sign_in(8457) & VN_data_in(8457);
  VN1409_in4 <= VN_sign_in(8458) & VN_data_in(8458);
  VN1409_in5 <= VN_sign_in(8459) & VN_data_in(8459);
  VN1410_in0 <= VN_sign_in(8460) & VN_data_in(8460);
  VN1410_in1 <= VN_sign_in(8461) & VN_data_in(8461);
  VN1410_in2 <= VN_sign_in(8462) & VN_data_in(8462);
  VN1410_in3 <= VN_sign_in(8463) & VN_data_in(8463);
  VN1410_in4 <= VN_sign_in(8464) & VN_data_in(8464);
  VN1410_in5 <= VN_sign_in(8465) & VN_data_in(8465);
  VN1411_in0 <= VN_sign_in(8466) & VN_data_in(8466);
  VN1411_in1 <= VN_sign_in(8467) & VN_data_in(8467);
  VN1411_in2 <= VN_sign_in(8468) & VN_data_in(8468);
  VN1411_in3 <= VN_sign_in(8469) & VN_data_in(8469);
  VN1411_in4 <= VN_sign_in(8470) & VN_data_in(8470);
  VN1411_in5 <= VN_sign_in(8471) & VN_data_in(8471);
  VN1412_in0 <= VN_sign_in(8472) & VN_data_in(8472);
  VN1412_in1 <= VN_sign_in(8473) & VN_data_in(8473);
  VN1412_in2 <= VN_sign_in(8474) & VN_data_in(8474);
  VN1412_in3 <= VN_sign_in(8475) & VN_data_in(8475);
  VN1412_in4 <= VN_sign_in(8476) & VN_data_in(8476);
  VN1412_in5 <= VN_sign_in(8477) & VN_data_in(8477);
  VN1413_in0 <= VN_sign_in(8478) & VN_data_in(8478);
  VN1413_in1 <= VN_sign_in(8479) & VN_data_in(8479);
  VN1413_in2 <= VN_sign_in(8480) & VN_data_in(8480);
  VN1413_in3 <= VN_sign_in(8481) & VN_data_in(8481);
  VN1413_in4 <= VN_sign_in(8482) & VN_data_in(8482);
  VN1413_in5 <= VN_sign_in(8483) & VN_data_in(8483);
  VN1414_in0 <= VN_sign_in(8484) & VN_data_in(8484);
  VN1414_in1 <= VN_sign_in(8485) & VN_data_in(8485);
  VN1414_in2 <= VN_sign_in(8486) & VN_data_in(8486);
  VN1414_in3 <= VN_sign_in(8487) & VN_data_in(8487);
  VN1414_in4 <= VN_sign_in(8488) & VN_data_in(8488);
  VN1414_in5 <= VN_sign_in(8489) & VN_data_in(8489);
  VN1415_in0 <= VN_sign_in(8490) & VN_data_in(8490);
  VN1415_in1 <= VN_sign_in(8491) & VN_data_in(8491);
  VN1415_in2 <= VN_sign_in(8492) & VN_data_in(8492);
  VN1415_in3 <= VN_sign_in(8493) & VN_data_in(8493);
  VN1415_in4 <= VN_sign_in(8494) & VN_data_in(8494);
  VN1415_in5 <= VN_sign_in(8495) & VN_data_in(8495);
  VN1416_in0 <= VN_sign_in(8496) & VN_data_in(8496);
  VN1416_in1 <= VN_sign_in(8497) & VN_data_in(8497);
  VN1416_in2 <= VN_sign_in(8498) & VN_data_in(8498);
  VN1416_in3 <= VN_sign_in(8499) & VN_data_in(8499);
  VN1416_in4 <= VN_sign_in(8500) & VN_data_in(8500);
  VN1416_in5 <= VN_sign_in(8501) & VN_data_in(8501);
  VN1417_in0 <= VN_sign_in(8502) & VN_data_in(8502);
  VN1417_in1 <= VN_sign_in(8503) & VN_data_in(8503);
  VN1417_in2 <= VN_sign_in(8504) & VN_data_in(8504);
  VN1417_in3 <= VN_sign_in(8505) & VN_data_in(8505);
  VN1417_in4 <= VN_sign_in(8506) & VN_data_in(8506);
  VN1417_in5 <= VN_sign_in(8507) & VN_data_in(8507);
  VN1418_in0 <= VN_sign_in(8508) & VN_data_in(8508);
  VN1418_in1 <= VN_sign_in(8509) & VN_data_in(8509);
  VN1418_in2 <= VN_sign_in(8510) & VN_data_in(8510);
  VN1418_in3 <= VN_sign_in(8511) & VN_data_in(8511);
  VN1418_in4 <= VN_sign_in(8512) & VN_data_in(8512);
  VN1418_in5 <= VN_sign_in(8513) & VN_data_in(8513);
  VN1419_in0 <= VN_sign_in(8514) & VN_data_in(8514);
  VN1419_in1 <= VN_sign_in(8515) & VN_data_in(8515);
  VN1419_in2 <= VN_sign_in(8516) & VN_data_in(8516);
  VN1419_in3 <= VN_sign_in(8517) & VN_data_in(8517);
  VN1419_in4 <= VN_sign_in(8518) & VN_data_in(8518);
  VN1419_in5 <= VN_sign_in(8519) & VN_data_in(8519);
  VN1420_in0 <= VN_sign_in(8520) & VN_data_in(8520);
  VN1420_in1 <= VN_sign_in(8521) & VN_data_in(8521);
  VN1420_in2 <= VN_sign_in(8522) & VN_data_in(8522);
  VN1420_in3 <= VN_sign_in(8523) & VN_data_in(8523);
  VN1420_in4 <= VN_sign_in(8524) & VN_data_in(8524);
  VN1420_in5 <= VN_sign_in(8525) & VN_data_in(8525);
  VN1421_in0 <= VN_sign_in(8526) & VN_data_in(8526);
  VN1421_in1 <= VN_sign_in(8527) & VN_data_in(8527);
  VN1421_in2 <= VN_sign_in(8528) & VN_data_in(8528);
  VN1421_in3 <= VN_sign_in(8529) & VN_data_in(8529);
  VN1421_in4 <= VN_sign_in(8530) & VN_data_in(8530);
  VN1421_in5 <= VN_sign_in(8531) & VN_data_in(8531);
  VN1422_in0 <= VN_sign_in(8532) & VN_data_in(8532);
  VN1422_in1 <= VN_sign_in(8533) & VN_data_in(8533);
  VN1422_in2 <= VN_sign_in(8534) & VN_data_in(8534);
  VN1422_in3 <= VN_sign_in(8535) & VN_data_in(8535);
  VN1422_in4 <= VN_sign_in(8536) & VN_data_in(8536);
  VN1422_in5 <= VN_sign_in(8537) & VN_data_in(8537);
  VN1423_in0 <= VN_sign_in(8538) & VN_data_in(8538);
  VN1423_in1 <= VN_sign_in(8539) & VN_data_in(8539);
  VN1423_in2 <= VN_sign_in(8540) & VN_data_in(8540);
  VN1423_in3 <= VN_sign_in(8541) & VN_data_in(8541);
  VN1423_in4 <= VN_sign_in(8542) & VN_data_in(8542);
  VN1423_in5 <= VN_sign_in(8543) & VN_data_in(8543);
  VN1424_in0 <= VN_sign_in(8544) & VN_data_in(8544);
  VN1424_in1 <= VN_sign_in(8545) & VN_data_in(8545);
  VN1424_in2 <= VN_sign_in(8546) & VN_data_in(8546);
  VN1424_in3 <= VN_sign_in(8547) & VN_data_in(8547);
  VN1424_in4 <= VN_sign_in(8548) & VN_data_in(8548);
  VN1424_in5 <= VN_sign_in(8549) & VN_data_in(8549);
  VN1425_in0 <= VN_sign_in(8550) & VN_data_in(8550);
  VN1425_in1 <= VN_sign_in(8551) & VN_data_in(8551);
  VN1425_in2 <= VN_sign_in(8552) & VN_data_in(8552);
  VN1425_in3 <= VN_sign_in(8553) & VN_data_in(8553);
  VN1425_in4 <= VN_sign_in(8554) & VN_data_in(8554);
  VN1425_in5 <= VN_sign_in(8555) & VN_data_in(8555);
  VN1426_in0 <= VN_sign_in(8556) & VN_data_in(8556);
  VN1426_in1 <= VN_sign_in(8557) & VN_data_in(8557);
  VN1426_in2 <= VN_sign_in(8558) & VN_data_in(8558);
  VN1426_in3 <= VN_sign_in(8559) & VN_data_in(8559);
  VN1426_in4 <= VN_sign_in(8560) & VN_data_in(8560);
  VN1426_in5 <= VN_sign_in(8561) & VN_data_in(8561);
  VN1427_in0 <= VN_sign_in(8562) & VN_data_in(8562);
  VN1427_in1 <= VN_sign_in(8563) & VN_data_in(8563);
  VN1427_in2 <= VN_sign_in(8564) & VN_data_in(8564);
  VN1427_in3 <= VN_sign_in(8565) & VN_data_in(8565);
  VN1427_in4 <= VN_sign_in(8566) & VN_data_in(8566);
  VN1427_in5 <= VN_sign_in(8567) & VN_data_in(8567);
  VN1428_in0 <= VN_sign_in(8568) & VN_data_in(8568);
  VN1428_in1 <= VN_sign_in(8569) & VN_data_in(8569);
  VN1428_in2 <= VN_sign_in(8570) & VN_data_in(8570);
  VN1428_in3 <= VN_sign_in(8571) & VN_data_in(8571);
  VN1428_in4 <= VN_sign_in(8572) & VN_data_in(8572);
  VN1428_in5 <= VN_sign_in(8573) & VN_data_in(8573);
  VN1429_in0 <= VN_sign_in(8574) & VN_data_in(8574);
  VN1429_in1 <= VN_sign_in(8575) & VN_data_in(8575);
  VN1429_in2 <= VN_sign_in(8576) & VN_data_in(8576);
  VN1429_in3 <= VN_sign_in(8577) & VN_data_in(8577);
  VN1429_in4 <= VN_sign_in(8578) & VN_data_in(8578);
  VN1429_in5 <= VN_sign_in(8579) & VN_data_in(8579);
  VN1430_in0 <= VN_sign_in(8580) & VN_data_in(8580);
  VN1430_in1 <= VN_sign_in(8581) & VN_data_in(8581);
  VN1430_in2 <= VN_sign_in(8582) & VN_data_in(8582);
  VN1430_in3 <= VN_sign_in(8583) & VN_data_in(8583);
  VN1430_in4 <= VN_sign_in(8584) & VN_data_in(8584);
  VN1430_in5 <= VN_sign_in(8585) & VN_data_in(8585);
  VN1431_in0 <= VN_sign_in(8586) & VN_data_in(8586);
  VN1431_in1 <= VN_sign_in(8587) & VN_data_in(8587);
  VN1431_in2 <= VN_sign_in(8588) & VN_data_in(8588);
  VN1431_in3 <= VN_sign_in(8589) & VN_data_in(8589);
  VN1431_in4 <= VN_sign_in(8590) & VN_data_in(8590);
  VN1431_in5 <= VN_sign_in(8591) & VN_data_in(8591);
  VN1432_in0 <= VN_sign_in(8592) & VN_data_in(8592);
  VN1432_in1 <= VN_sign_in(8593) & VN_data_in(8593);
  VN1432_in2 <= VN_sign_in(8594) & VN_data_in(8594);
  VN1432_in3 <= VN_sign_in(8595) & VN_data_in(8595);
  VN1432_in4 <= VN_sign_in(8596) & VN_data_in(8596);
  VN1432_in5 <= VN_sign_in(8597) & VN_data_in(8597);
  VN1433_in0 <= VN_sign_in(8598) & VN_data_in(8598);
  VN1433_in1 <= VN_sign_in(8599) & VN_data_in(8599);
  VN1433_in2 <= VN_sign_in(8600) & VN_data_in(8600);
  VN1433_in3 <= VN_sign_in(8601) & VN_data_in(8601);
  VN1433_in4 <= VN_sign_in(8602) & VN_data_in(8602);
  VN1433_in5 <= VN_sign_in(8603) & VN_data_in(8603);
  VN1434_in0 <= VN_sign_in(8604) & VN_data_in(8604);
  VN1434_in1 <= VN_sign_in(8605) & VN_data_in(8605);
  VN1434_in2 <= VN_sign_in(8606) & VN_data_in(8606);
  VN1434_in3 <= VN_sign_in(8607) & VN_data_in(8607);
  VN1434_in4 <= VN_sign_in(8608) & VN_data_in(8608);
  VN1434_in5 <= VN_sign_in(8609) & VN_data_in(8609);
  VN1435_in0 <= VN_sign_in(8610) & VN_data_in(8610);
  VN1435_in1 <= VN_sign_in(8611) & VN_data_in(8611);
  VN1435_in2 <= VN_sign_in(8612) & VN_data_in(8612);
  VN1435_in3 <= VN_sign_in(8613) & VN_data_in(8613);
  VN1435_in4 <= VN_sign_in(8614) & VN_data_in(8614);
  VN1435_in5 <= VN_sign_in(8615) & VN_data_in(8615);
  VN1436_in0 <= VN_sign_in(8616) & VN_data_in(8616);
  VN1436_in1 <= VN_sign_in(8617) & VN_data_in(8617);
  VN1436_in2 <= VN_sign_in(8618) & VN_data_in(8618);
  VN1436_in3 <= VN_sign_in(8619) & VN_data_in(8619);
  VN1436_in4 <= VN_sign_in(8620) & VN_data_in(8620);
  VN1436_in5 <= VN_sign_in(8621) & VN_data_in(8621);
  VN1437_in0 <= VN_sign_in(8622) & VN_data_in(8622);
  VN1437_in1 <= VN_sign_in(8623) & VN_data_in(8623);
  VN1437_in2 <= VN_sign_in(8624) & VN_data_in(8624);
  VN1437_in3 <= VN_sign_in(8625) & VN_data_in(8625);
  VN1437_in4 <= VN_sign_in(8626) & VN_data_in(8626);
  VN1437_in5 <= VN_sign_in(8627) & VN_data_in(8627);
  VN1438_in0 <= VN_sign_in(8628) & VN_data_in(8628);
  VN1438_in1 <= VN_sign_in(8629) & VN_data_in(8629);
  VN1438_in2 <= VN_sign_in(8630) & VN_data_in(8630);
  VN1438_in3 <= VN_sign_in(8631) & VN_data_in(8631);
  VN1438_in4 <= VN_sign_in(8632) & VN_data_in(8632);
  VN1438_in5 <= VN_sign_in(8633) & VN_data_in(8633);
  VN1439_in0 <= VN_sign_in(8634) & VN_data_in(8634);
  VN1439_in1 <= VN_sign_in(8635) & VN_data_in(8635);
  VN1439_in2 <= VN_sign_in(8636) & VN_data_in(8636);
  VN1439_in3 <= VN_sign_in(8637) & VN_data_in(8637);
  VN1439_in4 <= VN_sign_in(8638) & VN_data_in(8638);
  VN1439_in5 <= VN_sign_in(8639) & VN_data_in(8639);
  VN1440_in0 <= VN_sign_in(8640) & VN_data_in(8640);
  VN1440_in1 <= VN_sign_in(8641) & VN_data_in(8641);
  VN1440_in2 <= VN_sign_in(8642) & VN_data_in(8642);
  VN1440_in3 <= VN_sign_in(8643) & VN_data_in(8643);
  VN1440_in4 <= VN_sign_in(8644) & VN_data_in(8644);
  VN1440_in5 <= VN_sign_in(8645) & VN_data_in(8645);
  VN1441_in0 <= VN_sign_in(8646) & VN_data_in(8646);
  VN1441_in1 <= VN_sign_in(8647) & VN_data_in(8647);
  VN1441_in2 <= VN_sign_in(8648) & VN_data_in(8648);
  VN1441_in3 <= VN_sign_in(8649) & VN_data_in(8649);
  VN1441_in4 <= VN_sign_in(8650) & VN_data_in(8650);
  VN1441_in5 <= VN_sign_in(8651) & VN_data_in(8651);
  VN1442_in0 <= VN_sign_in(8652) & VN_data_in(8652);
  VN1442_in1 <= VN_sign_in(8653) & VN_data_in(8653);
  VN1442_in2 <= VN_sign_in(8654) & VN_data_in(8654);
  VN1442_in3 <= VN_sign_in(8655) & VN_data_in(8655);
  VN1442_in4 <= VN_sign_in(8656) & VN_data_in(8656);
  VN1442_in5 <= VN_sign_in(8657) & VN_data_in(8657);
  VN1443_in0 <= VN_sign_in(8658) & VN_data_in(8658);
  VN1443_in1 <= VN_sign_in(8659) & VN_data_in(8659);
  VN1443_in2 <= VN_sign_in(8660) & VN_data_in(8660);
  VN1443_in3 <= VN_sign_in(8661) & VN_data_in(8661);
  VN1443_in4 <= VN_sign_in(8662) & VN_data_in(8662);
  VN1443_in5 <= VN_sign_in(8663) & VN_data_in(8663);
  VN1444_in0 <= VN_sign_in(8664) & VN_data_in(8664);
  VN1444_in1 <= VN_sign_in(8665) & VN_data_in(8665);
  VN1444_in2 <= VN_sign_in(8666) & VN_data_in(8666);
  VN1444_in3 <= VN_sign_in(8667) & VN_data_in(8667);
  VN1444_in4 <= VN_sign_in(8668) & VN_data_in(8668);
  VN1444_in5 <= VN_sign_in(8669) & VN_data_in(8669);
  VN1445_in0 <= VN_sign_in(8670) & VN_data_in(8670);
  VN1445_in1 <= VN_sign_in(8671) & VN_data_in(8671);
  VN1445_in2 <= VN_sign_in(8672) & VN_data_in(8672);
  VN1445_in3 <= VN_sign_in(8673) & VN_data_in(8673);
  VN1445_in4 <= VN_sign_in(8674) & VN_data_in(8674);
  VN1445_in5 <= VN_sign_in(8675) & VN_data_in(8675);
  VN1446_in0 <= VN_sign_in(8676) & VN_data_in(8676);
  VN1446_in1 <= VN_sign_in(8677) & VN_data_in(8677);
  VN1446_in2 <= VN_sign_in(8678) & VN_data_in(8678);
  VN1446_in3 <= VN_sign_in(8679) & VN_data_in(8679);
  VN1446_in4 <= VN_sign_in(8680) & VN_data_in(8680);
  VN1446_in5 <= VN_sign_in(8681) & VN_data_in(8681);
  VN1447_in0 <= VN_sign_in(8682) & VN_data_in(8682);
  VN1447_in1 <= VN_sign_in(8683) & VN_data_in(8683);
  VN1447_in2 <= VN_sign_in(8684) & VN_data_in(8684);
  VN1447_in3 <= VN_sign_in(8685) & VN_data_in(8685);
  VN1447_in4 <= VN_sign_in(8686) & VN_data_in(8686);
  VN1447_in5 <= VN_sign_in(8687) & VN_data_in(8687);
  VN1448_in0 <= VN_sign_in(8688) & VN_data_in(8688);
  VN1448_in1 <= VN_sign_in(8689) & VN_data_in(8689);
  VN1448_in2 <= VN_sign_in(8690) & VN_data_in(8690);
  VN1448_in3 <= VN_sign_in(8691) & VN_data_in(8691);
  VN1448_in4 <= VN_sign_in(8692) & VN_data_in(8692);
  VN1448_in5 <= VN_sign_in(8693) & VN_data_in(8693);
  VN1449_in0 <= VN_sign_in(8694) & VN_data_in(8694);
  VN1449_in1 <= VN_sign_in(8695) & VN_data_in(8695);
  VN1449_in2 <= VN_sign_in(8696) & VN_data_in(8696);
  VN1449_in3 <= VN_sign_in(8697) & VN_data_in(8697);
  VN1449_in4 <= VN_sign_in(8698) & VN_data_in(8698);
  VN1449_in5 <= VN_sign_in(8699) & VN_data_in(8699);
  VN1450_in0 <= VN_sign_in(8700) & VN_data_in(8700);
  VN1450_in1 <= VN_sign_in(8701) & VN_data_in(8701);
  VN1450_in2 <= VN_sign_in(8702) & VN_data_in(8702);
  VN1450_in3 <= VN_sign_in(8703) & VN_data_in(8703);
  VN1450_in4 <= VN_sign_in(8704) & VN_data_in(8704);
  VN1450_in5 <= VN_sign_in(8705) & VN_data_in(8705);
  VN1451_in0 <= VN_sign_in(8706) & VN_data_in(8706);
  VN1451_in1 <= VN_sign_in(8707) & VN_data_in(8707);
  VN1451_in2 <= VN_sign_in(8708) & VN_data_in(8708);
  VN1451_in3 <= VN_sign_in(8709) & VN_data_in(8709);
  VN1451_in4 <= VN_sign_in(8710) & VN_data_in(8710);
  VN1451_in5 <= VN_sign_in(8711) & VN_data_in(8711);
  VN1452_in0 <= VN_sign_in(8712) & VN_data_in(8712);
  VN1452_in1 <= VN_sign_in(8713) & VN_data_in(8713);
  VN1452_in2 <= VN_sign_in(8714) & VN_data_in(8714);
  VN1452_in3 <= VN_sign_in(8715) & VN_data_in(8715);
  VN1452_in4 <= VN_sign_in(8716) & VN_data_in(8716);
  VN1452_in5 <= VN_sign_in(8717) & VN_data_in(8717);
  VN1453_in0 <= VN_sign_in(8718) & VN_data_in(8718);
  VN1453_in1 <= VN_sign_in(8719) & VN_data_in(8719);
  VN1453_in2 <= VN_sign_in(8720) & VN_data_in(8720);
  VN1453_in3 <= VN_sign_in(8721) & VN_data_in(8721);
  VN1453_in4 <= VN_sign_in(8722) & VN_data_in(8722);
  VN1453_in5 <= VN_sign_in(8723) & VN_data_in(8723);
  VN1454_in0 <= VN_sign_in(8724) & VN_data_in(8724);
  VN1454_in1 <= VN_sign_in(8725) & VN_data_in(8725);
  VN1454_in2 <= VN_sign_in(8726) & VN_data_in(8726);
  VN1454_in3 <= VN_sign_in(8727) & VN_data_in(8727);
  VN1454_in4 <= VN_sign_in(8728) & VN_data_in(8728);
  VN1454_in5 <= VN_sign_in(8729) & VN_data_in(8729);
  VN1455_in0 <= VN_sign_in(8730) & VN_data_in(8730);
  VN1455_in1 <= VN_sign_in(8731) & VN_data_in(8731);
  VN1455_in2 <= VN_sign_in(8732) & VN_data_in(8732);
  VN1455_in3 <= VN_sign_in(8733) & VN_data_in(8733);
  VN1455_in4 <= VN_sign_in(8734) & VN_data_in(8734);
  VN1455_in5 <= VN_sign_in(8735) & VN_data_in(8735);
  VN1456_in0 <= VN_sign_in(8736) & VN_data_in(8736);
  VN1456_in1 <= VN_sign_in(8737) & VN_data_in(8737);
  VN1456_in2 <= VN_sign_in(8738) & VN_data_in(8738);
  VN1456_in3 <= VN_sign_in(8739) & VN_data_in(8739);
  VN1456_in4 <= VN_sign_in(8740) & VN_data_in(8740);
  VN1456_in5 <= VN_sign_in(8741) & VN_data_in(8741);
  VN1457_in0 <= VN_sign_in(8742) & VN_data_in(8742);
  VN1457_in1 <= VN_sign_in(8743) & VN_data_in(8743);
  VN1457_in2 <= VN_sign_in(8744) & VN_data_in(8744);
  VN1457_in3 <= VN_sign_in(8745) & VN_data_in(8745);
  VN1457_in4 <= VN_sign_in(8746) & VN_data_in(8746);
  VN1457_in5 <= VN_sign_in(8747) & VN_data_in(8747);
  VN1458_in0 <= VN_sign_in(8748) & VN_data_in(8748);
  VN1458_in1 <= VN_sign_in(8749) & VN_data_in(8749);
  VN1458_in2 <= VN_sign_in(8750) & VN_data_in(8750);
  VN1458_in3 <= VN_sign_in(8751) & VN_data_in(8751);
  VN1458_in4 <= VN_sign_in(8752) & VN_data_in(8752);
  VN1458_in5 <= VN_sign_in(8753) & VN_data_in(8753);
  VN1459_in0 <= VN_sign_in(8754) & VN_data_in(8754);
  VN1459_in1 <= VN_sign_in(8755) & VN_data_in(8755);
  VN1459_in2 <= VN_sign_in(8756) & VN_data_in(8756);
  VN1459_in3 <= VN_sign_in(8757) & VN_data_in(8757);
  VN1459_in4 <= VN_sign_in(8758) & VN_data_in(8758);
  VN1459_in5 <= VN_sign_in(8759) & VN_data_in(8759);
  VN1460_in0 <= VN_sign_in(8760) & VN_data_in(8760);
  VN1460_in1 <= VN_sign_in(8761) & VN_data_in(8761);
  VN1460_in2 <= VN_sign_in(8762) & VN_data_in(8762);
  VN1460_in3 <= VN_sign_in(8763) & VN_data_in(8763);
  VN1460_in4 <= VN_sign_in(8764) & VN_data_in(8764);
  VN1460_in5 <= VN_sign_in(8765) & VN_data_in(8765);
  VN1461_in0 <= VN_sign_in(8766) & VN_data_in(8766);
  VN1461_in1 <= VN_sign_in(8767) & VN_data_in(8767);
  VN1461_in2 <= VN_sign_in(8768) & VN_data_in(8768);
  VN1461_in3 <= VN_sign_in(8769) & VN_data_in(8769);
  VN1461_in4 <= VN_sign_in(8770) & VN_data_in(8770);
  VN1461_in5 <= VN_sign_in(8771) & VN_data_in(8771);
  VN1462_in0 <= VN_sign_in(8772) & VN_data_in(8772);
  VN1462_in1 <= VN_sign_in(8773) & VN_data_in(8773);
  VN1462_in2 <= VN_sign_in(8774) & VN_data_in(8774);
  VN1462_in3 <= VN_sign_in(8775) & VN_data_in(8775);
  VN1462_in4 <= VN_sign_in(8776) & VN_data_in(8776);
  VN1462_in5 <= VN_sign_in(8777) & VN_data_in(8777);
  VN1463_in0 <= VN_sign_in(8778) & VN_data_in(8778);
  VN1463_in1 <= VN_sign_in(8779) & VN_data_in(8779);
  VN1463_in2 <= VN_sign_in(8780) & VN_data_in(8780);
  VN1463_in3 <= VN_sign_in(8781) & VN_data_in(8781);
  VN1463_in4 <= VN_sign_in(8782) & VN_data_in(8782);
  VN1463_in5 <= VN_sign_in(8783) & VN_data_in(8783);
  VN1464_in0 <= VN_sign_in(8784) & VN_data_in(8784);
  VN1464_in1 <= VN_sign_in(8785) & VN_data_in(8785);
  VN1464_in2 <= VN_sign_in(8786) & VN_data_in(8786);
  VN1464_in3 <= VN_sign_in(8787) & VN_data_in(8787);
  VN1464_in4 <= VN_sign_in(8788) & VN_data_in(8788);
  VN1464_in5 <= VN_sign_in(8789) & VN_data_in(8789);
  VN1465_in0 <= VN_sign_in(8790) & VN_data_in(8790);
  VN1465_in1 <= VN_sign_in(8791) & VN_data_in(8791);
  VN1465_in2 <= VN_sign_in(8792) & VN_data_in(8792);
  VN1465_in3 <= VN_sign_in(8793) & VN_data_in(8793);
  VN1465_in4 <= VN_sign_in(8794) & VN_data_in(8794);
  VN1465_in5 <= VN_sign_in(8795) & VN_data_in(8795);
  VN1466_in0 <= VN_sign_in(8796) & VN_data_in(8796);
  VN1466_in1 <= VN_sign_in(8797) & VN_data_in(8797);
  VN1466_in2 <= VN_sign_in(8798) & VN_data_in(8798);
  VN1466_in3 <= VN_sign_in(8799) & VN_data_in(8799);
  VN1466_in4 <= VN_sign_in(8800) & VN_data_in(8800);
  VN1466_in5 <= VN_sign_in(8801) & VN_data_in(8801);
  VN1467_in0 <= VN_sign_in(8802) & VN_data_in(8802);
  VN1467_in1 <= VN_sign_in(8803) & VN_data_in(8803);
  VN1467_in2 <= VN_sign_in(8804) & VN_data_in(8804);
  VN1467_in3 <= VN_sign_in(8805) & VN_data_in(8805);
  VN1467_in4 <= VN_sign_in(8806) & VN_data_in(8806);
  VN1467_in5 <= VN_sign_in(8807) & VN_data_in(8807);
  VN1468_in0 <= VN_sign_in(8808) & VN_data_in(8808);
  VN1468_in1 <= VN_sign_in(8809) & VN_data_in(8809);
  VN1468_in2 <= VN_sign_in(8810) & VN_data_in(8810);
  VN1468_in3 <= VN_sign_in(8811) & VN_data_in(8811);
  VN1468_in4 <= VN_sign_in(8812) & VN_data_in(8812);
  VN1468_in5 <= VN_sign_in(8813) & VN_data_in(8813);
  VN1469_in0 <= VN_sign_in(8814) & VN_data_in(8814);
  VN1469_in1 <= VN_sign_in(8815) & VN_data_in(8815);
  VN1469_in2 <= VN_sign_in(8816) & VN_data_in(8816);
  VN1469_in3 <= VN_sign_in(8817) & VN_data_in(8817);
  VN1469_in4 <= VN_sign_in(8818) & VN_data_in(8818);
  VN1469_in5 <= VN_sign_in(8819) & VN_data_in(8819);
  VN1470_in0 <= VN_sign_in(8820) & VN_data_in(8820);
  VN1470_in1 <= VN_sign_in(8821) & VN_data_in(8821);
  VN1470_in2 <= VN_sign_in(8822) & VN_data_in(8822);
  VN1470_in3 <= VN_sign_in(8823) & VN_data_in(8823);
  VN1470_in4 <= VN_sign_in(8824) & VN_data_in(8824);
  VN1470_in5 <= VN_sign_in(8825) & VN_data_in(8825);
  VN1471_in0 <= VN_sign_in(8826) & VN_data_in(8826);
  VN1471_in1 <= VN_sign_in(8827) & VN_data_in(8827);
  VN1471_in2 <= VN_sign_in(8828) & VN_data_in(8828);
  VN1471_in3 <= VN_sign_in(8829) & VN_data_in(8829);
  VN1471_in4 <= VN_sign_in(8830) & VN_data_in(8830);
  VN1471_in5 <= VN_sign_in(8831) & VN_data_in(8831);
  VN1472_in0 <= VN_sign_in(8832) & VN_data_in(8832);
  VN1472_in1 <= VN_sign_in(8833) & VN_data_in(8833);
  VN1472_in2 <= VN_sign_in(8834) & VN_data_in(8834);
  VN1472_in3 <= VN_sign_in(8835) & VN_data_in(8835);
  VN1472_in4 <= VN_sign_in(8836) & VN_data_in(8836);
  VN1472_in5 <= VN_sign_in(8837) & VN_data_in(8837);
  VN1473_in0 <= VN_sign_in(8838) & VN_data_in(8838);
  VN1473_in1 <= VN_sign_in(8839) & VN_data_in(8839);
  VN1473_in2 <= VN_sign_in(8840) & VN_data_in(8840);
  VN1473_in3 <= VN_sign_in(8841) & VN_data_in(8841);
  VN1473_in4 <= VN_sign_in(8842) & VN_data_in(8842);
  VN1473_in5 <= VN_sign_in(8843) & VN_data_in(8843);
  VN1474_in0 <= VN_sign_in(8844) & VN_data_in(8844);
  VN1474_in1 <= VN_sign_in(8845) & VN_data_in(8845);
  VN1474_in2 <= VN_sign_in(8846) & VN_data_in(8846);
  VN1474_in3 <= VN_sign_in(8847) & VN_data_in(8847);
  VN1474_in4 <= VN_sign_in(8848) & VN_data_in(8848);
  VN1474_in5 <= VN_sign_in(8849) & VN_data_in(8849);
  VN1475_in0 <= VN_sign_in(8850) & VN_data_in(8850);
  VN1475_in1 <= VN_sign_in(8851) & VN_data_in(8851);
  VN1475_in2 <= VN_sign_in(8852) & VN_data_in(8852);
  VN1475_in3 <= VN_sign_in(8853) & VN_data_in(8853);
  VN1475_in4 <= VN_sign_in(8854) & VN_data_in(8854);
  VN1475_in5 <= VN_sign_in(8855) & VN_data_in(8855);
  VN1476_in0 <= VN_sign_in(8856) & VN_data_in(8856);
  VN1476_in1 <= VN_sign_in(8857) & VN_data_in(8857);
  VN1476_in2 <= VN_sign_in(8858) & VN_data_in(8858);
  VN1476_in3 <= VN_sign_in(8859) & VN_data_in(8859);
  VN1476_in4 <= VN_sign_in(8860) & VN_data_in(8860);
  VN1476_in5 <= VN_sign_in(8861) & VN_data_in(8861);
  VN1477_in0 <= VN_sign_in(8862) & VN_data_in(8862);
  VN1477_in1 <= VN_sign_in(8863) & VN_data_in(8863);
  VN1477_in2 <= VN_sign_in(8864) & VN_data_in(8864);
  VN1477_in3 <= VN_sign_in(8865) & VN_data_in(8865);
  VN1477_in4 <= VN_sign_in(8866) & VN_data_in(8866);
  VN1477_in5 <= VN_sign_in(8867) & VN_data_in(8867);
  VN1478_in0 <= VN_sign_in(8868) & VN_data_in(8868);
  VN1478_in1 <= VN_sign_in(8869) & VN_data_in(8869);
  VN1478_in2 <= VN_sign_in(8870) & VN_data_in(8870);
  VN1478_in3 <= VN_sign_in(8871) & VN_data_in(8871);
  VN1478_in4 <= VN_sign_in(8872) & VN_data_in(8872);
  VN1478_in5 <= VN_sign_in(8873) & VN_data_in(8873);
  VN1479_in0 <= VN_sign_in(8874) & VN_data_in(8874);
  VN1479_in1 <= VN_sign_in(8875) & VN_data_in(8875);
  VN1479_in2 <= VN_sign_in(8876) & VN_data_in(8876);
  VN1479_in3 <= VN_sign_in(8877) & VN_data_in(8877);
  VN1479_in4 <= VN_sign_in(8878) & VN_data_in(8878);
  VN1479_in5 <= VN_sign_in(8879) & VN_data_in(8879);
  VN1480_in0 <= VN_sign_in(8880) & VN_data_in(8880);
  VN1480_in1 <= VN_sign_in(8881) & VN_data_in(8881);
  VN1480_in2 <= VN_sign_in(8882) & VN_data_in(8882);
  VN1480_in3 <= VN_sign_in(8883) & VN_data_in(8883);
  VN1480_in4 <= VN_sign_in(8884) & VN_data_in(8884);
  VN1480_in5 <= VN_sign_in(8885) & VN_data_in(8885);
  VN1481_in0 <= VN_sign_in(8886) & VN_data_in(8886);
  VN1481_in1 <= VN_sign_in(8887) & VN_data_in(8887);
  VN1481_in2 <= VN_sign_in(8888) & VN_data_in(8888);
  VN1481_in3 <= VN_sign_in(8889) & VN_data_in(8889);
  VN1481_in4 <= VN_sign_in(8890) & VN_data_in(8890);
  VN1481_in5 <= VN_sign_in(8891) & VN_data_in(8891);
  VN1482_in0 <= VN_sign_in(8892) & VN_data_in(8892);
  VN1482_in1 <= VN_sign_in(8893) & VN_data_in(8893);
  VN1482_in2 <= VN_sign_in(8894) & VN_data_in(8894);
  VN1482_in3 <= VN_sign_in(8895) & VN_data_in(8895);
  VN1482_in4 <= VN_sign_in(8896) & VN_data_in(8896);
  VN1482_in5 <= VN_sign_in(8897) & VN_data_in(8897);
  VN1483_in0 <= VN_sign_in(8898) & VN_data_in(8898);
  VN1483_in1 <= VN_sign_in(8899) & VN_data_in(8899);
  VN1483_in2 <= VN_sign_in(8900) & VN_data_in(8900);
  VN1483_in3 <= VN_sign_in(8901) & VN_data_in(8901);
  VN1483_in4 <= VN_sign_in(8902) & VN_data_in(8902);
  VN1483_in5 <= VN_sign_in(8903) & VN_data_in(8903);
  VN1484_in0 <= VN_sign_in(8904) & VN_data_in(8904);
  VN1484_in1 <= VN_sign_in(8905) & VN_data_in(8905);
  VN1484_in2 <= VN_sign_in(8906) & VN_data_in(8906);
  VN1484_in3 <= VN_sign_in(8907) & VN_data_in(8907);
  VN1484_in4 <= VN_sign_in(8908) & VN_data_in(8908);
  VN1484_in5 <= VN_sign_in(8909) & VN_data_in(8909);
  VN1485_in0 <= VN_sign_in(8910) & VN_data_in(8910);
  VN1485_in1 <= VN_sign_in(8911) & VN_data_in(8911);
  VN1485_in2 <= VN_sign_in(8912) & VN_data_in(8912);
  VN1485_in3 <= VN_sign_in(8913) & VN_data_in(8913);
  VN1485_in4 <= VN_sign_in(8914) & VN_data_in(8914);
  VN1485_in5 <= VN_sign_in(8915) & VN_data_in(8915);
  VN1486_in0 <= VN_sign_in(8916) & VN_data_in(8916);
  VN1486_in1 <= VN_sign_in(8917) & VN_data_in(8917);
  VN1486_in2 <= VN_sign_in(8918) & VN_data_in(8918);
  VN1486_in3 <= VN_sign_in(8919) & VN_data_in(8919);
  VN1486_in4 <= VN_sign_in(8920) & VN_data_in(8920);
  VN1486_in5 <= VN_sign_in(8921) & VN_data_in(8921);
  VN1487_in0 <= VN_sign_in(8922) & VN_data_in(8922);
  VN1487_in1 <= VN_sign_in(8923) & VN_data_in(8923);
  VN1487_in2 <= VN_sign_in(8924) & VN_data_in(8924);
  VN1487_in3 <= VN_sign_in(8925) & VN_data_in(8925);
  VN1487_in4 <= VN_sign_in(8926) & VN_data_in(8926);
  VN1487_in5 <= VN_sign_in(8927) & VN_data_in(8927);
  VN1488_in0 <= VN_sign_in(8928) & VN_data_in(8928);
  VN1488_in1 <= VN_sign_in(8929) & VN_data_in(8929);
  VN1488_in2 <= VN_sign_in(8930) & VN_data_in(8930);
  VN1488_in3 <= VN_sign_in(8931) & VN_data_in(8931);
  VN1488_in4 <= VN_sign_in(8932) & VN_data_in(8932);
  VN1488_in5 <= VN_sign_in(8933) & VN_data_in(8933);
  VN1489_in0 <= VN_sign_in(8934) & VN_data_in(8934);
  VN1489_in1 <= VN_sign_in(8935) & VN_data_in(8935);
  VN1489_in2 <= VN_sign_in(8936) & VN_data_in(8936);
  VN1489_in3 <= VN_sign_in(8937) & VN_data_in(8937);
  VN1489_in4 <= VN_sign_in(8938) & VN_data_in(8938);
  VN1489_in5 <= VN_sign_in(8939) & VN_data_in(8939);
  VN1490_in0 <= VN_sign_in(8940) & VN_data_in(8940);
  VN1490_in1 <= VN_sign_in(8941) & VN_data_in(8941);
  VN1490_in2 <= VN_sign_in(8942) & VN_data_in(8942);
  VN1490_in3 <= VN_sign_in(8943) & VN_data_in(8943);
  VN1490_in4 <= VN_sign_in(8944) & VN_data_in(8944);
  VN1490_in5 <= VN_sign_in(8945) & VN_data_in(8945);
  VN1491_in0 <= VN_sign_in(8946) & VN_data_in(8946);
  VN1491_in1 <= VN_sign_in(8947) & VN_data_in(8947);
  VN1491_in2 <= VN_sign_in(8948) & VN_data_in(8948);
  VN1491_in3 <= VN_sign_in(8949) & VN_data_in(8949);
  VN1491_in4 <= VN_sign_in(8950) & VN_data_in(8950);
  VN1491_in5 <= VN_sign_in(8951) & VN_data_in(8951);
  VN1492_in0 <= VN_sign_in(8952) & VN_data_in(8952);
  VN1492_in1 <= VN_sign_in(8953) & VN_data_in(8953);
  VN1492_in2 <= VN_sign_in(8954) & VN_data_in(8954);
  VN1492_in3 <= VN_sign_in(8955) & VN_data_in(8955);
  VN1492_in4 <= VN_sign_in(8956) & VN_data_in(8956);
  VN1492_in5 <= VN_sign_in(8957) & VN_data_in(8957);
  VN1493_in0 <= VN_sign_in(8958) & VN_data_in(8958);
  VN1493_in1 <= VN_sign_in(8959) & VN_data_in(8959);
  VN1493_in2 <= VN_sign_in(8960) & VN_data_in(8960);
  VN1493_in3 <= VN_sign_in(8961) & VN_data_in(8961);
  VN1493_in4 <= VN_sign_in(8962) & VN_data_in(8962);
  VN1493_in5 <= VN_sign_in(8963) & VN_data_in(8963);
  VN1494_in0 <= VN_sign_in(8964) & VN_data_in(8964);
  VN1494_in1 <= VN_sign_in(8965) & VN_data_in(8965);
  VN1494_in2 <= VN_sign_in(8966) & VN_data_in(8966);
  VN1494_in3 <= VN_sign_in(8967) & VN_data_in(8967);
  VN1494_in4 <= VN_sign_in(8968) & VN_data_in(8968);
  VN1494_in5 <= VN_sign_in(8969) & VN_data_in(8969);
  VN1495_in0 <= VN_sign_in(8970) & VN_data_in(8970);
  VN1495_in1 <= VN_sign_in(8971) & VN_data_in(8971);
  VN1495_in2 <= VN_sign_in(8972) & VN_data_in(8972);
  VN1495_in3 <= VN_sign_in(8973) & VN_data_in(8973);
  VN1495_in4 <= VN_sign_in(8974) & VN_data_in(8974);
  VN1495_in5 <= VN_sign_in(8975) & VN_data_in(8975);
  VN1496_in0 <= VN_sign_in(8976) & VN_data_in(8976);
  VN1496_in1 <= VN_sign_in(8977) & VN_data_in(8977);
  VN1496_in2 <= VN_sign_in(8978) & VN_data_in(8978);
  VN1496_in3 <= VN_sign_in(8979) & VN_data_in(8979);
  VN1496_in4 <= VN_sign_in(8980) & VN_data_in(8980);
  VN1496_in5 <= VN_sign_in(8981) & VN_data_in(8981);
  VN1497_in0 <= VN_sign_in(8982) & VN_data_in(8982);
  VN1497_in1 <= VN_sign_in(8983) & VN_data_in(8983);
  VN1497_in2 <= VN_sign_in(8984) & VN_data_in(8984);
  VN1497_in3 <= VN_sign_in(8985) & VN_data_in(8985);
  VN1497_in4 <= VN_sign_in(8986) & VN_data_in(8986);
  VN1497_in5 <= VN_sign_in(8987) & VN_data_in(8987);
  VN1498_in0 <= VN_sign_in(8988) & VN_data_in(8988);
  VN1498_in1 <= VN_sign_in(8989) & VN_data_in(8989);
  VN1498_in2 <= VN_sign_in(8990) & VN_data_in(8990);
  VN1498_in3 <= VN_sign_in(8991) & VN_data_in(8991);
  VN1498_in4 <= VN_sign_in(8992) & VN_data_in(8992);
  VN1498_in5 <= VN_sign_in(8993) & VN_data_in(8993);
  VN1499_in0 <= VN_sign_in(8994) & VN_data_in(8994);
  VN1499_in1 <= VN_sign_in(8995) & VN_data_in(8995);
  VN1499_in2 <= VN_sign_in(8996) & VN_data_in(8996);
  VN1499_in3 <= VN_sign_in(8997) & VN_data_in(8997);
  VN1499_in4 <= VN_sign_in(8998) & VN_data_in(8998);
  VN1499_in5 <= VN_sign_in(8999) & VN_data_in(8999);
  VN1500_in0 <= VN_sign_in(9000) & VN_data_in(9000);
  VN1500_in1 <= VN_sign_in(9001) & VN_data_in(9001);
  VN1500_in2 <= VN_sign_in(9002) & VN_data_in(9002);
  VN1500_in3 <= VN_sign_in(9003) & VN_data_in(9003);
  VN1500_in4 <= VN_sign_in(9004) & VN_data_in(9004);
  VN1500_in5 <= VN_sign_in(9005) & VN_data_in(9005);
  VN1501_in0 <= VN_sign_in(9006) & VN_data_in(9006);
  VN1501_in1 <= VN_sign_in(9007) & VN_data_in(9007);
  VN1501_in2 <= VN_sign_in(9008) & VN_data_in(9008);
  VN1501_in3 <= VN_sign_in(9009) & VN_data_in(9009);
  VN1501_in4 <= VN_sign_in(9010) & VN_data_in(9010);
  VN1501_in5 <= VN_sign_in(9011) & VN_data_in(9011);
  VN1502_in0 <= VN_sign_in(9012) & VN_data_in(9012);
  VN1502_in1 <= VN_sign_in(9013) & VN_data_in(9013);
  VN1502_in2 <= VN_sign_in(9014) & VN_data_in(9014);
  VN1502_in3 <= VN_sign_in(9015) & VN_data_in(9015);
  VN1502_in4 <= VN_sign_in(9016) & VN_data_in(9016);
  VN1502_in5 <= VN_sign_in(9017) & VN_data_in(9017);
  VN1503_in0 <= VN_sign_in(9018) & VN_data_in(9018);
  VN1503_in1 <= VN_sign_in(9019) & VN_data_in(9019);
  VN1503_in2 <= VN_sign_in(9020) & VN_data_in(9020);
  VN1503_in3 <= VN_sign_in(9021) & VN_data_in(9021);
  VN1503_in4 <= VN_sign_in(9022) & VN_data_in(9022);
  VN1503_in5 <= VN_sign_in(9023) & VN_data_in(9023);
  VN1504_in0 <= VN_sign_in(9024) & VN_data_in(9024);
  VN1504_in1 <= VN_sign_in(9025) & VN_data_in(9025);
  VN1504_in2 <= VN_sign_in(9026) & VN_data_in(9026);
  VN1504_in3 <= VN_sign_in(9027) & VN_data_in(9027);
  VN1504_in4 <= VN_sign_in(9028) & VN_data_in(9028);
  VN1504_in5 <= VN_sign_in(9029) & VN_data_in(9029);
  VN1505_in0 <= VN_sign_in(9030) & VN_data_in(9030);
  VN1505_in1 <= VN_sign_in(9031) & VN_data_in(9031);
  VN1505_in2 <= VN_sign_in(9032) & VN_data_in(9032);
  VN1505_in3 <= VN_sign_in(9033) & VN_data_in(9033);
  VN1505_in4 <= VN_sign_in(9034) & VN_data_in(9034);
  VN1505_in5 <= VN_sign_in(9035) & VN_data_in(9035);
  VN1506_in0 <= VN_sign_in(9036) & VN_data_in(9036);
  VN1506_in1 <= VN_sign_in(9037) & VN_data_in(9037);
  VN1506_in2 <= VN_sign_in(9038) & VN_data_in(9038);
  VN1506_in3 <= VN_sign_in(9039) & VN_data_in(9039);
  VN1506_in4 <= VN_sign_in(9040) & VN_data_in(9040);
  VN1506_in5 <= VN_sign_in(9041) & VN_data_in(9041);
  VN1507_in0 <= VN_sign_in(9042) & VN_data_in(9042);
  VN1507_in1 <= VN_sign_in(9043) & VN_data_in(9043);
  VN1507_in2 <= VN_sign_in(9044) & VN_data_in(9044);
  VN1507_in3 <= VN_sign_in(9045) & VN_data_in(9045);
  VN1507_in4 <= VN_sign_in(9046) & VN_data_in(9046);
  VN1507_in5 <= VN_sign_in(9047) & VN_data_in(9047);
  VN1508_in0 <= VN_sign_in(9048) & VN_data_in(9048);
  VN1508_in1 <= VN_sign_in(9049) & VN_data_in(9049);
  VN1508_in2 <= VN_sign_in(9050) & VN_data_in(9050);
  VN1508_in3 <= VN_sign_in(9051) & VN_data_in(9051);
  VN1508_in4 <= VN_sign_in(9052) & VN_data_in(9052);
  VN1508_in5 <= VN_sign_in(9053) & VN_data_in(9053);
  VN1509_in0 <= VN_sign_in(9054) & VN_data_in(9054);
  VN1509_in1 <= VN_sign_in(9055) & VN_data_in(9055);
  VN1509_in2 <= VN_sign_in(9056) & VN_data_in(9056);
  VN1509_in3 <= VN_sign_in(9057) & VN_data_in(9057);
  VN1509_in4 <= VN_sign_in(9058) & VN_data_in(9058);
  VN1509_in5 <= VN_sign_in(9059) & VN_data_in(9059);
  VN1510_in0 <= VN_sign_in(9060) & VN_data_in(9060);
  VN1510_in1 <= VN_sign_in(9061) & VN_data_in(9061);
  VN1510_in2 <= VN_sign_in(9062) & VN_data_in(9062);
  VN1510_in3 <= VN_sign_in(9063) & VN_data_in(9063);
  VN1510_in4 <= VN_sign_in(9064) & VN_data_in(9064);
  VN1510_in5 <= VN_sign_in(9065) & VN_data_in(9065);
  VN1511_in0 <= VN_sign_in(9066) & VN_data_in(9066);
  VN1511_in1 <= VN_sign_in(9067) & VN_data_in(9067);
  VN1511_in2 <= VN_sign_in(9068) & VN_data_in(9068);
  VN1511_in3 <= VN_sign_in(9069) & VN_data_in(9069);
  VN1511_in4 <= VN_sign_in(9070) & VN_data_in(9070);
  VN1511_in5 <= VN_sign_in(9071) & VN_data_in(9071);
  VN1512_in0 <= VN_sign_in(9072) & VN_data_in(9072);
  VN1512_in1 <= VN_sign_in(9073) & VN_data_in(9073);
  VN1512_in2 <= VN_sign_in(9074) & VN_data_in(9074);
  VN1512_in3 <= VN_sign_in(9075) & VN_data_in(9075);
  VN1512_in4 <= VN_sign_in(9076) & VN_data_in(9076);
  VN1512_in5 <= VN_sign_in(9077) & VN_data_in(9077);
  VN1513_in0 <= VN_sign_in(9078) & VN_data_in(9078);
  VN1513_in1 <= VN_sign_in(9079) & VN_data_in(9079);
  VN1513_in2 <= VN_sign_in(9080) & VN_data_in(9080);
  VN1513_in3 <= VN_sign_in(9081) & VN_data_in(9081);
  VN1513_in4 <= VN_sign_in(9082) & VN_data_in(9082);
  VN1513_in5 <= VN_sign_in(9083) & VN_data_in(9083);
  VN1514_in0 <= VN_sign_in(9084) & VN_data_in(9084);
  VN1514_in1 <= VN_sign_in(9085) & VN_data_in(9085);
  VN1514_in2 <= VN_sign_in(9086) & VN_data_in(9086);
  VN1514_in3 <= VN_sign_in(9087) & VN_data_in(9087);
  VN1514_in4 <= VN_sign_in(9088) & VN_data_in(9088);
  VN1514_in5 <= VN_sign_in(9089) & VN_data_in(9089);
  VN1515_in0 <= VN_sign_in(9090) & VN_data_in(9090);
  VN1515_in1 <= VN_sign_in(9091) & VN_data_in(9091);
  VN1515_in2 <= VN_sign_in(9092) & VN_data_in(9092);
  VN1515_in3 <= VN_sign_in(9093) & VN_data_in(9093);
  VN1515_in4 <= VN_sign_in(9094) & VN_data_in(9094);
  VN1515_in5 <= VN_sign_in(9095) & VN_data_in(9095);
  VN1516_in0 <= VN_sign_in(9096) & VN_data_in(9096);
  VN1516_in1 <= VN_sign_in(9097) & VN_data_in(9097);
  VN1516_in2 <= VN_sign_in(9098) & VN_data_in(9098);
  VN1516_in3 <= VN_sign_in(9099) & VN_data_in(9099);
  VN1516_in4 <= VN_sign_in(9100) & VN_data_in(9100);
  VN1516_in5 <= VN_sign_in(9101) & VN_data_in(9101);
  VN1517_in0 <= VN_sign_in(9102) & VN_data_in(9102);
  VN1517_in1 <= VN_sign_in(9103) & VN_data_in(9103);
  VN1517_in2 <= VN_sign_in(9104) & VN_data_in(9104);
  VN1517_in3 <= VN_sign_in(9105) & VN_data_in(9105);
  VN1517_in4 <= VN_sign_in(9106) & VN_data_in(9106);
  VN1517_in5 <= VN_sign_in(9107) & VN_data_in(9107);
  VN1518_in0 <= VN_sign_in(9108) & VN_data_in(9108);
  VN1518_in1 <= VN_sign_in(9109) & VN_data_in(9109);
  VN1518_in2 <= VN_sign_in(9110) & VN_data_in(9110);
  VN1518_in3 <= VN_sign_in(9111) & VN_data_in(9111);
  VN1518_in4 <= VN_sign_in(9112) & VN_data_in(9112);
  VN1518_in5 <= VN_sign_in(9113) & VN_data_in(9113);
  VN1519_in0 <= VN_sign_in(9114) & VN_data_in(9114);
  VN1519_in1 <= VN_sign_in(9115) & VN_data_in(9115);
  VN1519_in2 <= VN_sign_in(9116) & VN_data_in(9116);
  VN1519_in3 <= VN_sign_in(9117) & VN_data_in(9117);
  VN1519_in4 <= VN_sign_in(9118) & VN_data_in(9118);
  VN1519_in5 <= VN_sign_in(9119) & VN_data_in(9119);
  VN1520_in0 <= VN_sign_in(9120) & VN_data_in(9120);
  VN1520_in1 <= VN_sign_in(9121) & VN_data_in(9121);
  VN1520_in2 <= VN_sign_in(9122) & VN_data_in(9122);
  VN1520_in3 <= VN_sign_in(9123) & VN_data_in(9123);
  VN1520_in4 <= VN_sign_in(9124) & VN_data_in(9124);
  VN1520_in5 <= VN_sign_in(9125) & VN_data_in(9125);
  VN1521_in0 <= VN_sign_in(9126) & VN_data_in(9126);
  VN1521_in1 <= VN_sign_in(9127) & VN_data_in(9127);
  VN1521_in2 <= VN_sign_in(9128) & VN_data_in(9128);
  VN1521_in3 <= VN_sign_in(9129) & VN_data_in(9129);
  VN1521_in4 <= VN_sign_in(9130) & VN_data_in(9130);
  VN1521_in5 <= VN_sign_in(9131) & VN_data_in(9131);
  VN1522_in0 <= VN_sign_in(9132) & VN_data_in(9132);
  VN1522_in1 <= VN_sign_in(9133) & VN_data_in(9133);
  VN1522_in2 <= VN_sign_in(9134) & VN_data_in(9134);
  VN1522_in3 <= VN_sign_in(9135) & VN_data_in(9135);
  VN1522_in4 <= VN_sign_in(9136) & VN_data_in(9136);
  VN1522_in5 <= VN_sign_in(9137) & VN_data_in(9137);
  VN1523_in0 <= VN_sign_in(9138) & VN_data_in(9138);
  VN1523_in1 <= VN_sign_in(9139) & VN_data_in(9139);
  VN1523_in2 <= VN_sign_in(9140) & VN_data_in(9140);
  VN1523_in3 <= VN_sign_in(9141) & VN_data_in(9141);
  VN1523_in4 <= VN_sign_in(9142) & VN_data_in(9142);
  VN1523_in5 <= VN_sign_in(9143) & VN_data_in(9143);
  VN1524_in0 <= VN_sign_in(9144) & VN_data_in(9144);
  VN1524_in1 <= VN_sign_in(9145) & VN_data_in(9145);
  VN1524_in2 <= VN_sign_in(9146) & VN_data_in(9146);
  VN1524_in3 <= VN_sign_in(9147) & VN_data_in(9147);
  VN1524_in4 <= VN_sign_in(9148) & VN_data_in(9148);
  VN1524_in5 <= VN_sign_in(9149) & VN_data_in(9149);
  VN1525_in0 <= VN_sign_in(9150) & VN_data_in(9150);
  VN1525_in1 <= VN_sign_in(9151) & VN_data_in(9151);
  VN1525_in2 <= VN_sign_in(9152) & VN_data_in(9152);
  VN1525_in3 <= VN_sign_in(9153) & VN_data_in(9153);
  VN1525_in4 <= VN_sign_in(9154) & VN_data_in(9154);
  VN1525_in5 <= VN_sign_in(9155) & VN_data_in(9155);
  VN1526_in0 <= VN_sign_in(9156) & VN_data_in(9156);
  VN1526_in1 <= VN_sign_in(9157) & VN_data_in(9157);
  VN1526_in2 <= VN_sign_in(9158) & VN_data_in(9158);
  VN1526_in3 <= VN_sign_in(9159) & VN_data_in(9159);
  VN1526_in4 <= VN_sign_in(9160) & VN_data_in(9160);
  VN1526_in5 <= VN_sign_in(9161) & VN_data_in(9161);
  VN1527_in0 <= VN_sign_in(9162) & VN_data_in(9162);
  VN1527_in1 <= VN_sign_in(9163) & VN_data_in(9163);
  VN1527_in2 <= VN_sign_in(9164) & VN_data_in(9164);
  VN1527_in3 <= VN_sign_in(9165) & VN_data_in(9165);
  VN1527_in4 <= VN_sign_in(9166) & VN_data_in(9166);
  VN1527_in5 <= VN_sign_in(9167) & VN_data_in(9167);
  VN1528_in0 <= VN_sign_in(9168) & VN_data_in(9168);
  VN1528_in1 <= VN_sign_in(9169) & VN_data_in(9169);
  VN1528_in2 <= VN_sign_in(9170) & VN_data_in(9170);
  VN1528_in3 <= VN_sign_in(9171) & VN_data_in(9171);
  VN1528_in4 <= VN_sign_in(9172) & VN_data_in(9172);
  VN1528_in5 <= VN_sign_in(9173) & VN_data_in(9173);
  VN1529_in0 <= VN_sign_in(9174) & VN_data_in(9174);
  VN1529_in1 <= VN_sign_in(9175) & VN_data_in(9175);
  VN1529_in2 <= VN_sign_in(9176) & VN_data_in(9176);
  VN1529_in3 <= VN_sign_in(9177) & VN_data_in(9177);
  VN1529_in4 <= VN_sign_in(9178) & VN_data_in(9178);
  VN1529_in5 <= VN_sign_in(9179) & VN_data_in(9179);
  VN1530_in0 <= VN_sign_in(9180) & VN_data_in(9180);
  VN1530_in1 <= VN_sign_in(9181) & VN_data_in(9181);
  VN1530_in2 <= VN_sign_in(9182) & VN_data_in(9182);
  VN1530_in3 <= VN_sign_in(9183) & VN_data_in(9183);
  VN1530_in4 <= VN_sign_in(9184) & VN_data_in(9184);
  VN1530_in5 <= VN_sign_in(9185) & VN_data_in(9185);
  VN1531_in0 <= VN_sign_in(9186) & VN_data_in(9186);
  VN1531_in1 <= VN_sign_in(9187) & VN_data_in(9187);
  VN1531_in2 <= VN_sign_in(9188) & VN_data_in(9188);
  VN1531_in3 <= VN_sign_in(9189) & VN_data_in(9189);
  VN1531_in4 <= VN_sign_in(9190) & VN_data_in(9190);
  VN1531_in5 <= VN_sign_in(9191) & VN_data_in(9191);
  VN1532_in0 <= VN_sign_in(9192) & VN_data_in(9192);
  VN1532_in1 <= VN_sign_in(9193) & VN_data_in(9193);
  VN1532_in2 <= VN_sign_in(9194) & VN_data_in(9194);
  VN1532_in3 <= VN_sign_in(9195) & VN_data_in(9195);
  VN1532_in4 <= VN_sign_in(9196) & VN_data_in(9196);
  VN1532_in5 <= VN_sign_in(9197) & VN_data_in(9197);
  VN1533_in0 <= VN_sign_in(9198) & VN_data_in(9198);
  VN1533_in1 <= VN_sign_in(9199) & VN_data_in(9199);
  VN1533_in2 <= VN_sign_in(9200) & VN_data_in(9200);
  VN1533_in3 <= VN_sign_in(9201) & VN_data_in(9201);
  VN1533_in4 <= VN_sign_in(9202) & VN_data_in(9202);
  VN1533_in5 <= VN_sign_in(9203) & VN_data_in(9203);
  VN1534_in0 <= VN_sign_in(9204) & VN_data_in(9204);
  VN1534_in1 <= VN_sign_in(9205) & VN_data_in(9205);
  VN1534_in2 <= VN_sign_in(9206) & VN_data_in(9206);
  VN1534_in3 <= VN_sign_in(9207) & VN_data_in(9207);
  VN1534_in4 <= VN_sign_in(9208) & VN_data_in(9208);
  VN1534_in5 <= VN_sign_in(9209) & VN_data_in(9209);
  VN1535_in0 <= VN_sign_in(9210) & VN_data_in(9210);
  VN1535_in1 <= VN_sign_in(9211) & VN_data_in(9211);
  VN1535_in2 <= VN_sign_in(9212) & VN_data_in(9212);
  VN1535_in3 <= VN_sign_in(9213) & VN_data_in(9213);
  VN1535_in4 <= VN_sign_in(9214) & VN_data_in(9214);
  VN1535_in5 <= VN_sign_in(9215) & VN_data_in(9215);
  VN1536_in0 <= VN_sign_in(9216) & VN_data_in(9216);
  VN1536_in1 <= VN_sign_in(9217) & VN_data_in(9217);
  VN1536_in2 <= VN_sign_in(9218) & VN_data_in(9218);
  VN1536_in3 <= VN_sign_in(9219) & VN_data_in(9219);
  VN1536_in4 <= VN_sign_in(9220) & VN_data_in(9220);
  VN1536_in5 <= VN_sign_in(9221) & VN_data_in(9221);
  VN1537_in0 <= VN_sign_in(9222) & VN_data_in(9222);
  VN1537_in1 <= VN_sign_in(9223) & VN_data_in(9223);
  VN1537_in2 <= VN_sign_in(9224) & VN_data_in(9224);
  VN1537_in3 <= VN_sign_in(9225) & VN_data_in(9225);
  VN1537_in4 <= VN_sign_in(9226) & VN_data_in(9226);
  VN1537_in5 <= VN_sign_in(9227) & VN_data_in(9227);
  VN1538_in0 <= VN_sign_in(9228) & VN_data_in(9228);
  VN1538_in1 <= VN_sign_in(9229) & VN_data_in(9229);
  VN1538_in2 <= VN_sign_in(9230) & VN_data_in(9230);
  VN1538_in3 <= VN_sign_in(9231) & VN_data_in(9231);
  VN1538_in4 <= VN_sign_in(9232) & VN_data_in(9232);
  VN1538_in5 <= VN_sign_in(9233) & VN_data_in(9233);
  VN1539_in0 <= VN_sign_in(9234) & VN_data_in(9234);
  VN1539_in1 <= VN_sign_in(9235) & VN_data_in(9235);
  VN1539_in2 <= VN_sign_in(9236) & VN_data_in(9236);
  VN1539_in3 <= VN_sign_in(9237) & VN_data_in(9237);
  VN1539_in4 <= VN_sign_in(9238) & VN_data_in(9238);
  VN1539_in5 <= VN_sign_in(9239) & VN_data_in(9239);
  VN1540_in0 <= VN_sign_in(9240) & VN_data_in(9240);
  VN1540_in1 <= VN_sign_in(9241) & VN_data_in(9241);
  VN1540_in2 <= VN_sign_in(9242) & VN_data_in(9242);
  VN1540_in3 <= VN_sign_in(9243) & VN_data_in(9243);
  VN1540_in4 <= VN_sign_in(9244) & VN_data_in(9244);
  VN1540_in5 <= VN_sign_in(9245) & VN_data_in(9245);
  VN1541_in0 <= VN_sign_in(9246) & VN_data_in(9246);
  VN1541_in1 <= VN_sign_in(9247) & VN_data_in(9247);
  VN1541_in2 <= VN_sign_in(9248) & VN_data_in(9248);
  VN1541_in3 <= VN_sign_in(9249) & VN_data_in(9249);
  VN1541_in4 <= VN_sign_in(9250) & VN_data_in(9250);
  VN1541_in5 <= VN_sign_in(9251) & VN_data_in(9251);
  VN1542_in0 <= VN_sign_in(9252) & VN_data_in(9252);
  VN1542_in1 <= VN_sign_in(9253) & VN_data_in(9253);
  VN1542_in2 <= VN_sign_in(9254) & VN_data_in(9254);
  VN1542_in3 <= VN_sign_in(9255) & VN_data_in(9255);
  VN1542_in4 <= VN_sign_in(9256) & VN_data_in(9256);
  VN1542_in5 <= VN_sign_in(9257) & VN_data_in(9257);
  VN1543_in0 <= VN_sign_in(9258) & VN_data_in(9258);
  VN1543_in1 <= VN_sign_in(9259) & VN_data_in(9259);
  VN1543_in2 <= VN_sign_in(9260) & VN_data_in(9260);
  VN1543_in3 <= VN_sign_in(9261) & VN_data_in(9261);
  VN1543_in4 <= VN_sign_in(9262) & VN_data_in(9262);
  VN1543_in5 <= VN_sign_in(9263) & VN_data_in(9263);
  VN1544_in0 <= VN_sign_in(9264) & VN_data_in(9264);
  VN1544_in1 <= VN_sign_in(9265) & VN_data_in(9265);
  VN1544_in2 <= VN_sign_in(9266) & VN_data_in(9266);
  VN1544_in3 <= VN_sign_in(9267) & VN_data_in(9267);
  VN1544_in4 <= VN_sign_in(9268) & VN_data_in(9268);
  VN1544_in5 <= VN_sign_in(9269) & VN_data_in(9269);
  VN1545_in0 <= VN_sign_in(9270) & VN_data_in(9270);
  VN1545_in1 <= VN_sign_in(9271) & VN_data_in(9271);
  VN1545_in2 <= VN_sign_in(9272) & VN_data_in(9272);
  VN1545_in3 <= VN_sign_in(9273) & VN_data_in(9273);
  VN1545_in4 <= VN_sign_in(9274) & VN_data_in(9274);
  VN1545_in5 <= VN_sign_in(9275) & VN_data_in(9275);
  VN1546_in0 <= VN_sign_in(9276) & VN_data_in(9276);
  VN1546_in1 <= VN_sign_in(9277) & VN_data_in(9277);
  VN1546_in2 <= VN_sign_in(9278) & VN_data_in(9278);
  VN1546_in3 <= VN_sign_in(9279) & VN_data_in(9279);
  VN1546_in4 <= VN_sign_in(9280) & VN_data_in(9280);
  VN1546_in5 <= VN_sign_in(9281) & VN_data_in(9281);
  VN1547_in0 <= VN_sign_in(9282) & VN_data_in(9282);
  VN1547_in1 <= VN_sign_in(9283) & VN_data_in(9283);
  VN1547_in2 <= VN_sign_in(9284) & VN_data_in(9284);
  VN1547_in3 <= VN_sign_in(9285) & VN_data_in(9285);
  VN1547_in4 <= VN_sign_in(9286) & VN_data_in(9286);
  VN1547_in5 <= VN_sign_in(9287) & VN_data_in(9287);
  VN1548_in0 <= VN_sign_in(9288) & VN_data_in(9288);
  VN1548_in1 <= VN_sign_in(9289) & VN_data_in(9289);
  VN1548_in2 <= VN_sign_in(9290) & VN_data_in(9290);
  VN1548_in3 <= VN_sign_in(9291) & VN_data_in(9291);
  VN1548_in4 <= VN_sign_in(9292) & VN_data_in(9292);
  VN1548_in5 <= VN_sign_in(9293) & VN_data_in(9293);
  VN1549_in0 <= VN_sign_in(9294) & VN_data_in(9294);
  VN1549_in1 <= VN_sign_in(9295) & VN_data_in(9295);
  VN1549_in2 <= VN_sign_in(9296) & VN_data_in(9296);
  VN1549_in3 <= VN_sign_in(9297) & VN_data_in(9297);
  VN1549_in4 <= VN_sign_in(9298) & VN_data_in(9298);
  VN1549_in5 <= VN_sign_in(9299) & VN_data_in(9299);
  VN1550_in0 <= VN_sign_in(9300) & VN_data_in(9300);
  VN1550_in1 <= VN_sign_in(9301) & VN_data_in(9301);
  VN1550_in2 <= VN_sign_in(9302) & VN_data_in(9302);
  VN1550_in3 <= VN_sign_in(9303) & VN_data_in(9303);
  VN1550_in4 <= VN_sign_in(9304) & VN_data_in(9304);
  VN1550_in5 <= VN_sign_in(9305) & VN_data_in(9305);
  VN1551_in0 <= VN_sign_in(9306) & VN_data_in(9306);
  VN1551_in1 <= VN_sign_in(9307) & VN_data_in(9307);
  VN1551_in2 <= VN_sign_in(9308) & VN_data_in(9308);
  VN1551_in3 <= VN_sign_in(9309) & VN_data_in(9309);
  VN1551_in4 <= VN_sign_in(9310) & VN_data_in(9310);
  VN1551_in5 <= VN_sign_in(9311) & VN_data_in(9311);
  VN1552_in0 <= VN_sign_in(9312) & VN_data_in(9312);
  VN1552_in1 <= VN_sign_in(9313) & VN_data_in(9313);
  VN1552_in2 <= VN_sign_in(9314) & VN_data_in(9314);
  VN1552_in3 <= VN_sign_in(9315) & VN_data_in(9315);
  VN1552_in4 <= VN_sign_in(9316) & VN_data_in(9316);
  VN1552_in5 <= VN_sign_in(9317) & VN_data_in(9317);
  VN1553_in0 <= VN_sign_in(9318) & VN_data_in(9318);
  VN1553_in1 <= VN_sign_in(9319) & VN_data_in(9319);
  VN1553_in2 <= VN_sign_in(9320) & VN_data_in(9320);
  VN1553_in3 <= VN_sign_in(9321) & VN_data_in(9321);
  VN1553_in4 <= VN_sign_in(9322) & VN_data_in(9322);
  VN1553_in5 <= VN_sign_in(9323) & VN_data_in(9323);
  VN1554_in0 <= VN_sign_in(9324) & VN_data_in(9324);
  VN1554_in1 <= VN_sign_in(9325) & VN_data_in(9325);
  VN1554_in2 <= VN_sign_in(9326) & VN_data_in(9326);
  VN1554_in3 <= VN_sign_in(9327) & VN_data_in(9327);
  VN1554_in4 <= VN_sign_in(9328) & VN_data_in(9328);
  VN1554_in5 <= VN_sign_in(9329) & VN_data_in(9329);
  VN1555_in0 <= VN_sign_in(9330) & VN_data_in(9330);
  VN1555_in1 <= VN_sign_in(9331) & VN_data_in(9331);
  VN1555_in2 <= VN_sign_in(9332) & VN_data_in(9332);
  VN1555_in3 <= VN_sign_in(9333) & VN_data_in(9333);
  VN1555_in4 <= VN_sign_in(9334) & VN_data_in(9334);
  VN1555_in5 <= VN_sign_in(9335) & VN_data_in(9335);
  VN1556_in0 <= VN_sign_in(9336) & VN_data_in(9336);
  VN1556_in1 <= VN_sign_in(9337) & VN_data_in(9337);
  VN1556_in2 <= VN_sign_in(9338) & VN_data_in(9338);
  VN1556_in3 <= VN_sign_in(9339) & VN_data_in(9339);
  VN1556_in4 <= VN_sign_in(9340) & VN_data_in(9340);
  VN1556_in5 <= VN_sign_in(9341) & VN_data_in(9341);
  VN1557_in0 <= VN_sign_in(9342) & VN_data_in(9342);
  VN1557_in1 <= VN_sign_in(9343) & VN_data_in(9343);
  VN1557_in2 <= VN_sign_in(9344) & VN_data_in(9344);
  VN1557_in3 <= VN_sign_in(9345) & VN_data_in(9345);
  VN1557_in4 <= VN_sign_in(9346) & VN_data_in(9346);
  VN1557_in5 <= VN_sign_in(9347) & VN_data_in(9347);
  VN1558_in0 <= VN_sign_in(9348) & VN_data_in(9348);
  VN1558_in1 <= VN_sign_in(9349) & VN_data_in(9349);
  VN1558_in2 <= VN_sign_in(9350) & VN_data_in(9350);
  VN1558_in3 <= VN_sign_in(9351) & VN_data_in(9351);
  VN1558_in4 <= VN_sign_in(9352) & VN_data_in(9352);
  VN1558_in5 <= VN_sign_in(9353) & VN_data_in(9353);
  VN1559_in0 <= VN_sign_in(9354) & VN_data_in(9354);
  VN1559_in1 <= VN_sign_in(9355) & VN_data_in(9355);
  VN1559_in2 <= VN_sign_in(9356) & VN_data_in(9356);
  VN1559_in3 <= VN_sign_in(9357) & VN_data_in(9357);
  VN1559_in4 <= VN_sign_in(9358) & VN_data_in(9358);
  VN1559_in5 <= VN_sign_in(9359) & VN_data_in(9359);
  VN1560_in0 <= VN_sign_in(9360) & VN_data_in(9360);
  VN1560_in1 <= VN_sign_in(9361) & VN_data_in(9361);
  VN1560_in2 <= VN_sign_in(9362) & VN_data_in(9362);
  VN1560_in3 <= VN_sign_in(9363) & VN_data_in(9363);
  VN1560_in4 <= VN_sign_in(9364) & VN_data_in(9364);
  VN1560_in5 <= VN_sign_in(9365) & VN_data_in(9365);
  VN1561_in0 <= VN_sign_in(9366) & VN_data_in(9366);
  VN1561_in1 <= VN_sign_in(9367) & VN_data_in(9367);
  VN1561_in2 <= VN_sign_in(9368) & VN_data_in(9368);
  VN1561_in3 <= VN_sign_in(9369) & VN_data_in(9369);
  VN1561_in4 <= VN_sign_in(9370) & VN_data_in(9370);
  VN1561_in5 <= VN_sign_in(9371) & VN_data_in(9371);
  VN1562_in0 <= VN_sign_in(9372) & VN_data_in(9372);
  VN1562_in1 <= VN_sign_in(9373) & VN_data_in(9373);
  VN1562_in2 <= VN_sign_in(9374) & VN_data_in(9374);
  VN1562_in3 <= VN_sign_in(9375) & VN_data_in(9375);
  VN1562_in4 <= VN_sign_in(9376) & VN_data_in(9376);
  VN1562_in5 <= VN_sign_in(9377) & VN_data_in(9377);
  VN1563_in0 <= VN_sign_in(9378) & VN_data_in(9378);
  VN1563_in1 <= VN_sign_in(9379) & VN_data_in(9379);
  VN1563_in2 <= VN_sign_in(9380) & VN_data_in(9380);
  VN1563_in3 <= VN_sign_in(9381) & VN_data_in(9381);
  VN1563_in4 <= VN_sign_in(9382) & VN_data_in(9382);
  VN1563_in5 <= VN_sign_in(9383) & VN_data_in(9383);
  VN1564_in0 <= VN_sign_in(9384) & VN_data_in(9384);
  VN1564_in1 <= VN_sign_in(9385) & VN_data_in(9385);
  VN1564_in2 <= VN_sign_in(9386) & VN_data_in(9386);
  VN1564_in3 <= VN_sign_in(9387) & VN_data_in(9387);
  VN1564_in4 <= VN_sign_in(9388) & VN_data_in(9388);
  VN1564_in5 <= VN_sign_in(9389) & VN_data_in(9389);
  VN1565_in0 <= VN_sign_in(9390) & VN_data_in(9390);
  VN1565_in1 <= VN_sign_in(9391) & VN_data_in(9391);
  VN1565_in2 <= VN_sign_in(9392) & VN_data_in(9392);
  VN1565_in3 <= VN_sign_in(9393) & VN_data_in(9393);
  VN1565_in4 <= VN_sign_in(9394) & VN_data_in(9394);
  VN1565_in5 <= VN_sign_in(9395) & VN_data_in(9395);
  VN1566_in0 <= VN_sign_in(9396) & VN_data_in(9396);
  VN1566_in1 <= VN_sign_in(9397) & VN_data_in(9397);
  VN1566_in2 <= VN_sign_in(9398) & VN_data_in(9398);
  VN1566_in3 <= VN_sign_in(9399) & VN_data_in(9399);
  VN1566_in4 <= VN_sign_in(9400) & VN_data_in(9400);
  VN1566_in5 <= VN_sign_in(9401) & VN_data_in(9401);
  VN1567_in0 <= VN_sign_in(9402) & VN_data_in(9402);
  VN1567_in1 <= VN_sign_in(9403) & VN_data_in(9403);
  VN1567_in2 <= VN_sign_in(9404) & VN_data_in(9404);
  VN1567_in3 <= VN_sign_in(9405) & VN_data_in(9405);
  VN1567_in4 <= VN_sign_in(9406) & VN_data_in(9406);
  VN1567_in5 <= VN_sign_in(9407) & VN_data_in(9407);
  VN1568_in0 <= VN_sign_in(9408) & VN_data_in(9408);
  VN1568_in1 <= VN_sign_in(9409) & VN_data_in(9409);
  VN1568_in2 <= VN_sign_in(9410) & VN_data_in(9410);
  VN1568_in3 <= VN_sign_in(9411) & VN_data_in(9411);
  VN1568_in4 <= VN_sign_in(9412) & VN_data_in(9412);
  VN1568_in5 <= VN_sign_in(9413) & VN_data_in(9413);
  VN1569_in0 <= VN_sign_in(9414) & VN_data_in(9414);
  VN1569_in1 <= VN_sign_in(9415) & VN_data_in(9415);
  VN1569_in2 <= VN_sign_in(9416) & VN_data_in(9416);
  VN1569_in3 <= VN_sign_in(9417) & VN_data_in(9417);
  VN1569_in4 <= VN_sign_in(9418) & VN_data_in(9418);
  VN1569_in5 <= VN_sign_in(9419) & VN_data_in(9419);
  VN1570_in0 <= VN_sign_in(9420) & VN_data_in(9420);
  VN1570_in1 <= VN_sign_in(9421) & VN_data_in(9421);
  VN1570_in2 <= VN_sign_in(9422) & VN_data_in(9422);
  VN1570_in3 <= VN_sign_in(9423) & VN_data_in(9423);
  VN1570_in4 <= VN_sign_in(9424) & VN_data_in(9424);
  VN1570_in5 <= VN_sign_in(9425) & VN_data_in(9425);
  VN1571_in0 <= VN_sign_in(9426) & VN_data_in(9426);
  VN1571_in1 <= VN_sign_in(9427) & VN_data_in(9427);
  VN1571_in2 <= VN_sign_in(9428) & VN_data_in(9428);
  VN1571_in3 <= VN_sign_in(9429) & VN_data_in(9429);
  VN1571_in4 <= VN_sign_in(9430) & VN_data_in(9430);
  VN1571_in5 <= VN_sign_in(9431) & VN_data_in(9431);
  VN1572_in0 <= VN_sign_in(9432) & VN_data_in(9432);
  VN1572_in1 <= VN_sign_in(9433) & VN_data_in(9433);
  VN1572_in2 <= VN_sign_in(9434) & VN_data_in(9434);
  VN1572_in3 <= VN_sign_in(9435) & VN_data_in(9435);
  VN1572_in4 <= VN_sign_in(9436) & VN_data_in(9436);
  VN1572_in5 <= VN_sign_in(9437) & VN_data_in(9437);
  VN1573_in0 <= VN_sign_in(9438) & VN_data_in(9438);
  VN1573_in1 <= VN_sign_in(9439) & VN_data_in(9439);
  VN1573_in2 <= VN_sign_in(9440) & VN_data_in(9440);
  VN1573_in3 <= VN_sign_in(9441) & VN_data_in(9441);
  VN1573_in4 <= VN_sign_in(9442) & VN_data_in(9442);
  VN1573_in5 <= VN_sign_in(9443) & VN_data_in(9443);
  VN1574_in0 <= VN_sign_in(9444) & VN_data_in(9444);
  VN1574_in1 <= VN_sign_in(9445) & VN_data_in(9445);
  VN1574_in2 <= VN_sign_in(9446) & VN_data_in(9446);
  VN1574_in3 <= VN_sign_in(9447) & VN_data_in(9447);
  VN1574_in4 <= VN_sign_in(9448) & VN_data_in(9448);
  VN1574_in5 <= VN_sign_in(9449) & VN_data_in(9449);
  VN1575_in0 <= VN_sign_in(9450) & VN_data_in(9450);
  VN1575_in1 <= VN_sign_in(9451) & VN_data_in(9451);
  VN1575_in2 <= VN_sign_in(9452) & VN_data_in(9452);
  VN1575_in3 <= VN_sign_in(9453) & VN_data_in(9453);
  VN1575_in4 <= VN_sign_in(9454) & VN_data_in(9454);
  VN1575_in5 <= VN_sign_in(9455) & VN_data_in(9455);
  VN1576_in0 <= VN_sign_in(9456) & VN_data_in(9456);
  VN1576_in1 <= VN_sign_in(9457) & VN_data_in(9457);
  VN1576_in2 <= VN_sign_in(9458) & VN_data_in(9458);
  VN1576_in3 <= VN_sign_in(9459) & VN_data_in(9459);
  VN1576_in4 <= VN_sign_in(9460) & VN_data_in(9460);
  VN1576_in5 <= VN_sign_in(9461) & VN_data_in(9461);
  VN1577_in0 <= VN_sign_in(9462) & VN_data_in(9462);
  VN1577_in1 <= VN_sign_in(9463) & VN_data_in(9463);
  VN1577_in2 <= VN_sign_in(9464) & VN_data_in(9464);
  VN1577_in3 <= VN_sign_in(9465) & VN_data_in(9465);
  VN1577_in4 <= VN_sign_in(9466) & VN_data_in(9466);
  VN1577_in5 <= VN_sign_in(9467) & VN_data_in(9467);
  VN1578_in0 <= VN_sign_in(9468) & VN_data_in(9468);
  VN1578_in1 <= VN_sign_in(9469) & VN_data_in(9469);
  VN1578_in2 <= VN_sign_in(9470) & VN_data_in(9470);
  VN1578_in3 <= VN_sign_in(9471) & VN_data_in(9471);
  VN1578_in4 <= VN_sign_in(9472) & VN_data_in(9472);
  VN1578_in5 <= VN_sign_in(9473) & VN_data_in(9473);
  VN1579_in0 <= VN_sign_in(9474) & VN_data_in(9474);
  VN1579_in1 <= VN_sign_in(9475) & VN_data_in(9475);
  VN1579_in2 <= VN_sign_in(9476) & VN_data_in(9476);
  VN1579_in3 <= VN_sign_in(9477) & VN_data_in(9477);
  VN1579_in4 <= VN_sign_in(9478) & VN_data_in(9478);
  VN1579_in5 <= VN_sign_in(9479) & VN_data_in(9479);
  VN1580_in0 <= VN_sign_in(9480) & VN_data_in(9480);
  VN1580_in1 <= VN_sign_in(9481) & VN_data_in(9481);
  VN1580_in2 <= VN_sign_in(9482) & VN_data_in(9482);
  VN1580_in3 <= VN_sign_in(9483) & VN_data_in(9483);
  VN1580_in4 <= VN_sign_in(9484) & VN_data_in(9484);
  VN1580_in5 <= VN_sign_in(9485) & VN_data_in(9485);
  VN1581_in0 <= VN_sign_in(9486) & VN_data_in(9486);
  VN1581_in1 <= VN_sign_in(9487) & VN_data_in(9487);
  VN1581_in2 <= VN_sign_in(9488) & VN_data_in(9488);
  VN1581_in3 <= VN_sign_in(9489) & VN_data_in(9489);
  VN1581_in4 <= VN_sign_in(9490) & VN_data_in(9490);
  VN1581_in5 <= VN_sign_in(9491) & VN_data_in(9491);
  VN1582_in0 <= VN_sign_in(9492) & VN_data_in(9492);
  VN1582_in1 <= VN_sign_in(9493) & VN_data_in(9493);
  VN1582_in2 <= VN_sign_in(9494) & VN_data_in(9494);
  VN1582_in3 <= VN_sign_in(9495) & VN_data_in(9495);
  VN1582_in4 <= VN_sign_in(9496) & VN_data_in(9496);
  VN1582_in5 <= VN_sign_in(9497) & VN_data_in(9497);
  VN1583_in0 <= VN_sign_in(9498) & VN_data_in(9498);
  VN1583_in1 <= VN_sign_in(9499) & VN_data_in(9499);
  VN1583_in2 <= VN_sign_in(9500) & VN_data_in(9500);
  VN1583_in3 <= VN_sign_in(9501) & VN_data_in(9501);
  VN1583_in4 <= VN_sign_in(9502) & VN_data_in(9502);
  VN1583_in5 <= VN_sign_in(9503) & VN_data_in(9503);
  VN1584_in0 <= VN_sign_in(9504) & VN_data_in(9504);
  VN1584_in1 <= VN_sign_in(9505) & VN_data_in(9505);
  VN1584_in2 <= VN_sign_in(9506) & VN_data_in(9506);
  VN1584_in3 <= VN_sign_in(9507) & VN_data_in(9507);
  VN1584_in4 <= VN_sign_in(9508) & VN_data_in(9508);
  VN1584_in5 <= VN_sign_in(9509) & VN_data_in(9509);
  VN1585_in0 <= VN_sign_in(9510) & VN_data_in(9510);
  VN1585_in1 <= VN_sign_in(9511) & VN_data_in(9511);
  VN1585_in2 <= VN_sign_in(9512) & VN_data_in(9512);
  VN1585_in3 <= VN_sign_in(9513) & VN_data_in(9513);
  VN1585_in4 <= VN_sign_in(9514) & VN_data_in(9514);
  VN1585_in5 <= VN_sign_in(9515) & VN_data_in(9515);
  VN1586_in0 <= VN_sign_in(9516) & VN_data_in(9516);
  VN1586_in1 <= VN_sign_in(9517) & VN_data_in(9517);
  VN1586_in2 <= VN_sign_in(9518) & VN_data_in(9518);
  VN1586_in3 <= VN_sign_in(9519) & VN_data_in(9519);
  VN1586_in4 <= VN_sign_in(9520) & VN_data_in(9520);
  VN1586_in5 <= VN_sign_in(9521) & VN_data_in(9521);
  VN1587_in0 <= VN_sign_in(9522) & VN_data_in(9522);
  VN1587_in1 <= VN_sign_in(9523) & VN_data_in(9523);
  VN1587_in2 <= VN_sign_in(9524) & VN_data_in(9524);
  VN1587_in3 <= VN_sign_in(9525) & VN_data_in(9525);
  VN1587_in4 <= VN_sign_in(9526) & VN_data_in(9526);
  VN1587_in5 <= VN_sign_in(9527) & VN_data_in(9527);
  VN1588_in0 <= VN_sign_in(9528) & VN_data_in(9528);
  VN1588_in1 <= VN_sign_in(9529) & VN_data_in(9529);
  VN1588_in2 <= VN_sign_in(9530) & VN_data_in(9530);
  VN1588_in3 <= VN_sign_in(9531) & VN_data_in(9531);
  VN1588_in4 <= VN_sign_in(9532) & VN_data_in(9532);
  VN1588_in5 <= VN_sign_in(9533) & VN_data_in(9533);
  VN1589_in0 <= VN_sign_in(9534) & VN_data_in(9534);
  VN1589_in1 <= VN_sign_in(9535) & VN_data_in(9535);
  VN1589_in2 <= VN_sign_in(9536) & VN_data_in(9536);
  VN1589_in3 <= VN_sign_in(9537) & VN_data_in(9537);
  VN1589_in4 <= VN_sign_in(9538) & VN_data_in(9538);
  VN1589_in5 <= VN_sign_in(9539) & VN_data_in(9539);
  VN1590_in0 <= VN_sign_in(9540) & VN_data_in(9540);
  VN1590_in1 <= VN_sign_in(9541) & VN_data_in(9541);
  VN1590_in2 <= VN_sign_in(9542) & VN_data_in(9542);
  VN1590_in3 <= VN_sign_in(9543) & VN_data_in(9543);
  VN1590_in4 <= VN_sign_in(9544) & VN_data_in(9544);
  VN1590_in5 <= VN_sign_in(9545) & VN_data_in(9545);
  VN1591_in0 <= VN_sign_in(9546) & VN_data_in(9546);
  VN1591_in1 <= VN_sign_in(9547) & VN_data_in(9547);
  VN1591_in2 <= VN_sign_in(9548) & VN_data_in(9548);
  VN1591_in3 <= VN_sign_in(9549) & VN_data_in(9549);
  VN1591_in4 <= VN_sign_in(9550) & VN_data_in(9550);
  VN1591_in5 <= VN_sign_in(9551) & VN_data_in(9551);
  VN1592_in0 <= VN_sign_in(9552) & VN_data_in(9552);
  VN1592_in1 <= VN_sign_in(9553) & VN_data_in(9553);
  VN1592_in2 <= VN_sign_in(9554) & VN_data_in(9554);
  VN1592_in3 <= VN_sign_in(9555) & VN_data_in(9555);
  VN1592_in4 <= VN_sign_in(9556) & VN_data_in(9556);
  VN1592_in5 <= VN_sign_in(9557) & VN_data_in(9557);
  VN1593_in0 <= VN_sign_in(9558) & VN_data_in(9558);
  VN1593_in1 <= VN_sign_in(9559) & VN_data_in(9559);
  VN1593_in2 <= VN_sign_in(9560) & VN_data_in(9560);
  VN1593_in3 <= VN_sign_in(9561) & VN_data_in(9561);
  VN1593_in4 <= VN_sign_in(9562) & VN_data_in(9562);
  VN1593_in5 <= VN_sign_in(9563) & VN_data_in(9563);
  VN1594_in0 <= VN_sign_in(9564) & VN_data_in(9564);
  VN1594_in1 <= VN_sign_in(9565) & VN_data_in(9565);
  VN1594_in2 <= VN_sign_in(9566) & VN_data_in(9566);
  VN1594_in3 <= VN_sign_in(9567) & VN_data_in(9567);
  VN1594_in4 <= VN_sign_in(9568) & VN_data_in(9568);
  VN1594_in5 <= VN_sign_in(9569) & VN_data_in(9569);
  VN1595_in0 <= VN_sign_in(9570) & VN_data_in(9570);
  VN1595_in1 <= VN_sign_in(9571) & VN_data_in(9571);
  VN1595_in2 <= VN_sign_in(9572) & VN_data_in(9572);
  VN1595_in3 <= VN_sign_in(9573) & VN_data_in(9573);
  VN1595_in4 <= VN_sign_in(9574) & VN_data_in(9574);
  VN1595_in5 <= VN_sign_in(9575) & VN_data_in(9575);
  VN1596_in0 <= VN_sign_in(9576) & VN_data_in(9576);
  VN1596_in1 <= VN_sign_in(9577) & VN_data_in(9577);
  VN1596_in2 <= VN_sign_in(9578) & VN_data_in(9578);
  VN1596_in3 <= VN_sign_in(9579) & VN_data_in(9579);
  VN1596_in4 <= VN_sign_in(9580) & VN_data_in(9580);
  VN1596_in5 <= VN_sign_in(9581) & VN_data_in(9581);
  VN1597_in0 <= VN_sign_in(9582) & VN_data_in(9582);
  VN1597_in1 <= VN_sign_in(9583) & VN_data_in(9583);
  VN1597_in2 <= VN_sign_in(9584) & VN_data_in(9584);
  VN1597_in3 <= VN_sign_in(9585) & VN_data_in(9585);
  VN1597_in4 <= VN_sign_in(9586) & VN_data_in(9586);
  VN1597_in5 <= VN_sign_in(9587) & VN_data_in(9587);
  VN1598_in0 <= VN_sign_in(9588) & VN_data_in(9588);
  VN1598_in1 <= VN_sign_in(9589) & VN_data_in(9589);
  VN1598_in2 <= VN_sign_in(9590) & VN_data_in(9590);
  VN1598_in3 <= VN_sign_in(9591) & VN_data_in(9591);
  VN1598_in4 <= VN_sign_in(9592) & VN_data_in(9592);
  VN1598_in5 <= VN_sign_in(9593) & VN_data_in(9593);
  VN1599_in0 <= VN_sign_in(9594) & VN_data_in(9594);
  VN1599_in1 <= VN_sign_in(9595) & VN_data_in(9595);
  VN1599_in2 <= VN_sign_in(9596) & VN_data_in(9596);
  VN1599_in3 <= VN_sign_in(9597) & VN_data_in(9597);
  VN1599_in4 <= VN_sign_in(9598) & VN_data_in(9598);
  VN1599_in5 <= VN_sign_in(9599) & VN_data_in(9599);
  VN1600_in0 <= VN_sign_in(9600) & VN_data_in(9600);
  VN1600_in1 <= VN_sign_in(9601) & VN_data_in(9601);
  VN1600_in2 <= VN_sign_in(9602) & VN_data_in(9602);
  VN1600_in3 <= VN_sign_in(9603) & VN_data_in(9603);
  VN1600_in4 <= VN_sign_in(9604) & VN_data_in(9604);
  VN1600_in5 <= VN_sign_in(9605) & VN_data_in(9605);
  VN1601_in0 <= VN_sign_in(9606) & VN_data_in(9606);
  VN1601_in1 <= VN_sign_in(9607) & VN_data_in(9607);
  VN1601_in2 <= VN_sign_in(9608) & VN_data_in(9608);
  VN1601_in3 <= VN_sign_in(9609) & VN_data_in(9609);
  VN1601_in4 <= VN_sign_in(9610) & VN_data_in(9610);
  VN1601_in5 <= VN_sign_in(9611) & VN_data_in(9611);
  VN1602_in0 <= VN_sign_in(9612) & VN_data_in(9612);
  VN1602_in1 <= VN_sign_in(9613) & VN_data_in(9613);
  VN1602_in2 <= VN_sign_in(9614) & VN_data_in(9614);
  VN1602_in3 <= VN_sign_in(9615) & VN_data_in(9615);
  VN1602_in4 <= VN_sign_in(9616) & VN_data_in(9616);
  VN1602_in5 <= VN_sign_in(9617) & VN_data_in(9617);
  VN1603_in0 <= VN_sign_in(9618) & VN_data_in(9618);
  VN1603_in1 <= VN_sign_in(9619) & VN_data_in(9619);
  VN1603_in2 <= VN_sign_in(9620) & VN_data_in(9620);
  VN1603_in3 <= VN_sign_in(9621) & VN_data_in(9621);
  VN1603_in4 <= VN_sign_in(9622) & VN_data_in(9622);
  VN1603_in5 <= VN_sign_in(9623) & VN_data_in(9623);
  VN1604_in0 <= VN_sign_in(9624) & VN_data_in(9624);
  VN1604_in1 <= VN_sign_in(9625) & VN_data_in(9625);
  VN1604_in2 <= VN_sign_in(9626) & VN_data_in(9626);
  VN1604_in3 <= VN_sign_in(9627) & VN_data_in(9627);
  VN1604_in4 <= VN_sign_in(9628) & VN_data_in(9628);
  VN1604_in5 <= VN_sign_in(9629) & VN_data_in(9629);
  VN1605_in0 <= VN_sign_in(9630) & VN_data_in(9630);
  VN1605_in1 <= VN_sign_in(9631) & VN_data_in(9631);
  VN1605_in2 <= VN_sign_in(9632) & VN_data_in(9632);
  VN1605_in3 <= VN_sign_in(9633) & VN_data_in(9633);
  VN1605_in4 <= VN_sign_in(9634) & VN_data_in(9634);
  VN1605_in5 <= VN_sign_in(9635) & VN_data_in(9635);
  VN1606_in0 <= VN_sign_in(9636) & VN_data_in(9636);
  VN1606_in1 <= VN_sign_in(9637) & VN_data_in(9637);
  VN1606_in2 <= VN_sign_in(9638) & VN_data_in(9638);
  VN1606_in3 <= VN_sign_in(9639) & VN_data_in(9639);
  VN1606_in4 <= VN_sign_in(9640) & VN_data_in(9640);
  VN1606_in5 <= VN_sign_in(9641) & VN_data_in(9641);
  VN1607_in0 <= VN_sign_in(9642) & VN_data_in(9642);
  VN1607_in1 <= VN_sign_in(9643) & VN_data_in(9643);
  VN1607_in2 <= VN_sign_in(9644) & VN_data_in(9644);
  VN1607_in3 <= VN_sign_in(9645) & VN_data_in(9645);
  VN1607_in4 <= VN_sign_in(9646) & VN_data_in(9646);
  VN1607_in5 <= VN_sign_in(9647) & VN_data_in(9647);
  VN1608_in0 <= VN_sign_in(9648) & VN_data_in(9648);
  VN1608_in1 <= VN_sign_in(9649) & VN_data_in(9649);
  VN1608_in2 <= VN_sign_in(9650) & VN_data_in(9650);
  VN1608_in3 <= VN_sign_in(9651) & VN_data_in(9651);
  VN1608_in4 <= VN_sign_in(9652) & VN_data_in(9652);
  VN1608_in5 <= VN_sign_in(9653) & VN_data_in(9653);
  VN1609_in0 <= VN_sign_in(9654) & VN_data_in(9654);
  VN1609_in1 <= VN_sign_in(9655) & VN_data_in(9655);
  VN1609_in2 <= VN_sign_in(9656) & VN_data_in(9656);
  VN1609_in3 <= VN_sign_in(9657) & VN_data_in(9657);
  VN1609_in4 <= VN_sign_in(9658) & VN_data_in(9658);
  VN1609_in5 <= VN_sign_in(9659) & VN_data_in(9659);
  VN1610_in0 <= VN_sign_in(9660) & VN_data_in(9660);
  VN1610_in1 <= VN_sign_in(9661) & VN_data_in(9661);
  VN1610_in2 <= VN_sign_in(9662) & VN_data_in(9662);
  VN1610_in3 <= VN_sign_in(9663) & VN_data_in(9663);
  VN1610_in4 <= VN_sign_in(9664) & VN_data_in(9664);
  VN1610_in5 <= VN_sign_in(9665) & VN_data_in(9665);
  VN1611_in0 <= VN_sign_in(9666) & VN_data_in(9666);
  VN1611_in1 <= VN_sign_in(9667) & VN_data_in(9667);
  VN1611_in2 <= VN_sign_in(9668) & VN_data_in(9668);
  VN1611_in3 <= VN_sign_in(9669) & VN_data_in(9669);
  VN1611_in4 <= VN_sign_in(9670) & VN_data_in(9670);
  VN1611_in5 <= VN_sign_in(9671) & VN_data_in(9671);
  VN1612_in0 <= VN_sign_in(9672) & VN_data_in(9672);
  VN1612_in1 <= VN_sign_in(9673) & VN_data_in(9673);
  VN1612_in2 <= VN_sign_in(9674) & VN_data_in(9674);
  VN1612_in3 <= VN_sign_in(9675) & VN_data_in(9675);
  VN1612_in4 <= VN_sign_in(9676) & VN_data_in(9676);
  VN1612_in5 <= VN_sign_in(9677) & VN_data_in(9677);
  VN1613_in0 <= VN_sign_in(9678) & VN_data_in(9678);
  VN1613_in1 <= VN_sign_in(9679) & VN_data_in(9679);
  VN1613_in2 <= VN_sign_in(9680) & VN_data_in(9680);
  VN1613_in3 <= VN_sign_in(9681) & VN_data_in(9681);
  VN1613_in4 <= VN_sign_in(9682) & VN_data_in(9682);
  VN1613_in5 <= VN_sign_in(9683) & VN_data_in(9683);
  VN1614_in0 <= VN_sign_in(9684) & VN_data_in(9684);
  VN1614_in1 <= VN_sign_in(9685) & VN_data_in(9685);
  VN1614_in2 <= VN_sign_in(9686) & VN_data_in(9686);
  VN1614_in3 <= VN_sign_in(9687) & VN_data_in(9687);
  VN1614_in4 <= VN_sign_in(9688) & VN_data_in(9688);
  VN1614_in5 <= VN_sign_in(9689) & VN_data_in(9689);
  VN1615_in0 <= VN_sign_in(9690) & VN_data_in(9690);
  VN1615_in1 <= VN_sign_in(9691) & VN_data_in(9691);
  VN1615_in2 <= VN_sign_in(9692) & VN_data_in(9692);
  VN1615_in3 <= VN_sign_in(9693) & VN_data_in(9693);
  VN1615_in4 <= VN_sign_in(9694) & VN_data_in(9694);
  VN1615_in5 <= VN_sign_in(9695) & VN_data_in(9695);
  VN1616_in0 <= VN_sign_in(9696) & VN_data_in(9696);
  VN1616_in1 <= VN_sign_in(9697) & VN_data_in(9697);
  VN1616_in2 <= VN_sign_in(9698) & VN_data_in(9698);
  VN1616_in3 <= VN_sign_in(9699) & VN_data_in(9699);
  VN1616_in4 <= VN_sign_in(9700) & VN_data_in(9700);
  VN1616_in5 <= VN_sign_in(9701) & VN_data_in(9701);
  VN1617_in0 <= VN_sign_in(9702) & VN_data_in(9702);
  VN1617_in1 <= VN_sign_in(9703) & VN_data_in(9703);
  VN1617_in2 <= VN_sign_in(9704) & VN_data_in(9704);
  VN1617_in3 <= VN_sign_in(9705) & VN_data_in(9705);
  VN1617_in4 <= VN_sign_in(9706) & VN_data_in(9706);
  VN1617_in5 <= VN_sign_in(9707) & VN_data_in(9707);
  VN1618_in0 <= VN_sign_in(9708) & VN_data_in(9708);
  VN1618_in1 <= VN_sign_in(9709) & VN_data_in(9709);
  VN1618_in2 <= VN_sign_in(9710) & VN_data_in(9710);
  VN1618_in3 <= VN_sign_in(9711) & VN_data_in(9711);
  VN1618_in4 <= VN_sign_in(9712) & VN_data_in(9712);
  VN1618_in5 <= VN_sign_in(9713) & VN_data_in(9713);
  VN1619_in0 <= VN_sign_in(9714) & VN_data_in(9714);
  VN1619_in1 <= VN_sign_in(9715) & VN_data_in(9715);
  VN1619_in2 <= VN_sign_in(9716) & VN_data_in(9716);
  VN1619_in3 <= VN_sign_in(9717) & VN_data_in(9717);
  VN1619_in4 <= VN_sign_in(9718) & VN_data_in(9718);
  VN1619_in5 <= VN_sign_in(9719) & VN_data_in(9719);
  VN1620_in0 <= VN_sign_in(9720) & VN_data_in(9720);
  VN1620_in1 <= VN_sign_in(9721) & VN_data_in(9721);
  VN1620_in2 <= VN_sign_in(9722) & VN_data_in(9722);
  VN1620_in3 <= VN_sign_in(9723) & VN_data_in(9723);
  VN1620_in4 <= VN_sign_in(9724) & VN_data_in(9724);
  VN1620_in5 <= VN_sign_in(9725) & VN_data_in(9725);
  VN1621_in0 <= VN_sign_in(9726) & VN_data_in(9726);
  VN1621_in1 <= VN_sign_in(9727) & VN_data_in(9727);
  VN1621_in2 <= VN_sign_in(9728) & VN_data_in(9728);
  VN1621_in3 <= VN_sign_in(9729) & VN_data_in(9729);
  VN1621_in4 <= VN_sign_in(9730) & VN_data_in(9730);
  VN1621_in5 <= VN_sign_in(9731) & VN_data_in(9731);
  VN1622_in0 <= VN_sign_in(9732) & VN_data_in(9732);
  VN1622_in1 <= VN_sign_in(9733) & VN_data_in(9733);
  VN1622_in2 <= VN_sign_in(9734) & VN_data_in(9734);
  VN1622_in3 <= VN_sign_in(9735) & VN_data_in(9735);
  VN1622_in4 <= VN_sign_in(9736) & VN_data_in(9736);
  VN1622_in5 <= VN_sign_in(9737) & VN_data_in(9737);
  VN1623_in0 <= VN_sign_in(9738) & VN_data_in(9738);
  VN1623_in1 <= VN_sign_in(9739) & VN_data_in(9739);
  VN1623_in2 <= VN_sign_in(9740) & VN_data_in(9740);
  VN1623_in3 <= VN_sign_in(9741) & VN_data_in(9741);
  VN1623_in4 <= VN_sign_in(9742) & VN_data_in(9742);
  VN1623_in5 <= VN_sign_in(9743) & VN_data_in(9743);
  VN1624_in0 <= VN_sign_in(9744) & VN_data_in(9744);
  VN1624_in1 <= VN_sign_in(9745) & VN_data_in(9745);
  VN1624_in2 <= VN_sign_in(9746) & VN_data_in(9746);
  VN1624_in3 <= VN_sign_in(9747) & VN_data_in(9747);
  VN1624_in4 <= VN_sign_in(9748) & VN_data_in(9748);
  VN1624_in5 <= VN_sign_in(9749) & VN_data_in(9749);
  VN1625_in0 <= VN_sign_in(9750) & VN_data_in(9750);
  VN1625_in1 <= VN_sign_in(9751) & VN_data_in(9751);
  VN1625_in2 <= VN_sign_in(9752) & VN_data_in(9752);
  VN1625_in3 <= VN_sign_in(9753) & VN_data_in(9753);
  VN1625_in4 <= VN_sign_in(9754) & VN_data_in(9754);
  VN1625_in5 <= VN_sign_in(9755) & VN_data_in(9755);
  VN1626_in0 <= VN_sign_in(9756) & VN_data_in(9756);
  VN1626_in1 <= VN_sign_in(9757) & VN_data_in(9757);
  VN1626_in2 <= VN_sign_in(9758) & VN_data_in(9758);
  VN1626_in3 <= VN_sign_in(9759) & VN_data_in(9759);
  VN1626_in4 <= VN_sign_in(9760) & VN_data_in(9760);
  VN1626_in5 <= VN_sign_in(9761) & VN_data_in(9761);
  VN1627_in0 <= VN_sign_in(9762) & VN_data_in(9762);
  VN1627_in1 <= VN_sign_in(9763) & VN_data_in(9763);
  VN1627_in2 <= VN_sign_in(9764) & VN_data_in(9764);
  VN1627_in3 <= VN_sign_in(9765) & VN_data_in(9765);
  VN1627_in4 <= VN_sign_in(9766) & VN_data_in(9766);
  VN1627_in5 <= VN_sign_in(9767) & VN_data_in(9767);
  VN1628_in0 <= VN_sign_in(9768) & VN_data_in(9768);
  VN1628_in1 <= VN_sign_in(9769) & VN_data_in(9769);
  VN1628_in2 <= VN_sign_in(9770) & VN_data_in(9770);
  VN1628_in3 <= VN_sign_in(9771) & VN_data_in(9771);
  VN1628_in4 <= VN_sign_in(9772) & VN_data_in(9772);
  VN1628_in5 <= VN_sign_in(9773) & VN_data_in(9773);
  VN1629_in0 <= VN_sign_in(9774) & VN_data_in(9774);
  VN1629_in1 <= VN_sign_in(9775) & VN_data_in(9775);
  VN1629_in2 <= VN_sign_in(9776) & VN_data_in(9776);
  VN1629_in3 <= VN_sign_in(9777) & VN_data_in(9777);
  VN1629_in4 <= VN_sign_in(9778) & VN_data_in(9778);
  VN1629_in5 <= VN_sign_in(9779) & VN_data_in(9779);
  VN1630_in0 <= VN_sign_in(9780) & VN_data_in(9780);
  VN1630_in1 <= VN_sign_in(9781) & VN_data_in(9781);
  VN1630_in2 <= VN_sign_in(9782) & VN_data_in(9782);
  VN1630_in3 <= VN_sign_in(9783) & VN_data_in(9783);
  VN1630_in4 <= VN_sign_in(9784) & VN_data_in(9784);
  VN1630_in5 <= VN_sign_in(9785) & VN_data_in(9785);
  VN1631_in0 <= VN_sign_in(9786) & VN_data_in(9786);
  VN1631_in1 <= VN_sign_in(9787) & VN_data_in(9787);
  VN1631_in2 <= VN_sign_in(9788) & VN_data_in(9788);
  VN1631_in3 <= VN_sign_in(9789) & VN_data_in(9789);
  VN1631_in4 <= VN_sign_in(9790) & VN_data_in(9790);
  VN1631_in5 <= VN_sign_in(9791) & VN_data_in(9791);
  VN1632_in0 <= VN_sign_in(9792) & VN_data_in(9792);
  VN1632_in1 <= VN_sign_in(9793) & VN_data_in(9793);
  VN1632_in2 <= VN_sign_in(9794) & VN_data_in(9794);
  VN1632_in3 <= VN_sign_in(9795) & VN_data_in(9795);
  VN1632_in4 <= VN_sign_in(9796) & VN_data_in(9796);
  VN1632_in5 <= VN_sign_in(9797) & VN_data_in(9797);
  VN1633_in0 <= VN_sign_in(9798) & VN_data_in(9798);
  VN1633_in1 <= VN_sign_in(9799) & VN_data_in(9799);
  VN1633_in2 <= VN_sign_in(9800) & VN_data_in(9800);
  VN1633_in3 <= VN_sign_in(9801) & VN_data_in(9801);
  VN1633_in4 <= VN_sign_in(9802) & VN_data_in(9802);
  VN1633_in5 <= VN_sign_in(9803) & VN_data_in(9803);
  VN1634_in0 <= VN_sign_in(9804) & VN_data_in(9804);
  VN1634_in1 <= VN_sign_in(9805) & VN_data_in(9805);
  VN1634_in2 <= VN_sign_in(9806) & VN_data_in(9806);
  VN1634_in3 <= VN_sign_in(9807) & VN_data_in(9807);
  VN1634_in4 <= VN_sign_in(9808) & VN_data_in(9808);
  VN1634_in5 <= VN_sign_in(9809) & VN_data_in(9809);
  VN1635_in0 <= VN_sign_in(9810) & VN_data_in(9810);
  VN1635_in1 <= VN_sign_in(9811) & VN_data_in(9811);
  VN1635_in2 <= VN_sign_in(9812) & VN_data_in(9812);
  VN1635_in3 <= VN_sign_in(9813) & VN_data_in(9813);
  VN1635_in4 <= VN_sign_in(9814) & VN_data_in(9814);
  VN1635_in5 <= VN_sign_in(9815) & VN_data_in(9815);
  VN1636_in0 <= VN_sign_in(9816) & VN_data_in(9816);
  VN1636_in1 <= VN_sign_in(9817) & VN_data_in(9817);
  VN1636_in2 <= VN_sign_in(9818) & VN_data_in(9818);
  VN1636_in3 <= VN_sign_in(9819) & VN_data_in(9819);
  VN1636_in4 <= VN_sign_in(9820) & VN_data_in(9820);
  VN1636_in5 <= VN_sign_in(9821) & VN_data_in(9821);
  VN1637_in0 <= VN_sign_in(9822) & VN_data_in(9822);
  VN1637_in1 <= VN_sign_in(9823) & VN_data_in(9823);
  VN1637_in2 <= VN_sign_in(9824) & VN_data_in(9824);
  VN1637_in3 <= VN_sign_in(9825) & VN_data_in(9825);
  VN1637_in4 <= VN_sign_in(9826) & VN_data_in(9826);
  VN1637_in5 <= VN_sign_in(9827) & VN_data_in(9827);
  VN1638_in0 <= VN_sign_in(9828) & VN_data_in(9828);
  VN1638_in1 <= VN_sign_in(9829) & VN_data_in(9829);
  VN1638_in2 <= VN_sign_in(9830) & VN_data_in(9830);
  VN1638_in3 <= VN_sign_in(9831) & VN_data_in(9831);
  VN1638_in4 <= VN_sign_in(9832) & VN_data_in(9832);
  VN1638_in5 <= VN_sign_in(9833) & VN_data_in(9833);
  VN1639_in0 <= VN_sign_in(9834) & VN_data_in(9834);
  VN1639_in1 <= VN_sign_in(9835) & VN_data_in(9835);
  VN1639_in2 <= VN_sign_in(9836) & VN_data_in(9836);
  VN1639_in3 <= VN_sign_in(9837) & VN_data_in(9837);
  VN1639_in4 <= VN_sign_in(9838) & VN_data_in(9838);
  VN1639_in5 <= VN_sign_in(9839) & VN_data_in(9839);
  VN1640_in0 <= VN_sign_in(9840) & VN_data_in(9840);
  VN1640_in1 <= VN_sign_in(9841) & VN_data_in(9841);
  VN1640_in2 <= VN_sign_in(9842) & VN_data_in(9842);
  VN1640_in3 <= VN_sign_in(9843) & VN_data_in(9843);
  VN1640_in4 <= VN_sign_in(9844) & VN_data_in(9844);
  VN1640_in5 <= VN_sign_in(9845) & VN_data_in(9845);
  VN1641_in0 <= VN_sign_in(9846) & VN_data_in(9846);
  VN1641_in1 <= VN_sign_in(9847) & VN_data_in(9847);
  VN1641_in2 <= VN_sign_in(9848) & VN_data_in(9848);
  VN1641_in3 <= VN_sign_in(9849) & VN_data_in(9849);
  VN1641_in4 <= VN_sign_in(9850) & VN_data_in(9850);
  VN1641_in5 <= VN_sign_in(9851) & VN_data_in(9851);
  VN1642_in0 <= VN_sign_in(9852) & VN_data_in(9852);
  VN1642_in1 <= VN_sign_in(9853) & VN_data_in(9853);
  VN1642_in2 <= VN_sign_in(9854) & VN_data_in(9854);
  VN1642_in3 <= VN_sign_in(9855) & VN_data_in(9855);
  VN1642_in4 <= VN_sign_in(9856) & VN_data_in(9856);
  VN1642_in5 <= VN_sign_in(9857) & VN_data_in(9857);
  VN1643_in0 <= VN_sign_in(9858) & VN_data_in(9858);
  VN1643_in1 <= VN_sign_in(9859) & VN_data_in(9859);
  VN1643_in2 <= VN_sign_in(9860) & VN_data_in(9860);
  VN1643_in3 <= VN_sign_in(9861) & VN_data_in(9861);
  VN1643_in4 <= VN_sign_in(9862) & VN_data_in(9862);
  VN1643_in5 <= VN_sign_in(9863) & VN_data_in(9863);
  VN1644_in0 <= VN_sign_in(9864) & VN_data_in(9864);
  VN1644_in1 <= VN_sign_in(9865) & VN_data_in(9865);
  VN1644_in2 <= VN_sign_in(9866) & VN_data_in(9866);
  VN1644_in3 <= VN_sign_in(9867) & VN_data_in(9867);
  VN1644_in4 <= VN_sign_in(9868) & VN_data_in(9868);
  VN1644_in5 <= VN_sign_in(9869) & VN_data_in(9869);
  VN1645_in0 <= VN_sign_in(9870) & VN_data_in(9870);
  VN1645_in1 <= VN_sign_in(9871) & VN_data_in(9871);
  VN1645_in2 <= VN_sign_in(9872) & VN_data_in(9872);
  VN1645_in3 <= VN_sign_in(9873) & VN_data_in(9873);
  VN1645_in4 <= VN_sign_in(9874) & VN_data_in(9874);
  VN1645_in5 <= VN_sign_in(9875) & VN_data_in(9875);
  VN1646_in0 <= VN_sign_in(9876) & VN_data_in(9876);
  VN1646_in1 <= VN_sign_in(9877) & VN_data_in(9877);
  VN1646_in2 <= VN_sign_in(9878) & VN_data_in(9878);
  VN1646_in3 <= VN_sign_in(9879) & VN_data_in(9879);
  VN1646_in4 <= VN_sign_in(9880) & VN_data_in(9880);
  VN1646_in5 <= VN_sign_in(9881) & VN_data_in(9881);
  VN1647_in0 <= VN_sign_in(9882) & VN_data_in(9882);
  VN1647_in1 <= VN_sign_in(9883) & VN_data_in(9883);
  VN1647_in2 <= VN_sign_in(9884) & VN_data_in(9884);
  VN1647_in3 <= VN_sign_in(9885) & VN_data_in(9885);
  VN1647_in4 <= VN_sign_in(9886) & VN_data_in(9886);
  VN1647_in5 <= VN_sign_in(9887) & VN_data_in(9887);
  VN1648_in0 <= VN_sign_in(9888) & VN_data_in(9888);
  VN1648_in1 <= VN_sign_in(9889) & VN_data_in(9889);
  VN1648_in2 <= VN_sign_in(9890) & VN_data_in(9890);
  VN1648_in3 <= VN_sign_in(9891) & VN_data_in(9891);
  VN1648_in4 <= VN_sign_in(9892) & VN_data_in(9892);
  VN1648_in5 <= VN_sign_in(9893) & VN_data_in(9893);
  VN1649_in0 <= VN_sign_in(9894) & VN_data_in(9894);
  VN1649_in1 <= VN_sign_in(9895) & VN_data_in(9895);
  VN1649_in2 <= VN_sign_in(9896) & VN_data_in(9896);
  VN1649_in3 <= VN_sign_in(9897) & VN_data_in(9897);
  VN1649_in4 <= VN_sign_in(9898) & VN_data_in(9898);
  VN1649_in5 <= VN_sign_in(9899) & VN_data_in(9899);
  VN1650_in0 <= VN_sign_in(9900) & VN_data_in(9900);
  VN1650_in1 <= VN_sign_in(9901) & VN_data_in(9901);
  VN1650_in2 <= VN_sign_in(9902) & VN_data_in(9902);
  VN1650_in3 <= VN_sign_in(9903) & VN_data_in(9903);
  VN1650_in4 <= VN_sign_in(9904) & VN_data_in(9904);
  VN1650_in5 <= VN_sign_in(9905) & VN_data_in(9905);
  VN1651_in0 <= VN_sign_in(9906) & VN_data_in(9906);
  VN1651_in1 <= VN_sign_in(9907) & VN_data_in(9907);
  VN1651_in2 <= VN_sign_in(9908) & VN_data_in(9908);
  VN1651_in3 <= VN_sign_in(9909) & VN_data_in(9909);
  VN1651_in4 <= VN_sign_in(9910) & VN_data_in(9910);
  VN1651_in5 <= VN_sign_in(9911) & VN_data_in(9911);
  VN1652_in0 <= VN_sign_in(9912) & VN_data_in(9912);
  VN1652_in1 <= VN_sign_in(9913) & VN_data_in(9913);
  VN1652_in2 <= VN_sign_in(9914) & VN_data_in(9914);
  VN1652_in3 <= VN_sign_in(9915) & VN_data_in(9915);
  VN1652_in4 <= VN_sign_in(9916) & VN_data_in(9916);
  VN1652_in5 <= VN_sign_in(9917) & VN_data_in(9917);
  VN1653_in0 <= VN_sign_in(9918) & VN_data_in(9918);
  VN1653_in1 <= VN_sign_in(9919) & VN_data_in(9919);
  VN1653_in2 <= VN_sign_in(9920) & VN_data_in(9920);
  VN1653_in3 <= VN_sign_in(9921) & VN_data_in(9921);
  VN1653_in4 <= VN_sign_in(9922) & VN_data_in(9922);
  VN1653_in5 <= VN_sign_in(9923) & VN_data_in(9923);
  VN1654_in0 <= VN_sign_in(9924) & VN_data_in(9924);
  VN1654_in1 <= VN_sign_in(9925) & VN_data_in(9925);
  VN1654_in2 <= VN_sign_in(9926) & VN_data_in(9926);
  VN1654_in3 <= VN_sign_in(9927) & VN_data_in(9927);
  VN1654_in4 <= VN_sign_in(9928) & VN_data_in(9928);
  VN1654_in5 <= VN_sign_in(9929) & VN_data_in(9929);
  VN1655_in0 <= VN_sign_in(9930) & VN_data_in(9930);
  VN1655_in1 <= VN_sign_in(9931) & VN_data_in(9931);
  VN1655_in2 <= VN_sign_in(9932) & VN_data_in(9932);
  VN1655_in3 <= VN_sign_in(9933) & VN_data_in(9933);
  VN1655_in4 <= VN_sign_in(9934) & VN_data_in(9934);
  VN1655_in5 <= VN_sign_in(9935) & VN_data_in(9935);
  VN1656_in0 <= VN_sign_in(9936) & VN_data_in(9936);
  VN1656_in1 <= VN_sign_in(9937) & VN_data_in(9937);
  VN1656_in2 <= VN_sign_in(9938) & VN_data_in(9938);
  VN1656_in3 <= VN_sign_in(9939) & VN_data_in(9939);
  VN1656_in4 <= VN_sign_in(9940) & VN_data_in(9940);
  VN1656_in5 <= VN_sign_in(9941) & VN_data_in(9941);
  VN1657_in0 <= VN_sign_in(9942) & VN_data_in(9942);
  VN1657_in1 <= VN_sign_in(9943) & VN_data_in(9943);
  VN1657_in2 <= VN_sign_in(9944) & VN_data_in(9944);
  VN1657_in3 <= VN_sign_in(9945) & VN_data_in(9945);
  VN1657_in4 <= VN_sign_in(9946) & VN_data_in(9946);
  VN1657_in5 <= VN_sign_in(9947) & VN_data_in(9947);
  VN1658_in0 <= VN_sign_in(9948) & VN_data_in(9948);
  VN1658_in1 <= VN_sign_in(9949) & VN_data_in(9949);
  VN1658_in2 <= VN_sign_in(9950) & VN_data_in(9950);
  VN1658_in3 <= VN_sign_in(9951) & VN_data_in(9951);
  VN1658_in4 <= VN_sign_in(9952) & VN_data_in(9952);
  VN1658_in5 <= VN_sign_in(9953) & VN_data_in(9953);
  VN1659_in0 <= VN_sign_in(9954) & VN_data_in(9954);
  VN1659_in1 <= VN_sign_in(9955) & VN_data_in(9955);
  VN1659_in2 <= VN_sign_in(9956) & VN_data_in(9956);
  VN1659_in3 <= VN_sign_in(9957) & VN_data_in(9957);
  VN1659_in4 <= VN_sign_in(9958) & VN_data_in(9958);
  VN1659_in5 <= VN_sign_in(9959) & VN_data_in(9959);
  VN1660_in0 <= VN_sign_in(9960) & VN_data_in(9960);
  VN1660_in1 <= VN_sign_in(9961) & VN_data_in(9961);
  VN1660_in2 <= VN_sign_in(9962) & VN_data_in(9962);
  VN1660_in3 <= VN_sign_in(9963) & VN_data_in(9963);
  VN1660_in4 <= VN_sign_in(9964) & VN_data_in(9964);
  VN1660_in5 <= VN_sign_in(9965) & VN_data_in(9965);
  VN1661_in0 <= VN_sign_in(9966) & VN_data_in(9966);
  VN1661_in1 <= VN_sign_in(9967) & VN_data_in(9967);
  VN1661_in2 <= VN_sign_in(9968) & VN_data_in(9968);
  VN1661_in3 <= VN_sign_in(9969) & VN_data_in(9969);
  VN1661_in4 <= VN_sign_in(9970) & VN_data_in(9970);
  VN1661_in5 <= VN_sign_in(9971) & VN_data_in(9971);
  VN1662_in0 <= VN_sign_in(9972) & VN_data_in(9972);
  VN1662_in1 <= VN_sign_in(9973) & VN_data_in(9973);
  VN1662_in2 <= VN_sign_in(9974) & VN_data_in(9974);
  VN1662_in3 <= VN_sign_in(9975) & VN_data_in(9975);
  VN1662_in4 <= VN_sign_in(9976) & VN_data_in(9976);
  VN1662_in5 <= VN_sign_in(9977) & VN_data_in(9977);
  VN1663_in0 <= VN_sign_in(9978) & VN_data_in(9978);
  VN1663_in1 <= VN_sign_in(9979) & VN_data_in(9979);
  VN1663_in2 <= VN_sign_in(9980) & VN_data_in(9980);
  VN1663_in3 <= VN_sign_in(9981) & VN_data_in(9981);
  VN1663_in4 <= VN_sign_in(9982) & VN_data_in(9982);
  VN1663_in5 <= VN_sign_in(9983) & VN_data_in(9983);
  VN1664_in0 <= VN_sign_in(9984) & VN_data_in(9984);
  VN1664_in1 <= VN_sign_in(9985) & VN_data_in(9985);
  VN1664_in2 <= VN_sign_in(9986) & VN_data_in(9986);
  VN1664_in3 <= VN_sign_in(9987) & VN_data_in(9987);
  VN1664_in4 <= VN_sign_in(9988) & VN_data_in(9988);
  VN1664_in5 <= VN_sign_in(9989) & VN_data_in(9989);
  VN1665_in0 <= VN_sign_in(9990) & VN_data_in(9990);
  VN1665_in1 <= VN_sign_in(9991) & VN_data_in(9991);
  VN1665_in2 <= VN_sign_in(9992) & VN_data_in(9992);
  VN1665_in3 <= VN_sign_in(9993) & VN_data_in(9993);
  VN1665_in4 <= VN_sign_in(9994) & VN_data_in(9994);
  VN1665_in5 <= VN_sign_in(9995) & VN_data_in(9995);
  VN1666_in0 <= VN_sign_in(9996) & VN_data_in(9996);
  VN1666_in1 <= VN_sign_in(9997) & VN_data_in(9997);
  VN1666_in2 <= VN_sign_in(9998) & VN_data_in(9998);
  VN1666_in3 <= VN_sign_in(9999) & VN_data_in(9999);
  VN1666_in4 <= VN_sign_in(10000) & VN_data_in(10000);
  VN1666_in5 <= VN_sign_in(10001) & VN_data_in(10001);
  VN1667_in0 <= VN_sign_in(10002) & VN_data_in(10002);
  VN1667_in1 <= VN_sign_in(10003) & VN_data_in(10003);
  VN1667_in2 <= VN_sign_in(10004) & VN_data_in(10004);
  VN1667_in3 <= VN_sign_in(10005) & VN_data_in(10005);
  VN1667_in4 <= VN_sign_in(10006) & VN_data_in(10006);
  VN1667_in5 <= VN_sign_in(10007) & VN_data_in(10007);
  VN1668_in0 <= VN_sign_in(10008) & VN_data_in(10008);
  VN1668_in1 <= VN_sign_in(10009) & VN_data_in(10009);
  VN1668_in2 <= VN_sign_in(10010) & VN_data_in(10010);
  VN1668_in3 <= VN_sign_in(10011) & VN_data_in(10011);
  VN1668_in4 <= VN_sign_in(10012) & VN_data_in(10012);
  VN1668_in5 <= VN_sign_in(10013) & VN_data_in(10013);
  VN1669_in0 <= VN_sign_in(10014) & VN_data_in(10014);
  VN1669_in1 <= VN_sign_in(10015) & VN_data_in(10015);
  VN1669_in2 <= VN_sign_in(10016) & VN_data_in(10016);
  VN1669_in3 <= VN_sign_in(10017) & VN_data_in(10017);
  VN1669_in4 <= VN_sign_in(10018) & VN_data_in(10018);
  VN1669_in5 <= VN_sign_in(10019) & VN_data_in(10019);
  VN1670_in0 <= VN_sign_in(10020) & VN_data_in(10020);
  VN1670_in1 <= VN_sign_in(10021) & VN_data_in(10021);
  VN1670_in2 <= VN_sign_in(10022) & VN_data_in(10022);
  VN1670_in3 <= VN_sign_in(10023) & VN_data_in(10023);
  VN1670_in4 <= VN_sign_in(10024) & VN_data_in(10024);
  VN1670_in5 <= VN_sign_in(10025) & VN_data_in(10025);
  VN1671_in0 <= VN_sign_in(10026) & VN_data_in(10026);
  VN1671_in1 <= VN_sign_in(10027) & VN_data_in(10027);
  VN1671_in2 <= VN_sign_in(10028) & VN_data_in(10028);
  VN1671_in3 <= VN_sign_in(10029) & VN_data_in(10029);
  VN1671_in4 <= VN_sign_in(10030) & VN_data_in(10030);
  VN1671_in5 <= VN_sign_in(10031) & VN_data_in(10031);
  VN1672_in0 <= VN_sign_in(10032) & VN_data_in(10032);
  VN1672_in1 <= VN_sign_in(10033) & VN_data_in(10033);
  VN1672_in2 <= VN_sign_in(10034) & VN_data_in(10034);
  VN1672_in3 <= VN_sign_in(10035) & VN_data_in(10035);
  VN1672_in4 <= VN_sign_in(10036) & VN_data_in(10036);
  VN1672_in5 <= VN_sign_in(10037) & VN_data_in(10037);
  VN1673_in0 <= VN_sign_in(10038) & VN_data_in(10038);
  VN1673_in1 <= VN_sign_in(10039) & VN_data_in(10039);
  VN1673_in2 <= VN_sign_in(10040) & VN_data_in(10040);
  VN1673_in3 <= VN_sign_in(10041) & VN_data_in(10041);
  VN1673_in4 <= VN_sign_in(10042) & VN_data_in(10042);
  VN1673_in5 <= VN_sign_in(10043) & VN_data_in(10043);
  VN1674_in0 <= VN_sign_in(10044) & VN_data_in(10044);
  VN1674_in1 <= VN_sign_in(10045) & VN_data_in(10045);
  VN1674_in2 <= VN_sign_in(10046) & VN_data_in(10046);
  VN1674_in3 <= VN_sign_in(10047) & VN_data_in(10047);
  VN1674_in4 <= VN_sign_in(10048) & VN_data_in(10048);
  VN1674_in5 <= VN_sign_in(10049) & VN_data_in(10049);
  VN1675_in0 <= VN_sign_in(10050) & VN_data_in(10050);
  VN1675_in1 <= VN_sign_in(10051) & VN_data_in(10051);
  VN1675_in2 <= VN_sign_in(10052) & VN_data_in(10052);
  VN1675_in3 <= VN_sign_in(10053) & VN_data_in(10053);
  VN1675_in4 <= VN_sign_in(10054) & VN_data_in(10054);
  VN1675_in5 <= VN_sign_in(10055) & VN_data_in(10055);
  VN1676_in0 <= VN_sign_in(10056) & VN_data_in(10056);
  VN1676_in1 <= VN_sign_in(10057) & VN_data_in(10057);
  VN1676_in2 <= VN_sign_in(10058) & VN_data_in(10058);
  VN1676_in3 <= VN_sign_in(10059) & VN_data_in(10059);
  VN1676_in4 <= VN_sign_in(10060) & VN_data_in(10060);
  VN1676_in5 <= VN_sign_in(10061) & VN_data_in(10061);
  VN1677_in0 <= VN_sign_in(10062) & VN_data_in(10062);
  VN1677_in1 <= VN_sign_in(10063) & VN_data_in(10063);
  VN1677_in2 <= VN_sign_in(10064) & VN_data_in(10064);
  VN1677_in3 <= VN_sign_in(10065) & VN_data_in(10065);
  VN1677_in4 <= VN_sign_in(10066) & VN_data_in(10066);
  VN1677_in5 <= VN_sign_in(10067) & VN_data_in(10067);
  VN1678_in0 <= VN_sign_in(10068) & VN_data_in(10068);
  VN1678_in1 <= VN_sign_in(10069) & VN_data_in(10069);
  VN1678_in2 <= VN_sign_in(10070) & VN_data_in(10070);
  VN1678_in3 <= VN_sign_in(10071) & VN_data_in(10071);
  VN1678_in4 <= VN_sign_in(10072) & VN_data_in(10072);
  VN1678_in5 <= VN_sign_in(10073) & VN_data_in(10073);
  VN1679_in0 <= VN_sign_in(10074) & VN_data_in(10074);
  VN1679_in1 <= VN_sign_in(10075) & VN_data_in(10075);
  VN1679_in2 <= VN_sign_in(10076) & VN_data_in(10076);
  VN1679_in3 <= VN_sign_in(10077) & VN_data_in(10077);
  VN1679_in4 <= VN_sign_in(10078) & VN_data_in(10078);
  VN1679_in5 <= VN_sign_in(10079) & VN_data_in(10079);
  VN1680_in0 <= VN_sign_in(10080) & VN_data_in(10080);
  VN1680_in1 <= VN_sign_in(10081) & VN_data_in(10081);
  VN1680_in2 <= VN_sign_in(10082) & VN_data_in(10082);
  VN1680_in3 <= VN_sign_in(10083) & VN_data_in(10083);
  VN1680_in4 <= VN_sign_in(10084) & VN_data_in(10084);
  VN1680_in5 <= VN_sign_in(10085) & VN_data_in(10085);
  VN1681_in0 <= VN_sign_in(10086) & VN_data_in(10086);
  VN1681_in1 <= VN_sign_in(10087) & VN_data_in(10087);
  VN1681_in2 <= VN_sign_in(10088) & VN_data_in(10088);
  VN1681_in3 <= VN_sign_in(10089) & VN_data_in(10089);
  VN1681_in4 <= VN_sign_in(10090) & VN_data_in(10090);
  VN1681_in5 <= VN_sign_in(10091) & VN_data_in(10091);
  VN1682_in0 <= VN_sign_in(10092) & VN_data_in(10092);
  VN1682_in1 <= VN_sign_in(10093) & VN_data_in(10093);
  VN1682_in2 <= VN_sign_in(10094) & VN_data_in(10094);
  VN1682_in3 <= VN_sign_in(10095) & VN_data_in(10095);
  VN1682_in4 <= VN_sign_in(10096) & VN_data_in(10096);
  VN1682_in5 <= VN_sign_in(10097) & VN_data_in(10097);
  VN1683_in0 <= VN_sign_in(10098) & VN_data_in(10098);
  VN1683_in1 <= VN_sign_in(10099) & VN_data_in(10099);
  VN1683_in2 <= VN_sign_in(10100) & VN_data_in(10100);
  VN1683_in3 <= VN_sign_in(10101) & VN_data_in(10101);
  VN1683_in4 <= VN_sign_in(10102) & VN_data_in(10102);
  VN1683_in5 <= VN_sign_in(10103) & VN_data_in(10103);
  VN1684_in0 <= VN_sign_in(10104) & VN_data_in(10104);
  VN1684_in1 <= VN_sign_in(10105) & VN_data_in(10105);
  VN1684_in2 <= VN_sign_in(10106) & VN_data_in(10106);
  VN1684_in3 <= VN_sign_in(10107) & VN_data_in(10107);
  VN1684_in4 <= VN_sign_in(10108) & VN_data_in(10108);
  VN1684_in5 <= VN_sign_in(10109) & VN_data_in(10109);
  VN1685_in0 <= VN_sign_in(10110) & VN_data_in(10110);
  VN1685_in1 <= VN_sign_in(10111) & VN_data_in(10111);
  VN1685_in2 <= VN_sign_in(10112) & VN_data_in(10112);
  VN1685_in3 <= VN_sign_in(10113) & VN_data_in(10113);
  VN1685_in4 <= VN_sign_in(10114) & VN_data_in(10114);
  VN1685_in5 <= VN_sign_in(10115) & VN_data_in(10115);
  VN1686_in0 <= VN_sign_in(10116) & VN_data_in(10116);
  VN1686_in1 <= VN_sign_in(10117) & VN_data_in(10117);
  VN1686_in2 <= VN_sign_in(10118) & VN_data_in(10118);
  VN1686_in3 <= VN_sign_in(10119) & VN_data_in(10119);
  VN1686_in4 <= VN_sign_in(10120) & VN_data_in(10120);
  VN1686_in5 <= VN_sign_in(10121) & VN_data_in(10121);
  VN1687_in0 <= VN_sign_in(10122) & VN_data_in(10122);
  VN1687_in1 <= VN_sign_in(10123) & VN_data_in(10123);
  VN1687_in2 <= VN_sign_in(10124) & VN_data_in(10124);
  VN1687_in3 <= VN_sign_in(10125) & VN_data_in(10125);
  VN1687_in4 <= VN_sign_in(10126) & VN_data_in(10126);
  VN1687_in5 <= VN_sign_in(10127) & VN_data_in(10127);
  VN1688_in0 <= VN_sign_in(10128) & VN_data_in(10128);
  VN1688_in1 <= VN_sign_in(10129) & VN_data_in(10129);
  VN1688_in2 <= VN_sign_in(10130) & VN_data_in(10130);
  VN1688_in3 <= VN_sign_in(10131) & VN_data_in(10131);
  VN1688_in4 <= VN_sign_in(10132) & VN_data_in(10132);
  VN1688_in5 <= VN_sign_in(10133) & VN_data_in(10133);
  VN1689_in0 <= VN_sign_in(10134) & VN_data_in(10134);
  VN1689_in1 <= VN_sign_in(10135) & VN_data_in(10135);
  VN1689_in2 <= VN_sign_in(10136) & VN_data_in(10136);
  VN1689_in3 <= VN_sign_in(10137) & VN_data_in(10137);
  VN1689_in4 <= VN_sign_in(10138) & VN_data_in(10138);
  VN1689_in5 <= VN_sign_in(10139) & VN_data_in(10139);
  VN1690_in0 <= VN_sign_in(10140) & VN_data_in(10140);
  VN1690_in1 <= VN_sign_in(10141) & VN_data_in(10141);
  VN1690_in2 <= VN_sign_in(10142) & VN_data_in(10142);
  VN1690_in3 <= VN_sign_in(10143) & VN_data_in(10143);
  VN1690_in4 <= VN_sign_in(10144) & VN_data_in(10144);
  VN1690_in5 <= VN_sign_in(10145) & VN_data_in(10145);
  VN1691_in0 <= VN_sign_in(10146) & VN_data_in(10146);
  VN1691_in1 <= VN_sign_in(10147) & VN_data_in(10147);
  VN1691_in2 <= VN_sign_in(10148) & VN_data_in(10148);
  VN1691_in3 <= VN_sign_in(10149) & VN_data_in(10149);
  VN1691_in4 <= VN_sign_in(10150) & VN_data_in(10150);
  VN1691_in5 <= VN_sign_in(10151) & VN_data_in(10151);
  VN1692_in0 <= VN_sign_in(10152) & VN_data_in(10152);
  VN1692_in1 <= VN_sign_in(10153) & VN_data_in(10153);
  VN1692_in2 <= VN_sign_in(10154) & VN_data_in(10154);
  VN1692_in3 <= VN_sign_in(10155) & VN_data_in(10155);
  VN1692_in4 <= VN_sign_in(10156) & VN_data_in(10156);
  VN1692_in5 <= VN_sign_in(10157) & VN_data_in(10157);
  VN1693_in0 <= VN_sign_in(10158) & VN_data_in(10158);
  VN1693_in1 <= VN_sign_in(10159) & VN_data_in(10159);
  VN1693_in2 <= VN_sign_in(10160) & VN_data_in(10160);
  VN1693_in3 <= VN_sign_in(10161) & VN_data_in(10161);
  VN1693_in4 <= VN_sign_in(10162) & VN_data_in(10162);
  VN1693_in5 <= VN_sign_in(10163) & VN_data_in(10163);
  VN1694_in0 <= VN_sign_in(10164) & VN_data_in(10164);
  VN1694_in1 <= VN_sign_in(10165) & VN_data_in(10165);
  VN1694_in2 <= VN_sign_in(10166) & VN_data_in(10166);
  VN1694_in3 <= VN_sign_in(10167) & VN_data_in(10167);
  VN1694_in4 <= VN_sign_in(10168) & VN_data_in(10168);
  VN1694_in5 <= VN_sign_in(10169) & VN_data_in(10169);
  VN1695_in0 <= VN_sign_in(10170) & VN_data_in(10170);
  VN1695_in1 <= VN_sign_in(10171) & VN_data_in(10171);
  VN1695_in2 <= VN_sign_in(10172) & VN_data_in(10172);
  VN1695_in3 <= VN_sign_in(10173) & VN_data_in(10173);
  VN1695_in4 <= VN_sign_in(10174) & VN_data_in(10174);
  VN1695_in5 <= VN_sign_in(10175) & VN_data_in(10175);
  VN1696_in0 <= VN_sign_in(10176) & VN_data_in(10176);
  VN1696_in1 <= VN_sign_in(10177) & VN_data_in(10177);
  VN1696_in2 <= VN_sign_in(10178) & VN_data_in(10178);
  VN1696_in3 <= VN_sign_in(10179) & VN_data_in(10179);
  VN1696_in4 <= VN_sign_in(10180) & VN_data_in(10180);
  VN1696_in5 <= VN_sign_in(10181) & VN_data_in(10181);
  VN1697_in0 <= VN_sign_in(10182) & VN_data_in(10182);
  VN1697_in1 <= VN_sign_in(10183) & VN_data_in(10183);
  VN1697_in2 <= VN_sign_in(10184) & VN_data_in(10184);
  VN1697_in3 <= VN_sign_in(10185) & VN_data_in(10185);
  VN1697_in4 <= VN_sign_in(10186) & VN_data_in(10186);
  VN1697_in5 <= VN_sign_in(10187) & VN_data_in(10187);
  VN1698_in0 <= VN_sign_in(10188) & VN_data_in(10188);
  VN1698_in1 <= VN_sign_in(10189) & VN_data_in(10189);
  VN1698_in2 <= VN_sign_in(10190) & VN_data_in(10190);
  VN1698_in3 <= VN_sign_in(10191) & VN_data_in(10191);
  VN1698_in4 <= VN_sign_in(10192) & VN_data_in(10192);
  VN1698_in5 <= VN_sign_in(10193) & VN_data_in(10193);
  VN1699_in0 <= VN_sign_in(10194) & VN_data_in(10194);
  VN1699_in1 <= VN_sign_in(10195) & VN_data_in(10195);
  VN1699_in2 <= VN_sign_in(10196) & VN_data_in(10196);
  VN1699_in3 <= VN_sign_in(10197) & VN_data_in(10197);
  VN1699_in4 <= VN_sign_in(10198) & VN_data_in(10198);
  VN1699_in5 <= VN_sign_in(10199) & VN_data_in(10199);
  VN1700_in0 <= VN_sign_in(10200) & VN_data_in(10200);
  VN1700_in1 <= VN_sign_in(10201) & VN_data_in(10201);
  VN1700_in2 <= VN_sign_in(10202) & VN_data_in(10202);
  VN1700_in3 <= VN_sign_in(10203) & VN_data_in(10203);
  VN1700_in4 <= VN_sign_in(10204) & VN_data_in(10204);
  VN1700_in5 <= VN_sign_in(10205) & VN_data_in(10205);
  VN1701_in0 <= VN_sign_in(10206) & VN_data_in(10206);
  VN1701_in1 <= VN_sign_in(10207) & VN_data_in(10207);
  VN1701_in2 <= VN_sign_in(10208) & VN_data_in(10208);
  VN1701_in3 <= VN_sign_in(10209) & VN_data_in(10209);
  VN1701_in4 <= VN_sign_in(10210) & VN_data_in(10210);
  VN1701_in5 <= VN_sign_in(10211) & VN_data_in(10211);
  VN1702_in0 <= VN_sign_in(10212) & VN_data_in(10212);
  VN1702_in1 <= VN_sign_in(10213) & VN_data_in(10213);
  VN1702_in2 <= VN_sign_in(10214) & VN_data_in(10214);
  VN1702_in3 <= VN_sign_in(10215) & VN_data_in(10215);
  VN1702_in4 <= VN_sign_in(10216) & VN_data_in(10216);
  VN1702_in5 <= VN_sign_in(10217) & VN_data_in(10217);
  VN1703_in0 <= VN_sign_in(10218) & VN_data_in(10218);
  VN1703_in1 <= VN_sign_in(10219) & VN_data_in(10219);
  VN1703_in2 <= VN_sign_in(10220) & VN_data_in(10220);
  VN1703_in3 <= VN_sign_in(10221) & VN_data_in(10221);
  VN1703_in4 <= VN_sign_in(10222) & VN_data_in(10222);
  VN1703_in5 <= VN_sign_in(10223) & VN_data_in(10223);
  VN1704_in0 <= VN_sign_in(10224) & VN_data_in(10224);
  VN1704_in1 <= VN_sign_in(10225) & VN_data_in(10225);
  VN1704_in2 <= VN_sign_in(10226) & VN_data_in(10226);
  VN1704_in3 <= VN_sign_in(10227) & VN_data_in(10227);
  VN1704_in4 <= VN_sign_in(10228) & VN_data_in(10228);
  VN1704_in5 <= VN_sign_in(10229) & VN_data_in(10229);
  VN1705_in0 <= VN_sign_in(10230) & VN_data_in(10230);
  VN1705_in1 <= VN_sign_in(10231) & VN_data_in(10231);
  VN1705_in2 <= VN_sign_in(10232) & VN_data_in(10232);
  VN1705_in3 <= VN_sign_in(10233) & VN_data_in(10233);
  VN1705_in4 <= VN_sign_in(10234) & VN_data_in(10234);
  VN1705_in5 <= VN_sign_in(10235) & VN_data_in(10235);
  VN1706_in0 <= VN_sign_in(10236) & VN_data_in(10236);
  VN1706_in1 <= VN_sign_in(10237) & VN_data_in(10237);
  VN1706_in2 <= VN_sign_in(10238) & VN_data_in(10238);
  VN1706_in3 <= VN_sign_in(10239) & VN_data_in(10239);
  VN1706_in4 <= VN_sign_in(10240) & VN_data_in(10240);
  VN1706_in5 <= VN_sign_in(10241) & VN_data_in(10241);
  VN1707_in0 <= VN_sign_in(10242) & VN_data_in(10242);
  VN1707_in1 <= VN_sign_in(10243) & VN_data_in(10243);
  VN1707_in2 <= VN_sign_in(10244) & VN_data_in(10244);
  VN1707_in3 <= VN_sign_in(10245) & VN_data_in(10245);
  VN1707_in4 <= VN_sign_in(10246) & VN_data_in(10246);
  VN1707_in5 <= VN_sign_in(10247) & VN_data_in(10247);
  VN1708_in0 <= VN_sign_in(10248) & VN_data_in(10248);
  VN1708_in1 <= VN_sign_in(10249) & VN_data_in(10249);
  VN1708_in2 <= VN_sign_in(10250) & VN_data_in(10250);
  VN1708_in3 <= VN_sign_in(10251) & VN_data_in(10251);
  VN1708_in4 <= VN_sign_in(10252) & VN_data_in(10252);
  VN1708_in5 <= VN_sign_in(10253) & VN_data_in(10253);
  VN1709_in0 <= VN_sign_in(10254) & VN_data_in(10254);
  VN1709_in1 <= VN_sign_in(10255) & VN_data_in(10255);
  VN1709_in2 <= VN_sign_in(10256) & VN_data_in(10256);
  VN1709_in3 <= VN_sign_in(10257) & VN_data_in(10257);
  VN1709_in4 <= VN_sign_in(10258) & VN_data_in(10258);
  VN1709_in5 <= VN_sign_in(10259) & VN_data_in(10259);
  VN1710_in0 <= VN_sign_in(10260) & VN_data_in(10260);
  VN1710_in1 <= VN_sign_in(10261) & VN_data_in(10261);
  VN1710_in2 <= VN_sign_in(10262) & VN_data_in(10262);
  VN1710_in3 <= VN_sign_in(10263) & VN_data_in(10263);
  VN1710_in4 <= VN_sign_in(10264) & VN_data_in(10264);
  VN1710_in5 <= VN_sign_in(10265) & VN_data_in(10265);
  VN1711_in0 <= VN_sign_in(10266) & VN_data_in(10266);
  VN1711_in1 <= VN_sign_in(10267) & VN_data_in(10267);
  VN1711_in2 <= VN_sign_in(10268) & VN_data_in(10268);
  VN1711_in3 <= VN_sign_in(10269) & VN_data_in(10269);
  VN1711_in4 <= VN_sign_in(10270) & VN_data_in(10270);
  VN1711_in5 <= VN_sign_in(10271) & VN_data_in(10271);
  VN1712_in0 <= VN_sign_in(10272) & VN_data_in(10272);
  VN1712_in1 <= VN_sign_in(10273) & VN_data_in(10273);
  VN1712_in2 <= VN_sign_in(10274) & VN_data_in(10274);
  VN1712_in3 <= VN_sign_in(10275) & VN_data_in(10275);
  VN1712_in4 <= VN_sign_in(10276) & VN_data_in(10276);
  VN1712_in5 <= VN_sign_in(10277) & VN_data_in(10277);
  VN1713_in0 <= VN_sign_in(10278) & VN_data_in(10278);
  VN1713_in1 <= VN_sign_in(10279) & VN_data_in(10279);
  VN1713_in2 <= VN_sign_in(10280) & VN_data_in(10280);
  VN1713_in3 <= VN_sign_in(10281) & VN_data_in(10281);
  VN1713_in4 <= VN_sign_in(10282) & VN_data_in(10282);
  VN1713_in5 <= VN_sign_in(10283) & VN_data_in(10283);
  VN1714_in0 <= VN_sign_in(10284) & VN_data_in(10284);
  VN1714_in1 <= VN_sign_in(10285) & VN_data_in(10285);
  VN1714_in2 <= VN_sign_in(10286) & VN_data_in(10286);
  VN1714_in3 <= VN_sign_in(10287) & VN_data_in(10287);
  VN1714_in4 <= VN_sign_in(10288) & VN_data_in(10288);
  VN1714_in5 <= VN_sign_in(10289) & VN_data_in(10289);
  VN1715_in0 <= VN_sign_in(10290) & VN_data_in(10290);
  VN1715_in1 <= VN_sign_in(10291) & VN_data_in(10291);
  VN1715_in2 <= VN_sign_in(10292) & VN_data_in(10292);
  VN1715_in3 <= VN_sign_in(10293) & VN_data_in(10293);
  VN1715_in4 <= VN_sign_in(10294) & VN_data_in(10294);
  VN1715_in5 <= VN_sign_in(10295) & VN_data_in(10295);
  VN1716_in0 <= VN_sign_in(10296) & VN_data_in(10296);
  VN1716_in1 <= VN_sign_in(10297) & VN_data_in(10297);
  VN1716_in2 <= VN_sign_in(10298) & VN_data_in(10298);
  VN1716_in3 <= VN_sign_in(10299) & VN_data_in(10299);
  VN1716_in4 <= VN_sign_in(10300) & VN_data_in(10300);
  VN1716_in5 <= VN_sign_in(10301) & VN_data_in(10301);
  VN1717_in0 <= VN_sign_in(10302) & VN_data_in(10302);
  VN1717_in1 <= VN_sign_in(10303) & VN_data_in(10303);
  VN1717_in2 <= VN_sign_in(10304) & VN_data_in(10304);
  VN1717_in3 <= VN_sign_in(10305) & VN_data_in(10305);
  VN1717_in4 <= VN_sign_in(10306) & VN_data_in(10306);
  VN1717_in5 <= VN_sign_in(10307) & VN_data_in(10307);
  VN1718_in0 <= VN_sign_in(10308) & VN_data_in(10308);
  VN1718_in1 <= VN_sign_in(10309) & VN_data_in(10309);
  VN1718_in2 <= VN_sign_in(10310) & VN_data_in(10310);
  VN1718_in3 <= VN_sign_in(10311) & VN_data_in(10311);
  VN1718_in4 <= VN_sign_in(10312) & VN_data_in(10312);
  VN1718_in5 <= VN_sign_in(10313) & VN_data_in(10313);
  VN1719_in0 <= VN_sign_in(10314) & VN_data_in(10314);
  VN1719_in1 <= VN_sign_in(10315) & VN_data_in(10315);
  VN1719_in2 <= VN_sign_in(10316) & VN_data_in(10316);
  VN1719_in3 <= VN_sign_in(10317) & VN_data_in(10317);
  VN1719_in4 <= VN_sign_in(10318) & VN_data_in(10318);
  VN1719_in5 <= VN_sign_in(10319) & VN_data_in(10319);
  VN1720_in0 <= VN_sign_in(10320) & VN_data_in(10320);
  VN1720_in1 <= VN_sign_in(10321) & VN_data_in(10321);
  VN1720_in2 <= VN_sign_in(10322) & VN_data_in(10322);
  VN1720_in3 <= VN_sign_in(10323) & VN_data_in(10323);
  VN1720_in4 <= VN_sign_in(10324) & VN_data_in(10324);
  VN1720_in5 <= VN_sign_in(10325) & VN_data_in(10325);
  VN1721_in0 <= VN_sign_in(10326) & VN_data_in(10326);
  VN1721_in1 <= VN_sign_in(10327) & VN_data_in(10327);
  VN1721_in2 <= VN_sign_in(10328) & VN_data_in(10328);
  VN1721_in3 <= VN_sign_in(10329) & VN_data_in(10329);
  VN1721_in4 <= VN_sign_in(10330) & VN_data_in(10330);
  VN1721_in5 <= VN_sign_in(10331) & VN_data_in(10331);
  VN1722_in0 <= VN_sign_in(10332) & VN_data_in(10332);
  VN1722_in1 <= VN_sign_in(10333) & VN_data_in(10333);
  VN1722_in2 <= VN_sign_in(10334) & VN_data_in(10334);
  VN1722_in3 <= VN_sign_in(10335) & VN_data_in(10335);
  VN1722_in4 <= VN_sign_in(10336) & VN_data_in(10336);
  VN1722_in5 <= VN_sign_in(10337) & VN_data_in(10337);
  VN1723_in0 <= VN_sign_in(10338) & VN_data_in(10338);
  VN1723_in1 <= VN_sign_in(10339) & VN_data_in(10339);
  VN1723_in2 <= VN_sign_in(10340) & VN_data_in(10340);
  VN1723_in3 <= VN_sign_in(10341) & VN_data_in(10341);
  VN1723_in4 <= VN_sign_in(10342) & VN_data_in(10342);
  VN1723_in5 <= VN_sign_in(10343) & VN_data_in(10343);
  VN1724_in0 <= VN_sign_in(10344) & VN_data_in(10344);
  VN1724_in1 <= VN_sign_in(10345) & VN_data_in(10345);
  VN1724_in2 <= VN_sign_in(10346) & VN_data_in(10346);
  VN1724_in3 <= VN_sign_in(10347) & VN_data_in(10347);
  VN1724_in4 <= VN_sign_in(10348) & VN_data_in(10348);
  VN1724_in5 <= VN_sign_in(10349) & VN_data_in(10349);
  VN1725_in0 <= VN_sign_in(10350) & VN_data_in(10350);
  VN1725_in1 <= VN_sign_in(10351) & VN_data_in(10351);
  VN1725_in2 <= VN_sign_in(10352) & VN_data_in(10352);
  VN1725_in3 <= VN_sign_in(10353) & VN_data_in(10353);
  VN1725_in4 <= VN_sign_in(10354) & VN_data_in(10354);
  VN1725_in5 <= VN_sign_in(10355) & VN_data_in(10355);
  VN1726_in0 <= VN_sign_in(10356) & VN_data_in(10356);
  VN1726_in1 <= VN_sign_in(10357) & VN_data_in(10357);
  VN1726_in2 <= VN_sign_in(10358) & VN_data_in(10358);
  VN1726_in3 <= VN_sign_in(10359) & VN_data_in(10359);
  VN1726_in4 <= VN_sign_in(10360) & VN_data_in(10360);
  VN1726_in5 <= VN_sign_in(10361) & VN_data_in(10361);
  VN1727_in0 <= VN_sign_in(10362) & VN_data_in(10362);
  VN1727_in1 <= VN_sign_in(10363) & VN_data_in(10363);
  VN1727_in2 <= VN_sign_in(10364) & VN_data_in(10364);
  VN1727_in3 <= VN_sign_in(10365) & VN_data_in(10365);
  VN1727_in4 <= VN_sign_in(10366) & VN_data_in(10366);
  VN1727_in5 <= VN_sign_in(10367) & VN_data_in(10367);
  VN1728_in0 <= VN_sign_in(10368) & VN_data_in(10368);
  VN1728_in1 <= VN_sign_in(10369) & VN_data_in(10369);
  VN1728_in2 <= VN_sign_in(10370) & VN_data_in(10370);
  VN1728_in3 <= VN_sign_in(10371) & VN_data_in(10371);
  VN1728_in4 <= VN_sign_in(10372) & VN_data_in(10372);
  VN1728_in5 <= VN_sign_in(10373) & VN_data_in(10373);
  VN1729_in0 <= VN_sign_in(10374) & VN_data_in(10374);
  VN1729_in1 <= VN_sign_in(10375) & VN_data_in(10375);
  VN1729_in2 <= VN_sign_in(10376) & VN_data_in(10376);
  VN1729_in3 <= VN_sign_in(10377) & VN_data_in(10377);
  VN1729_in4 <= VN_sign_in(10378) & VN_data_in(10378);
  VN1729_in5 <= VN_sign_in(10379) & VN_data_in(10379);
  VN1730_in0 <= VN_sign_in(10380) & VN_data_in(10380);
  VN1730_in1 <= VN_sign_in(10381) & VN_data_in(10381);
  VN1730_in2 <= VN_sign_in(10382) & VN_data_in(10382);
  VN1730_in3 <= VN_sign_in(10383) & VN_data_in(10383);
  VN1730_in4 <= VN_sign_in(10384) & VN_data_in(10384);
  VN1730_in5 <= VN_sign_in(10385) & VN_data_in(10385);
  VN1731_in0 <= VN_sign_in(10386) & VN_data_in(10386);
  VN1731_in1 <= VN_sign_in(10387) & VN_data_in(10387);
  VN1731_in2 <= VN_sign_in(10388) & VN_data_in(10388);
  VN1731_in3 <= VN_sign_in(10389) & VN_data_in(10389);
  VN1731_in4 <= VN_sign_in(10390) & VN_data_in(10390);
  VN1731_in5 <= VN_sign_in(10391) & VN_data_in(10391);
  VN1732_in0 <= VN_sign_in(10392) & VN_data_in(10392);
  VN1732_in1 <= VN_sign_in(10393) & VN_data_in(10393);
  VN1732_in2 <= VN_sign_in(10394) & VN_data_in(10394);
  VN1732_in3 <= VN_sign_in(10395) & VN_data_in(10395);
  VN1732_in4 <= VN_sign_in(10396) & VN_data_in(10396);
  VN1732_in5 <= VN_sign_in(10397) & VN_data_in(10397);
  VN1733_in0 <= VN_sign_in(10398) & VN_data_in(10398);
  VN1733_in1 <= VN_sign_in(10399) & VN_data_in(10399);
  VN1733_in2 <= VN_sign_in(10400) & VN_data_in(10400);
  VN1733_in3 <= VN_sign_in(10401) & VN_data_in(10401);
  VN1733_in4 <= VN_sign_in(10402) & VN_data_in(10402);
  VN1733_in5 <= VN_sign_in(10403) & VN_data_in(10403);
  VN1734_in0 <= VN_sign_in(10404) & VN_data_in(10404);
  VN1734_in1 <= VN_sign_in(10405) & VN_data_in(10405);
  VN1734_in2 <= VN_sign_in(10406) & VN_data_in(10406);
  VN1734_in3 <= VN_sign_in(10407) & VN_data_in(10407);
  VN1734_in4 <= VN_sign_in(10408) & VN_data_in(10408);
  VN1734_in5 <= VN_sign_in(10409) & VN_data_in(10409);
  VN1735_in0 <= VN_sign_in(10410) & VN_data_in(10410);
  VN1735_in1 <= VN_sign_in(10411) & VN_data_in(10411);
  VN1735_in2 <= VN_sign_in(10412) & VN_data_in(10412);
  VN1735_in3 <= VN_sign_in(10413) & VN_data_in(10413);
  VN1735_in4 <= VN_sign_in(10414) & VN_data_in(10414);
  VN1735_in5 <= VN_sign_in(10415) & VN_data_in(10415);
  VN1736_in0 <= VN_sign_in(10416) & VN_data_in(10416);
  VN1736_in1 <= VN_sign_in(10417) & VN_data_in(10417);
  VN1736_in2 <= VN_sign_in(10418) & VN_data_in(10418);
  VN1736_in3 <= VN_sign_in(10419) & VN_data_in(10419);
  VN1736_in4 <= VN_sign_in(10420) & VN_data_in(10420);
  VN1736_in5 <= VN_sign_in(10421) & VN_data_in(10421);
  VN1737_in0 <= VN_sign_in(10422) & VN_data_in(10422);
  VN1737_in1 <= VN_sign_in(10423) & VN_data_in(10423);
  VN1737_in2 <= VN_sign_in(10424) & VN_data_in(10424);
  VN1737_in3 <= VN_sign_in(10425) & VN_data_in(10425);
  VN1737_in4 <= VN_sign_in(10426) & VN_data_in(10426);
  VN1737_in5 <= VN_sign_in(10427) & VN_data_in(10427);
  VN1738_in0 <= VN_sign_in(10428) & VN_data_in(10428);
  VN1738_in1 <= VN_sign_in(10429) & VN_data_in(10429);
  VN1738_in2 <= VN_sign_in(10430) & VN_data_in(10430);
  VN1738_in3 <= VN_sign_in(10431) & VN_data_in(10431);
  VN1738_in4 <= VN_sign_in(10432) & VN_data_in(10432);
  VN1738_in5 <= VN_sign_in(10433) & VN_data_in(10433);
  VN1739_in0 <= VN_sign_in(10434) & VN_data_in(10434);
  VN1739_in1 <= VN_sign_in(10435) & VN_data_in(10435);
  VN1739_in2 <= VN_sign_in(10436) & VN_data_in(10436);
  VN1739_in3 <= VN_sign_in(10437) & VN_data_in(10437);
  VN1739_in4 <= VN_sign_in(10438) & VN_data_in(10438);
  VN1739_in5 <= VN_sign_in(10439) & VN_data_in(10439);
  VN1740_in0 <= VN_sign_in(10440) & VN_data_in(10440);
  VN1740_in1 <= VN_sign_in(10441) & VN_data_in(10441);
  VN1740_in2 <= VN_sign_in(10442) & VN_data_in(10442);
  VN1740_in3 <= VN_sign_in(10443) & VN_data_in(10443);
  VN1740_in4 <= VN_sign_in(10444) & VN_data_in(10444);
  VN1740_in5 <= VN_sign_in(10445) & VN_data_in(10445);
  VN1741_in0 <= VN_sign_in(10446) & VN_data_in(10446);
  VN1741_in1 <= VN_sign_in(10447) & VN_data_in(10447);
  VN1741_in2 <= VN_sign_in(10448) & VN_data_in(10448);
  VN1741_in3 <= VN_sign_in(10449) & VN_data_in(10449);
  VN1741_in4 <= VN_sign_in(10450) & VN_data_in(10450);
  VN1741_in5 <= VN_sign_in(10451) & VN_data_in(10451);
  VN1742_in0 <= VN_sign_in(10452) & VN_data_in(10452);
  VN1742_in1 <= VN_sign_in(10453) & VN_data_in(10453);
  VN1742_in2 <= VN_sign_in(10454) & VN_data_in(10454);
  VN1742_in3 <= VN_sign_in(10455) & VN_data_in(10455);
  VN1742_in4 <= VN_sign_in(10456) & VN_data_in(10456);
  VN1742_in5 <= VN_sign_in(10457) & VN_data_in(10457);
  VN1743_in0 <= VN_sign_in(10458) & VN_data_in(10458);
  VN1743_in1 <= VN_sign_in(10459) & VN_data_in(10459);
  VN1743_in2 <= VN_sign_in(10460) & VN_data_in(10460);
  VN1743_in3 <= VN_sign_in(10461) & VN_data_in(10461);
  VN1743_in4 <= VN_sign_in(10462) & VN_data_in(10462);
  VN1743_in5 <= VN_sign_in(10463) & VN_data_in(10463);
  VN1744_in0 <= VN_sign_in(10464) & VN_data_in(10464);
  VN1744_in1 <= VN_sign_in(10465) & VN_data_in(10465);
  VN1744_in2 <= VN_sign_in(10466) & VN_data_in(10466);
  VN1744_in3 <= VN_sign_in(10467) & VN_data_in(10467);
  VN1744_in4 <= VN_sign_in(10468) & VN_data_in(10468);
  VN1744_in5 <= VN_sign_in(10469) & VN_data_in(10469);
  VN1745_in0 <= VN_sign_in(10470) & VN_data_in(10470);
  VN1745_in1 <= VN_sign_in(10471) & VN_data_in(10471);
  VN1745_in2 <= VN_sign_in(10472) & VN_data_in(10472);
  VN1745_in3 <= VN_sign_in(10473) & VN_data_in(10473);
  VN1745_in4 <= VN_sign_in(10474) & VN_data_in(10474);
  VN1745_in5 <= VN_sign_in(10475) & VN_data_in(10475);
  VN1746_in0 <= VN_sign_in(10476) & VN_data_in(10476);
  VN1746_in1 <= VN_sign_in(10477) & VN_data_in(10477);
  VN1746_in2 <= VN_sign_in(10478) & VN_data_in(10478);
  VN1746_in3 <= VN_sign_in(10479) & VN_data_in(10479);
  VN1746_in4 <= VN_sign_in(10480) & VN_data_in(10480);
  VN1746_in5 <= VN_sign_in(10481) & VN_data_in(10481);
  VN1747_in0 <= VN_sign_in(10482) & VN_data_in(10482);
  VN1747_in1 <= VN_sign_in(10483) & VN_data_in(10483);
  VN1747_in2 <= VN_sign_in(10484) & VN_data_in(10484);
  VN1747_in3 <= VN_sign_in(10485) & VN_data_in(10485);
  VN1747_in4 <= VN_sign_in(10486) & VN_data_in(10486);
  VN1747_in5 <= VN_sign_in(10487) & VN_data_in(10487);
  VN1748_in0 <= VN_sign_in(10488) & VN_data_in(10488);
  VN1748_in1 <= VN_sign_in(10489) & VN_data_in(10489);
  VN1748_in2 <= VN_sign_in(10490) & VN_data_in(10490);
  VN1748_in3 <= VN_sign_in(10491) & VN_data_in(10491);
  VN1748_in4 <= VN_sign_in(10492) & VN_data_in(10492);
  VN1748_in5 <= VN_sign_in(10493) & VN_data_in(10493);
  VN1749_in0 <= VN_sign_in(10494) & VN_data_in(10494);
  VN1749_in1 <= VN_sign_in(10495) & VN_data_in(10495);
  VN1749_in2 <= VN_sign_in(10496) & VN_data_in(10496);
  VN1749_in3 <= VN_sign_in(10497) & VN_data_in(10497);
  VN1749_in4 <= VN_sign_in(10498) & VN_data_in(10498);
  VN1749_in5 <= VN_sign_in(10499) & VN_data_in(10499);
  VN1750_in0 <= VN_sign_in(10500) & VN_data_in(10500);
  VN1750_in1 <= VN_sign_in(10501) & VN_data_in(10501);
  VN1750_in2 <= VN_sign_in(10502) & VN_data_in(10502);
  VN1750_in3 <= VN_sign_in(10503) & VN_data_in(10503);
  VN1750_in4 <= VN_sign_in(10504) & VN_data_in(10504);
  VN1750_in5 <= VN_sign_in(10505) & VN_data_in(10505);
  VN1751_in0 <= VN_sign_in(10506) & VN_data_in(10506);
  VN1751_in1 <= VN_sign_in(10507) & VN_data_in(10507);
  VN1751_in2 <= VN_sign_in(10508) & VN_data_in(10508);
  VN1751_in3 <= VN_sign_in(10509) & VN_data_in(10509);
  VN1751_in4 <= VN_sign_in(10510) & VN_data_in(10510);
  VN1751_in5 <= VN_sign_in(10511) & VN_data_in(10511);
  VN1752_in0 <= VN_sign_in(10512) & VN_data_in(10512);
  VN1752_in1 <= VN_sign_in(10513) & VN_data_in(10513);
  VN1752_in2 <= VN_sign_in(10514) & VN_data_in(10514);
  VN1752_in3 <= VN_sign_in(10515) & VN_data_in(10515);
  VN1752_in4 <= VN_sign_in(10516) & VN_data_in(10516);
  VN1752_in5 <= VN_sign_in(10517) & VN_data_in(10517);
  VN1753_in0 <= VN_sign_in(10518) & VN_data_in(10518);
  VN1753_in1 <= VN_sign_in(10519) & VN_data_in(10519);
  VN1753_in2 <= VN_sign_in(10520) & VN_data_in(10520);
  VN1753_in3 <= VN_sign_in(10521) & VN_data_in(10521);
  VN1753_in4 <= VN_sign_in(10522) & VN_data_in(10522);
  VN1753_in5 <= VN_sign_in(10523) & VN_data_in(10523);
  VN1754_in0 <= VN_sign_in(10524) & VN_data_in(10524);
  VN1754_in1 <= VN_sign_in(10525) & VN_data_in(10525);
  VN1754_in2 <= VN_sign_in(10526) & VN_data_in(10526);
  VN1754_in3 <= VN_sign_in(10527) & VN_data_in(10527);
  VN1754_in4 <= VN_sign_in(10528) & VN_data_in(10528);
  VN1754_in5 <= VN_sign_in(10529) & VN_data_in(10529);
  VN1755_in0 <= VN_sign_in(10530) & VN_data_in(10530);
  VN1755_in1 <= VN_sign_in(10531) & VN_data_in(10531);
  VN1755_in2 <= VN_sign_in(10532) & VN_data_in(10532);
  VN1755_in3 <= VN_sign_in(10533) & VN_data_in(10533);
  VN1755_in4 <= VN_sign_in(10534) & VN_data_in(10534);
  VN1755_in5 <= VN_sign_in(10535) & VN_data_in(10535);
  VN1756_in0 <= VN_sign_in(10536) & VN_data_in(10536);
  VN1756_in1 <= VN_sign_in(10537) & VN_data_in(10537);
  VN1756_in2 <= VN_sign_in(10538) & VN_data_in(10538);
  VN1756_in3 <= VN_sign_in(10539) & VN_data_in(10539);
  VN1756_in4 <= VN_sign_in(10540) & VN_data_in(10540);
  VN1756_in5 <= VN_sign_in(10541) & VN_data_in(10541);
  VN1757_in0 <= VN_sign_in(10542) & VN_data_in(10542);
  VN1757_in1 <= VN_sign_in(10543) & VN_data_in(10543);
  VN1757_in2 <= VN_sign_in(10544) & VN_data_in(10544);
  VN1757_in3 <= VN_sign_in(10545) & VN_data_in(10545);
  VN1757_in4 <= VN_sign_in(10546) & VN_data_in(10546);
  VN1757_in5 <= VN_sign_in(10547) & VN_data_in(10547);
  VN1758_in0 <= VN_sign_in(10548) & VN_data_in(10548);
  VN1758_in1 <= VN_sign_in(10549) & VN_data_in(10549);
  VN1758_in2 <= VN_sign_in(10550) & VN_data_in(10550);
  VN1758_in3 <= VN_sign_in(10551) & VN_data_in(10551);
  VN1758_in4 <= VN_sign_in(10552) & VN_data_in(10552);
  VN1758_in5 <= VN_sign_in(10553) & VN_data_in(10553);
  VN1759_in0 <= VN_sign_in(10554) & VN_data_in(10554);
  VN1759_in1 <= VN_sign_in(10555) & VN_data_in(10555);
  VN1759_in2 <= VN_sign_in(10556) & VN_data_in(10556);
  VN1759_in3 <= VN_sign_in(10557) & VN_data_in(10557);
  VN1759_in4 <= VN_sign_in(10558) & VN_data_in(10558);
  VN1759_in5 <= VN_sign_in(10559) & VN_data_in(10559);
  VN1760_in0 <= VN_sign_in(10560) & VN_data_in(10560);
  VN1760_in1 <= VN_sign_in(10561) & VN_data_in(10561);
  VN1760_in2 <= VN_sign_in(10562) & VN_data_in(10562);
  VN1760_in3 <= VN_sign_in(10563) & VN_data_in(10563);
  VN1760_in4 <= VN_sign_in(10564) & VN_data_in(10564);
  VN1760_in5 <= VN_sign_in(10565) & VN_data_in(10565);
  VN1761_in0 <= VN_sign_in(10566) & VN_data_in(10566);
  VN1761_in1 <= VN_sign_in(10567) & VN_data_in(10567);
  VN1761_in2 <= VN_sign_in(10568) & VN_data_in(10568);
  VN1761_in3 <= VN_sign_in(10569) & VN_data_in(10569);
  VN1761_in4 <= VN_sign_in(10570) & VN_data_in(10570);
  VN1761_in5 <= VN_sign_in(10571) & VN_data_in(10571);
  VN1762_in0 <= VN_sign_in(10572) & VN_data_in(10572);
  VN1762_in1 <= VN_sign_in(10573) & VN_data_in(10573);
  VN1762_in2 <= VN_sign_in(10574) & VN_data_in(10574);
  VN1762_in3 <= VN_sign_in(10575) & VN_data_in(10575);
  VN1762_in4 <= VN_sign_in(10576) & VN_data_in(10576);
  VN1762_in5 <= VN_sign_in(10577) & VN_data_in(10577);
  VN1763_in0 <= VN_sign_in(10578) & VN_data_in(10578);
  VN1763_in1 <= VN_sign_in(10579) & VN_data_in(10579);
  VN1763_in2 <= VN_sign_in(10580) & VN_data_in(10580);
  VN1763_in3 <= VN_sign_in(10581) & VN_data_in(10581);
  VN1763_in4 <= VN_sign_in(10582) & VN_data_in(10582);
  VN1763_in5 <= VN_sign_in(10583) & VN_data_in(10583);
  VN1764_in0 <= VN_sign_in(10584) & VN_data_in(10584);
  VN1764_in1 <= VN_sign_in(10585) & VN_data_in(10585);
  VN1764_in2 <= VN_sign_in(10586) & VN_data_in(10586);
  VN1764_in3 <= VN_sign_in(10587) & VN_data_in(10587);
  VN1764_in4 <= VN_sign_in(10588) & VN_data_in(10588);
  VN1764_in5 <= VN_sign_in(10589) & VN_data_in(10589);
  VN1765_in0 <= VN_sign_in(10590) & VN_data_in(10590);
  VN1765_in1 <= VN_sign_in(10591) & VN_data_in(10591);
  VN1765_in2 <= VN_sign_in(10592) & VN_data_in(10592);
  VN1765_in3 <= VN_sign_in(10593) & VN_data_in(10593);
  VN1765_in4 <= VN_sign_in(10594) & VN_data_in(10594);
  VN1765_in5 <= VN_sign_in(10595) & VN_data_in(10595);
  VN1766_in0 <= VN_sign_in(10596) & VN_data_in(10596);
  VN1766_in1 <= VN_sign_in(10597) & VN_data_in(10597);
  VN1766_in2 <= VN_sign_in(10598) & VN_data_in(10598);
  VN1766_in3 <= VN_sign_in(10599) & VN_data_in(10599);
  VN1766_in4 <= VN_sign_in(10600) & VN_data_in(10600);
  VN1766_in5 <= VN_sign_in(10601) & VN_data_in(10601);
  VN1767_in0 <= VN_sign_in(10602) & VN_data_in(10602);
  VN1767_in1 <= VN_sign_in(10603) & VN_data_in(10603);
  VN1767_in2 <= VN_sign_in(10604) & VN_data_in(10604);
  VN1767_in3 <= VN_sign_in(10605) & VN_data_in(10605);
  VN1767_in4 <= VN_sign_in(10606) & VN_data_in(10606);
  VN1767_in5 <= VN_sign_in(10607) & VN_data_in(10607);
  VN1768_in0 <= VN_sign_in(10608) & VN_data_in(10608);
  VN1768_in1 <= VN_sign_in(10609) & VN_data_in(10609);
  VN1768_in2 <= VN_sign_in(10610) & VN_data_in(10610);
  VN1768_in3 <= VN_sign_in(10611) & VN_data_in(10611);
  VN1768_in4 <= VN_sign_in(10612) & VN_data_in(10612);
  VN1768_in5 <= VN_sign_in(10613) & VN_data_in(10613);
  VN1769_in0 <= VN_sign_in(10614) & VN_data_in(10614);
  VN1769_in1 <= VN_sign_in(10615) & VN_data_in(10615);
  VN1769_in2 <= VN_sign_in(10616) & VN_data_in(10616);
  VN1769_in3 <= VN_sign_in(10617) & VN_data_in(10617);
  VN1769_in4 <= VN_sign_in(10618) & VN_data_in(10618);
  VN1769_in5 <= VN_sign_in(10619) & VN_data_in(10619);
  VN1770_in0 <= VN_sign_in(10620) & VN_data_in(10620);
  VN1770_in1 <= VN_sign_in(10621) & VN_data_in(10621);
  VN1770_in2 <= VN_sign_in(10622) & VN_data_in(10622);
  VN1770_in3 <= VN_sign_in(10623) & VN_data_in(10623);
  VN1770_in4 <= VN_sign_in(10624) & VN_data_in(10624);
  VN1770_in5 <= VN_sign_in(10625) & VN_data_in(10625);
  VN1771_in0 <= VN_sign_in(10626) & VN_data_in(10626);
  VN1771_in1 <= VN_sign_in(10627) & VN_data_in(10627);
  VN1771_in2 <= VN_sign_in(10628) & VN_data_in(10628);
  VN1771_in3 <= VN_sign_in(10629) & VN_data_in(10629);
  VN1771_in4 <= VN_sign_in(10630) & VN_data_in(10630);
  VN1771_in5 <= VN_sign_in(10631) & VN_data_in(10631);
  VN1772_in0 <= VN_sign_in(10632) & VN_data_in(10632);
  VN1772_in1 <= VN_sign_in(10633) & VN_data_in(10633);
  VN1772_in2 <= VN_sign_in(10634) & VN_data_in(10634);
  VN1772_in3 <= VN_sign_in(10635) & VN_data_in(10635);
  VN1772_in4 <= VN_sign_in(10636) & VN_data_in(10636);
  VN1772_in5 <= VN_sign_in(10637) & VN_data_in(10637);
  VN1773_in0 <= VN_sign_in(10638) & VN_data_in(10638);
  VN1773_in1 <= VN_sign_in(10639) & VN_data_in(10639);
  VN1773_in2 <= VN_sign_in(10640) & VN_data_in(10640);
  VN1773_in3 <= VN_sign_in(10641) & VN_data_in(10641);
  VN1773_in4 <= VN_sign_in(10642) & VN_data_in(10642);
  VN1773_in5 <= VN_sign_in(10643) & VN_data_in(10643);
  VN1774_in0 <= VN_sign_in(10644) & VN_data_in(10644);
  VN1774_in1 <= VN_sign_in(10645) & VN_data_in(10645);
  VN1774_in2 <= VN_sign_in(10646) & VN_data_in(10646);
  VN1774_in3 <= VN_sign_in(10647) & VN_data_in(10647);
  VN1774_in4 <= VN_sign_in(10648) & VN_data_in(10648);
  VN1774_in5 <= VN_sign_in(10649) & VN_data_in(10649);
  VN1775_in0 <= VN_sign_in(10650) & VN_data_in(10650);
  VN1775_in1 <= VN_sign_in(10651) & VN_data_in(10651);
  VN1775_in2 <= VN_sign_in(10652) & VN_data_in(10652);
  VN1775_in3 <= VN_sign_in(10653) & VN_data_in(10653);
  VN1775_in4 <= VN_sign_in(10654) & VN_data_in(10654);
  VN1775_in5 <= VN_sign_in(10655) & VN_data_in(10655);
  VN1776_in0 <= VN_sign_in(10656) & VN_data_in(10656);
  VN1776_in1 <= VN_sign_in(10657) & VN_data_in(10657);
  VN1776_in2 <= VN_sign_in(10658) & VN_data_in(10658);
  VN1776_in3 <= VN_sign_in(10659) & VN_data_in(10659);
  VN1776_in4 <= VN_sign_in(10660) & VN_data_in(10660);
  VN1776_in5 <= VN_sign_in(10661) & VN_data_in(10661);
  VN1777_in0 <= VN_sign_in(10662) & VN_data_in(10662);
  VN1777_in1 <= VN_sign_in(10663) & VN_data_in(10663);
  VN1777_in2 <= VN_sign_in(10664) & VN_data_in(10664);
  VN1777_in3 <= VN_sign_in(10665) & VN_data_in(10665);
  VN1777_in4 <= VN_sign_in(10666) & VN_data_in(10666);
  VN1777_in5 <= VN_sign_in(10667) & VN_data_in(10667);
  VN1778_in0 <= VN_sign_in(10668) & VN_data_in(10668);
  VN1778_in1 <= VN_sign_in(10669) & VN_data_in(10669);
  VN1778_in2 <= VN_sign_in(10670) & VN_data_in(10670);
  VN1778_in3 <= VN_sign_in(10671) & VN_data_in(10671);
  VN1778_in4 <= VN_sign_in(10672) & VN_data_in(10672);
  VN1778_in5 <= VN_sign_in(10673) & VN_data_in(10673);
  VN1779_in0 <= VN_sign_in(10674) & VN_data_in(10674);
  VN1779_in1 <= VN_sign_in(10675) & VN_data_in(10675);
  VN1779_in2 <= VN_sign_in(10676) & VN_data_in(10676);
  VN1779_in3 <= VN_sign_in(10677) & VN_data_in(10677);
  VN1779_in4 <= VN_sign_in(10678) & VN_data_in(10678);
  VN1779_in5 <= VN_sign_in(10679) & VN_data_in(10679);
  VN1780_in0 <= VN_sign_in(10680) & VN_data_in(10680);
  VN1780_in1 <= VN_sign_in(10681) & VN_data_in(10681);
  VN1780_in2 <= VN_sign_in(10682) & VN_data_in(10682);
  VN1780_in3 <= VN_sign_in(10683) & VN_data_in(10683);
  VN1780_in4 <= VN_sign_in(10684) & VN_data_in(10684);
  VN1780_in5 <= VN_sign_in(10685) & VN_data_in(10685);
  VN1781_in0 <= VN_sign_in(10686) & VN_data_in(10686);
  VN1781_in1 <= VN_sign_in(10687) & VN_data_in(10687);
  VN1781_in2 <= VN_sign_in(10688) & VN_data_in(10688);
  VN1781_in3 <= VN_sign_in(10689) & VN_data_in(10689);
  VN1781_in4 <= VN_sign_in(10690) & VN_data_in(10690);
  VN1781_in5 <= VN_sign_in(10691) & VN_data_in(10691);
  VN1782_in0 <= VN_sign_in(10692) & VN_data_in(10692);
  VN1782_in1 <= VN_sign_in(10693) & VN_data_in(10693);
  VN1782_in2 <= VN_sign_in(10694) & VN_data_in(10694);
  VN1782_in3 <= VN_sign_in(10695) & VN_data_in(10695);
  VN1782_in4 <= VN_sign_in(10696) & VN_data_in(10696);
  VN1782_in5 <= VN_sign_in(10697) & VN_data_in(10697);
  VN1783_in0 <= VN_sign_in(10698) & VN_data_in(10698);
  VN1783_in1 <= VN_sign_in(10699) & VN_data_in(10699);
  VN1783_in2 <= VN_sign_in(10700) & VN_data_in(10700);
  VN1783_in3 <= VN_sign_in(10701) & VN_data_in(10701);
  VN1783_in4 <= VN_sign_in(10702) & VN_data_in(10702);
  VN1783_in5 <= VN_sign_in(10703) & VN_data_in(10703);
  VN1784_in0 <= VN_sign_in(10704) & VN_data_in(10704);
  VN1784_in1 <= VN_sign_in(10705) & VN_data_in(10705);
  VN1784_in2 <= VN_sign_in(10706) & VN_data_in(10706);
  VN1784_in3 <= VN_sign_in(10707) & VN_data_in(10707);
  VN1784_in4 <= VN_sign_in(10708) & VN_data_in(10708);
  VN1784_in5 <= VN_sign_in(10709) & VN_data_in(10709);
  VN1785_in0 <= VN_sign_in(10710) & VN_data_in(10710);
  VN1785_in1 <= VN_sign_in(10711) & VN_data_in(10711);
  VN1785_in2 <= VN_sign_in(10712) & VN_data_in(10712);
  VN1785_in3 <= VN_sign_in(10713) & VN_data_in(10713);
  VN1785_in4 <= VN_sign_in(10714) & VN_data_in(10714);
  VN1785_in5 <= VN_sign_in(10715) & VN_data_in(10715);
  VN1786_in0 <= VN_sign_in(10716) & VN_data_in(10716);
  VN1786_in1 <= VN_sign_in(10717) & VN_data_in(10717);
  VN1786_in2 <= VN_sign_in(10718) & VN_data_in(10718);
  VN1786_in3 <= VN_sign_in(10719) & VN_data_in(10719);
  VN1786_in4 <= VN_sign_in(10720) & VN_data_in(10720);
  VN1786_in5 <= VN_sign_in(10721) & VN_data_in(10721);
  VN1787_in0 <= VN_sign_in(10722) & VN_data_in(10722);
  VN1787_in1 <= VN_sign_in(10723) & VN_data_in(10723);
  VN1787_in2 <= VN_sign_in(10724) & VN_data_in(10724);
  VN1787_in3 <= VN_sign_in(10725) & VN_data_in(10725);
  VN1787_in4 <= VN_sign_in(10726) & VN_data_in(10726);
  VN1787_in5 <= VN_sign_in(10727) & VN_data_in(10727);
  VN1788_in0 <= VN_sign_in(10728) & VN_data_in(10728);
  VN1788_in1 <= VN_sign_in(10729) & VN_data_in(10729);
  VN1788_in2 <= VN_sign_in(10730) & VN_data_in(10730);
  VN1788_in3 <= VN_sign_in(10731) & VN_data_in(10731);
  VN1788_in4 <= VN_sign_in(10732) & VN_data_in(10732);
  VN1788_in5 <= VN_sign_in(10733) & VN_data_in(10733);
  VN1789_in0 <= VN_sign_in(10734) & VN_data_in(10734);
  VN1789_in1 <= VN_sign_in(10735) & VN_data_in(10735);
  VN1789_in2 <= VN_sign_in(10736) & VN_data_in(10736);
  VN1789_in3 <= VN_sign_in(10737) & VN_data_in(10737);
  VN1789_in4 <= VN_sign_in(10738) & VN_data_in(10738);
  VN1789_in5 <= VN_sign_in(10739) & VN_data_in(10739);
  VN1790_in0 <= VN_sign_in(10740) & VN_data_in(10740);
  VN1790_in1 <= VN_sign_in(10741) & VN_data_in(10741);
  VN1790_in2 <= VN_sign_in(10742) & VN_data_in(10742);
  VN1790_in3 <= VN_sign_in(10743) & VN_data_in(10743);
  VN1790_in4 <= VN_sign_in(10744) & VN_data_in(10744);
  VN1790_in5 <= VN_sign_in(10745) & VN_data_in(10745);
  VN1791_in0 <= VN_sign_in(10746) & VN_data_in(10746);
  VN1791_in1 <= VN_sign_in(10747) & VN_data_in(10747);
  VN1791_in2 <= VN_sign_in(10748) & VN_data_in(10748);
  VN1791_in3 <= VN_sign_in(10749) & VN_data_in(10749);
  VN1791_in4 <= VN_sign_in(10750) & VN_data_in(10750);
  VN1791_in5 <= VN_sign_in(10751) & VN_data_in(10751);
  VN1792_in0 <= VN_sign_in(10752) & VN_data_in(10752);
  VN1792_in1 <= VN_sign_in(10753) & VN_data_in(10753);
  VN1792_in2 <= VN_sign_in(10754) & VN_data_in(10754);
  VN1792_in3 <= VN_sign_in(10755) & VN_data_in(10755);
  VN1792_in4 <= VN_sign_in(10756) & VN_data_in(10756);
  VN1792_in5 <= VN_sign_in(10757) & VN_data_in(10757);
  VN1793_in0 <= VN_sign_in(10758) & VN_data_in(10758);
  VN1793_in1 <= VN_sign_in(10759) & VN_data_in(10759);
  VN1793_in2 <= VN_sign_in(10760) & VN_data_in(10760);
  VN1793_in3 <= VN_sign_in(10761) & VN_data_in(10761);
  VN1793_in4 <= VN_sign_in(10762) & VN_data_in(10762);
  VN1793_in5 <= VN_sign_in(10763) & VN_data_in(10763);
  VN1794_in0 <= VN_sign_in(10764) & VN_data_in(10764);
  VN1794_in1 <= VN_sign_in(10765) & VN_data_in(10765);
  VN1794_in2 <= VN_sign_in(10766) & VN_data_in(10766);
  VN1794_in3 <= VN_sign_in(10767) & VN_data_in(10767);
  VN1794_in4 <= VN_sign_in(10768) & VN_data_in(10768);
  VN1794_in5 <= VN_sign_in(10769) & VN_data_in(10769);
  VN1795_in0 <= VN_sign_in(10770) & VN_data_in(10770);
  VN1795_in1 <= VN_sign_in(10771) & VN_data_in(10771);
  VN1795_in2 <= VN_sign_in(10772) & VN_data_in(10772);
  VN1795_in3 <= VN_sign_in(10773) & VN_data_in(10773);
  VN1795_in4 <= VN_sign_in(10774) & VN_data_in(10774);
  VN1795_in5 <= VN_sign_in(10775) & VN_data_in(10775);
  VN1796_in0 <= VN_sign_in(10776) & VN_data_in(10776);
  VN1796_in1 <= VN_sign_in(10777) & VN_data_in(10777);
  VN1796_in2 <= VN_sign_in(10778) & VN_data_in(10778);
  VN1796_in3 <= VN_sign_in(10779) & VN_data_in(10779);
  VN1796_in4 <= VN_sign_in(10780) & VN_data_in(10780);
  VN1796_in5 <= VN_sign_in(10781) & VN_data_in(10781);
  VN1797_in0 <= VN_sign_in(10782) & VN_data_in(10782);
  VN1797_in1 <= VN_sign_in(10783) & VN_data_in(10783);
  VN1797_in2 <= VN_sign_in(10784) & VN_data_in(10784);
  VN1797_in3 <= VN_sign_in(10785) & VN_data_in(10785);
  VN1797_in4 <= VN_sign_in(10786) & VN_data_in(10786);
  VN1797_in5 <= VN_sign_in(10787) & VN_data_in(10787);
  VN1798_in0 <= VN_sign_in(10788) & VN_data_in(10788);
  VN1798_in1 <= VN_sign_in(10789) & VN_data_in(10789);
  VN1798_in2 <= VN_sign_in(10790) & VN_data_in(10790);
  VN1798_in3 <= VN_sign_in(10791) & VN_data_in(10791);
  VN1798_in4 <= VN_sign_in(10792) & VN_data_in(10792);
  VN1798_in5 <= VN_sign_in(10793) & VN_data_in(10793);
  VN1799_in0 <= VN_sign_in(10794) & VN_data_in(10794);
  VN1799_in1 <= VN_sign_in(10795) & VN_data_in(10795);
  VN1799_in2 <= VN_sign_in(10796) & VN_data_in(10796);
  VN1799_in3 <= VN_sign_in(10797) & VN_data_in(10797);
  VN1799_in4 <= VN_sign_in(10798) & VN_data_in(10798);
  VN1799_in5 <= VN_sign_in(10799) & VN_data_in(10799);
  VN1800_in0 <= VN_sign_in(10800) & VN_data_in(10800);
  VN1800_in1 <= VN_sign_in(10801) & VN_data_in(10801);
  VN1800_in2 <= VN_sign_in(10802) & VN_data_in(10802);
  VN1800_in3 <= VN_sign_in(10803) & VN_data_in(10803);
  VN1800_in4 <= VN_sign_in(10804) & VN_data_in(10804);
  VN1800_in5 <= VN_sign_in(10805) & VN_data_in(10805);
  VN1801_in0 <= VN_sign_in(10806) & VN_data_in(10806);
  VN1801_in1 <= VN_sign_in(10807) & VN_data_in(10807);
  VN1801_in2 <= VN_sign_in(10808) & VN_data_in(10808);
  VN1801_in3 <= VN_sign_in(10809) & VN_data_in(10809);
  VN1801_in4 <= VN_sign_in(10810) & VN_data_in(10810);
  VN1801_in5 <= VN_sign_in(10811) & VN_data_in(10811);
  VN1802_in0 <= VN_sign_in(10812) & VN_data_in(10812);
  VN1802_in1 <= VN_sign_in(10813) & VN_data_in(10813);
  VN1802_in2 <= VN_sign_in(10814) & VN_data_in(10814);
  VN1802_in3 <= VN_sign_in(10815) & VN_data_in(10815);
  VN1802_in4 <= VN_sign_in(10816) & VN_data_in(10816);
  VN1802_in5 <= VN_sign_in(10817) & VN_data_in(10817);
  VN1803_in0 <= VN_sign_in(10818) & VN_data_in(10818);
  VN1803_in1 <= VN_sign_in(10819) & VN_data_in(10819);
  VN1803_in2 <= VN_sign_in(10820) & VN_data_in(10820);
  VN1803_in3 <= VN_sign_in(10821) & VN_data_in(10821);
  VN1803_in4 <= VN_sign_in(10822) & VN_data_in(10822);
  VN1803_in5 <= VN_sign_in(10823) & VN_data_in(10823);
  VN1804_in0 <= VN_sign_in(10824) & VN_data_in(10824);
  VN1804_in1 <= VN_sign_in(10825) & VN_data_in(10825);
  VN1804_in2 <= VN_sign_in(10826) & VN_data_in(10826);
  VN1804_in3 <= VN_sign_in(10827) & VN_data_in(10827);
  VN1804_in4 <= VN_sign_in(10828) & VN_data_in(10828);
  VN1804_in5 <= VN_sign_in(10829) & VN_data_in(10829);
  VN1805_in0 <= VN_sign_in(10830) & VN_data_in(10830);
  VN1805_in1 <= VN_sign_in(10831) & VN_data_in(10831);
  VN1805_in2 <= VN_sign_in(10832) & VN_data_in(10832);
  VN1805_in3 <= VN_sign_in(10833) & VN_data_in(10833);
  VN1805_in4 <= VN_sign_in(10834) & VN_data_in(10834);
  VN1805_in5 <= VN_sign_in(10835) & VN_data_in(10835);
  VN1806_in0 <= VN_sign_in(10836) & VN_data_in(10836);
  VN1806_in1 <= VN_sign_in(10837) & VN_data_in(10837);
  VN1806_in2 <= VN_sign_in(10838) & VN_data_in(10838);
  VN1806_in3 <= VN_sign_in(10839) & VN_data_in(10839);
  VN1806_in4 <= VN_sign_in(10840) & VN_data_in(10840);
  VN1806_in5 <= VN_sign_in(10841) & VN_data_in(10841);
  VN1807_in0 <= VN_sign_in(10842) & VN_data_in(10842);
  VN1807_in1 <= VN_sign_in(10843) & VN_data_in(10843);
  VN1807_in2 <= VN_sign_in(10844) & VN_data_in(10844);
  VN1807_in3 <= VN_sign_in(10845) & VN_data_in(10845);
  VN1807_in4 <= VN_sign_in(10846) & VN_data_in(10846);
  VN1807_in5 <= VN_sign_in(10847) & VN_data_in(10847);
  VN1808_in0 <= VN_sign_in(10848) & VN_data_in(10848);
  VN1808_in1 <= VN_sign_in(10849) & VN_data_in(10849);
  VN1808_in2 <= VN_sign_in(10850) & VN_data_in(10850);
  VN1808_in3 <= VN_sign_in(10851) & VN_data_in(10851);
  VN1808_in4 <= VN_sign_in(10852) & VN_data_in(10852);
  VN1808_in5 <= VN_sign_in(10853) & VN_data_in(10853);
  VN1809_in0 <= VN_sign_in(10854) & VN_data_in(10854);
  VN1809_in1 <= VN_sign_in(10855) & VN_data_in(10855);
  VN1809_in2 <= VN_sign_in(10856) & VN_data_in(10856);
  VN1809_in3 <= VN_sign_in(10857) & VN_data_in(10857);
  VN1809_in4 <= VN_sign_in(10858) & VN_data_in(10858);
  VN1809_in5 <= VN_sign_in(10859) & VN_data_in(10859);
  VN1810_in0 <= VN_sign_in(10860) & VN_data_in(10860);
  VN1810_in1 <= VN_sign_in(10861) & VN_data_in(10861);
  VN1810_in2 <= VN_sign_in(10862) & VN_data_in(10862);
  VN1810_in3 <= VN_sign_in(10863) & VN_data_in(10863);
  VN1810_in4 <= VN_sign_in(10864) & VN_data_in(10864);
  VN1810_in5 <= VN_sign_in(10865) & VN_data_in(10865);
  VN1811_in0 <= VN_sign_in(10866) & VN_data_in(10866);
  VN1811_in1 <= VN_sign_in(10867) & VN_data_in(10867);
  VN1811_in2 <= VN_sign_in(10868) & VN_data_in(10868);
  VN1811_in3 <= VN_sign_in(10869) & VN_data_in(10869);
  VN1811_in4 <= VN_sign_in(10870) & VN_data_in(10870);
  VN1811_in5 <= VN_sign_in(10871) & VN_data_in(10871);
  VN1812_in0 <= VN_sign_in(10872) & VN_data_in(10872);
  VN1812_in1 <= VN_sign_in(10873) & VN_data_in(10873);
  VN1812_in2 <= VN_sign_in(10874) & VN_data_in(10874);
  VN1812_in3 <= VN_sign_in(10875) & VN_data_in(10875);
  VN1812_in4 <= VN_sign_in(10876) & VN_data_in(10876);
  VN1812_in5 <= VN_sign_in(10877) & VN_data_in(10877);
  VN1813_in0 <= VN_sign_in(10878) & VN_data_in(10878);
  VN1813_in1 <= VN_sign_in(10879) & VN_data_in(10879);
  VN1813_in2 <= VN_sign_in(10880) & VN_data_in(10880);
  VN1813_in3 <= VN_sign_in(10881) & VN_data_in(10881);
  VN1813_in4 <= VN_sign_in(10882) & VN_data_in(10882);
  VN1813_in5 <= VN_sign_in(10883) & VN_data_in(10883);
  VN1814_in0 <= VN_sign_in(10884) & VN_data_in(10884);
  VN1814_in1 <= VN_sign_in(10885) & VN_data_in(10885);
  VN1814_in2 <= VN_sign_in(10886) & VN_data_in(10886);
  VN1814_in3 <= VN_sign_in(10887) & VN_data_in(10887);
  VN1814_in4 <= VN_sign_in(10888) & VN_data_in(10888);
  VN1814_in5 <= VN_sign_in(10889) & VN_data_in(10889);
  VN1815_in0 <= VN_sign_in(10890) & VN_data_in(10890);
  VN1815_in1 <= VN_sign_in(10891) & VN_data_in(10891);
  VN1815_in2 <= VN_sign_in(10892) & VN_data_in(10892);
  VN1815_in3 <= VN_sign_in(10893) & VN_data_in(10893);
  VN1815_in4 <= VN_sign_in(10894) & VN_data_in(10894);
  VN1815_in5 <= VN_sign_in(10895) & VN_data_in(10895);
  VN1816_in0 <= VN_sign_in(10896) & VN_data_in(10896);
  VN1816_in1 <= VN_sign_in(10897) & VN_data_in(10897);
  VN1816_in2 <= VN_sign_in(10898) & VN_data_in(10898);
  VN1816_in3 <= VN_sign_in(10899) & VN_data_in(10899);
  VN1816_in4 <= VN_sign_in(10900) & VN_data_in(10900);
  VN1816_in5 <= VN_sign_in(10901) & VN_data_in(10901);
  VN1817_in0 <= VN_sign_in(10902) & VN_data_in(10902);
  VN1817_in1 <= VN_sign_in(10903) & VN_data_in(10903);
  VN1817_in2 <= VN_sign_in(10904) & VN_data_in(10904);
  VN1817_in3 <= VN_sign_in(10905) & VN_data_in(10905);
  VN1817_in4 <= VN_sign_in(10906) & VN_data_in(10906);
  VN1817_in5 <= VN_sign_in(10907) & VN_data_in(10907);
  VN1818_in0 <= VN_sign_in(10908) & VN_data_in(10908);
  VN1818_in1 <= VN_sign_in(10909) & VN_data_in(10909);
  VN1818_in2 <= VN_sign_in(10910) & VN_data_in(10910);
  VN1818_in3 <= VN_sign_in(10911) & VN_data_in(10911);
  VN1818_in4 <= VN_sign_in(10912) & VN_data_in(10912);
  VN1818_in5 <= VN_sign_in(10913) & VN_data_in(10913);
  VN1819_in0 <= VN_sign_in(10914) & VN_data_in(10914);
  VN1819_in1 <= VN_sign_in(10915) & VN_data_in(10915);
  VN1819_in2 <= VN_sign_in(10916) & VN_data_in(10916);
  VN1819_in3 <= VN_sign_in(10917) & VN_data_in(10917);
  VN1819_in4 <= VN_sign_in(10918) & VN_data_in(10918);
  VN1819_in5 <= VN_sign_in(10919) & VN_data_in(10919);
  VN1820_in0 <= VN_sign_in(10920) & VN_data_in(10920);
  VN1820_in1 <= VN_sign_in(10921) & VN_data_in(10921);
  VN1820_in2 <= VN_sign_in(10922) & VN_data_in(10922);
  VN1820_in3 <= VN_sign_in(10923) & VN_data_in(10923);
  VN1820_in4 <= VN_sign_in(10924) & VN_data_in(10924);
  VN1820_in5 <= VN_sign_in(10925) & VN_data_in(10925);
  VN1821_in0 <= VN_sign_in(10926) & VN_data_in(10926);
  VN1821_in1 <= VN_sign_in(10927) & VN_data_in(10927);
  VN1821_in2 <= VN_sign_in(10928) & VN_data_in(10928);
  VN1821_in3 <= VN_sign_in(10929) & VN_data_in(10929);
  VN1821_in4 <= VN_sign_in(10930) & VN_data_in(10930);
  VN1821_in5 <= VN_sign_in(10931) & VN_data_in(10931);
  VN1822_in0 <= VN_sign_in(10932) & VN_data_in(10932);
  VN1822_in1 <= VN_sign_in(10933) & VN_data_in(10933);
  VN1822_in2 <= VN_sign_in(10934) & VN_data_in(10934);
  VN1822_in3 <= VN_sign_in(10935) & VN_data_in(10935);
  VN1822_in4 <= VN_sign_in(10936) & VN_data_in(10936);
  VN1822_in5 <= VN_sign_in(10937) & VN_data_in(10937);
  VN1823_in0 <= VN_sign_in(10938) & VN_data_in(10938);
  VN1823_in1 <= VN_sign_in(10939) & VN_data_in(10939);
  VN1823_in2 <= VN_sign_in(10940) & VN_data_in(10940);
  VN1823_in3 <= VN_sign_in(10941) & VN_data_in(10941);
  VN1823_in4 <= VN_sign_in(10942) & VN_data_in(10942);
  VN1823_in5 <= VN_sign_in(10943) & VN_data_in(10943);
  VN1824_in0 <= VN_sign_in(10944) & VN_data_in(10944);
  VN1824_in1 <= VN_sign_in(10945) & VN_data_in(10945);
  VN1824_in2 <= VN_sign_in(10946) & VN_data_in(10946);
  VN1824_in3 <= VN_sign_in(10947) & VN_data_in(10947);
  VN1824_in4 <= VN_sign_in(10948) & VN_data_in(10948);
  VN1824_in5 <= VN_sign_in(10949) & VN_data_in(10949);
  VN1825_in0 <= VN_sign_in(10950) & VN_data_in(10950);
  VN1825_in1 <= VN_sign_in(10951) & VN_data_in(10951);
  VN1825_in2 <= VN_sign_in(10952) & VN_data_in(10952);
  VN1825_in3 <= VN_sign_in(10953) & VN_data_in(10953);
  VN1825_in4 <= VN_sign_in(10954) & VN_data_in(10954);
  VN1825_in5 <= VN_sign_in(10955) & VN_data_in(10955);
  VN1826_in0 <= VN_sign_in(10956) & VN_data_in(10956);
  VN1826_in1 <= VN_sign_in(10957) & VN_data_in(10957);
  VN1826_in2 <= VN_sign_in(10958) & VN_data_in(10958);
  VN1826_in3 <= VN_sign_in(10959) & VN_data_in(10959);
  VN1826_in4 <= VN_sign_in(10960) & VN_data_in(10960);
  VN1826_in5 <= VN_sign_in(10961) & VN_data_in(10961);
  VN1827_in0 <= VN_sign_in(10962) & VN_data_in(10962);
  VN1827_in1 <= VN_sign_in(10963) & VN_data_in(10963);
  VN1827_in2 <= VN_sign_in(10964) & VN_data_in(10964);
  VN1827_in3 <= VN_sign_in(10965) & VN_data_in(10965);
  VN1827_in4 <= VN_sign_in(10966) & VN_data_in(10966);
  VN1827_in5 <= VN_sign_in(10967) & VN_data_in(10967);
  VN1828_in0 <= VN_sign_in(10968) & VN_data_in(10968);
  VN1828_in1 <= VN_sign_in(10969) & VN_data_in(10969);
  VN1828_in2 <= VN_sign_in(10970) & VN_data_in(10970);
  VN1828_in3 <= VN_sign_in(10971) & VN_data_in(10971);
  VN1828_in4 <= VN_sign_in(10972) & VN_data_in(10972);
  VN1828_in5 <= VN_sign_in(10973) & VN_data_in(10973);
  VN1829_in0 <= VN_sign_in(10974) & VN_data_in(10974);
  VN1829_in1 <= VN_sign_in(10975) & VN_data_in(10975);
  VN1829_in2 <= VN_sign_in(10976) & VN_data_in(10976);
  VN1829_in3 <= VN_sign_in(10977) & VN_data_in(10977);
  VN1829_in4 <= VN_sign_in(10978) & VN_data_in(10978);
  VN1829_in5 <= VN_sign_in(10979) & VN_data_in(10979);
  VN1830_in0 <= VN_sign_in(10980) & VN_data_in(10980);
  VN1830_in1 <= VN_sign_in(10981) & VN_data_in(10981);
  VN1830_in2 <= VN_sign_in(10982) & VN_data_in(10982);
  VN1830_in3 <= VN_sign_in(10983) & VN_data_in(10983);
  VN1830_in4 <= VN_sign_in(10984) & VN_data_in(10984);
  VN1830_in5 <= VN_sign_in(10985) & VN_data_in(10985);
  VN1831_in0 <= VN_sign_in(10986) & VN_data_in(10986);
  VN1831_in1 <= VN_sign_in(10987) & VN_data_in(10987);
  VN1831_in2 <= VN_sign_in(10988) & VN_data_in(10988);
  VN1831_in3 <= VN_sign_in(10989) & VN_data_in(10989);
  VN1831_in4 <= VN_sign_in(10990) & VN_data_in(10990);
  VN1831_in5 <= VN_sign_in(10991) & VN_data_in(10991);
  VN1832_in0 <= VN_sign_in(10992) & VN_data_in(10992);
  VN1832_in1 <= VN_sign_in(10993) & VN_data_in(10993);
  VN1832_in2 <= VN_sign_in(10994) & VN_data_in(10994);
  VN1832_in3 <= VN_sign_in(10995) & VN_data_in(10995);
  VN1832_in4 <= VN_sign_in(10996) & VN_data_in(10996);
  VN1832_in5 <= VN_sign_in(10997) & VN_data_in(10997);
  VN1833_in0 <= VN_sign_in(10998) & VN_data_in(10998);
  VN1833_in1 <= VN_sign_in(10999) & VN_data_in(10999);
  VN1833_in2 <= VN_sign_in(11000) & VN_data_in(11000);
  VN1833_in3 <= VN_sign_in(11001) & VN_data_in(11001);
  VN1833_in4 <= VN_sign_in(11002) & VN_data_in(11002);
  VN1833_in5 <= VN_sign_in(11003) & VN_data_in(11003);
  VN1834_in0 <= VN_sign_in(11004) & VN_data_in(11004);
  VN1834_in1 <= VN_sign_in(11005) & VN_data_in(11005);
  VN1834_in2 <= VN_sign_in(11006) & VN_data_in(11006);
  VN1834_in3 <= VN_sign_in(11007) & VN_data_in(11007);
  VN1834_in4 <= VN_sign_in(11008) & VN_data_in(11008);
  VN1834_in5 <= VN_sign_in(11009) & VN_data_in(11009);
  VN1835_in0 <= VN_sign_in(11010) & VN_data_in(11010);
  VN1835_in1 <= VN_sign_in(11011) & VN_data_in(11011);
  VN1835_in2 <= VN_sign_in(11012) & VN_data_in(11012);
  VN1835_in3 <= VN_sign_in(11013) & VN_data_in(11013);
  VN1835_in4 <= VN_sign_in(11014) & VN_data_in(11014);
  VN1835_in5 <= VN_sign_in(11015) & VN_data_in(11015);
  VN1836_in0 <= VN_sign_in(11016) & VN_data_in(11016);
  VN1836_in1 <= VN_sign_in(11017) & VN_data_in(11017);
  VN1836_in2 <= VN_sign_in(11018) & VN_data_in(11018);
  VN1836_in3 <= VN_sign_in(11019) & VN_data_in(11019);
  VN1836_in4 <= VN_sign_in(11020) & VN_data_in(11020);
  VN1836_in5 <= VN_sign_in(11021) & VN_data_in(11021);
  VN1837_in0 <= VN_sign_in(11022) & VN_data_in(11022);
  VN1837_in1 <= VN_sign_in(11023) & VN_data_in(11023);
  VN1837_in2 <= VN_sign_in(11024) & VN_data_in(11024);
  VN1837_in3 <= VN_sign_in(11025) & VN_data_in(11025);
  VN1837_in4 <= VN_sign_in(11026) & VN_data_in(11026);
  VN1837_in5 <= VN_sign_in(11027) & VN_data_in(11027);
  VN1838_in0 <= VN_sign_in(11028) & VN_data_in(11028);
  VN1838_in1 <= VN_sign_in(11029) & VN_data_in(11029);
  VN1838_in2 <= VN_sign_in(11030) & VN_data_in(11030);
  VN1838_in3 <= VN_sign_in(11031) & VN_data_in(11031);
  VN1838_in4 <= VN_sign_in(11032) & VN_data_in(11032);
  VN1838_in5 <= VN_sign_in(11033) & VN_data_in(11033);
  VN1839_in0 <= VN_sign_in(11034) & VN_data_in(11034);
  VN1839_in1 <= VN_sign_in(11035) & VN_data_in(11035);
  VN1839_in2 <= VN_sign_in(11036) & VN_data_in(11036);
  VN1839_in3 <= VN_sign_in(11037) & VN_data_in(11037);
  VN1839_in4 <= VN_sign_in(11038) & VN_data_in(11038);
  VN1839_in5 <= VN_sign_in(11039) & VN_data_in(11039);
  VN1840_in0 <= VN_sign_in(11040) & VN_data_in(11040);
  VN1840_in1 <= VN_sign_in(11041) & VN_data_in(11041);
  VN1840_in2 <= VN_sign_in(11042) & VN_data_in(11042);
  VN1840_in3 <= VN_sign_in(11043) & VN_data_in(11043);
  VN1840_in4 <= VN_sign_in(11044) & VN_data_in(11044);
  VN1840_in5 <= VN_sign_in(11045) & VN_data_in(11045);
  VN1841_in0 <= VN_sign_in(11046) & VN_data_in(11046);
  VN1841_in1 <= VN_sign_in(11047) & VN_data_in(11047);
  VN1841_in2 <= VN_sign_in(11048) & VN_data_in(11048);
  VN1841_in3 <= VN_sign_in(11049) & VN_data_in(11049);
  VN1841_in4 <= VN_sign_in(11050) & VN_data_in(11050);
  VN1841_in5 <= VN_sign_in(11051) & VN_data_in(11051);
  VN1842_in0 <= VN_sign_in(11052) & VN_data_in(11052);
  VN1842_in1 <= VN_sign_in(11053) & VN_data_in(11053);
  VN1842_in2 <= VN_sign_in(11054) & VN_data_in(11054);
  VN1842_in3 <= VN_sign_in(11055) & VN_data_in(11055);
  VN1842_in4 <= VN_sign_in(11056) & VN_data_in(11056);
  VN1842_in5 <= VN_sign_in(11057) & VN_data_in(11057);
  VN1843_in0 <= VN_sign_in(11058) & VN_data_in(11058);
  VN1843_in1 <= VN_sign_in(11059) & VN_data_in(11059);
  VN1843_in2 <= VN_sign_in(11060) & VN_data_in(11060);
  VN1843_in3 <= VN_sign_in(11061) & VN_data_in(11061);
  VN1843_in4 <= VN_sign_in(11062) & VN_data_in(11062);
  VN1843_in5 <= VN_sign_in(11063) & VN_data_in(11063);
  VN1844_in0 <= VN_sign_in(11064) & VN_data_in(11064);
  VN1844_in1 <= VN_sign_in(11065) & VN_data_in(11065);
  VN1844_in2 <= VN_sign_in(11066) & VN_data_in(11066);
  VN1844_in3 <= VN_sign_in(11067) & VN_data_in(11067);
  VN1844_in4 <= VN_sign_in(11068) & VN_data_in(11068);
  VN1844_in5 <= VN_sign_in(11069) & VN_data_in(11069);
  VN1845_in0 <= VN_sign_in(11070) & VN_data_in(11070);
  VN1845_in1 <= VN_sign_in(11071) & VN_data_in(11071);
  VN1845_in2 <= VN_sign_in(11072) & VN_data_in(11072);
  VN1845_in3 <= VN_sign_in(11073) & VN_data_in(11073);
  VN1845_in4 <= VN_sign_in(11074) & VN_data_in(11074);
  VN1845_in5 <= VN_sign_in(11075) & VN_data_in(11075);
  VN1846_in0 <= VN_sign_in(11076) & VN_data_in(11076);
  VN1846_in1 <= VN_sign_in(11077) & VN_data_in(11077);
  VN1846_in2 <= VN_sign_in(11078) & VN_data_in(11078);
  VN1846_in3 <= VN_sign_in(11079) & VN_data_in(11079);
  VN1846_in4 <= VN_sign_in(11080) & VN_data_in(11080);
  VN1846_in5 <= VN_sign_in(11081) & VN_data_in(11081);
  VN1847_in0 <= VN_sign_in(11082) & VN_data_in(11082);
  VN1847_in1 <= VN_sign_in(11083) & VN_data_in(11083);
  VN1847_in2 <= VN_sign_in(11084) & VN_data_in(11084);
  VN1847_in3 <= VN_sign_in(11085) & VN_data_in(11085);
  VN1847_in4 <= VN_sign_in(11086) & VN_data_in(11086);
  VN1847_in5 <= VN_sign_in(11087) & VN_data_in(11087);
  VN1848_in0 <= VN_sign_in(11088) & VN_data_in(11088);
  VN1848_in1 <= VN_sign_in(11089) & VN_data_in(11089);
  VN1848_in2 <= VN_sign_in(11090) & VN_data_in(11090);
  VN1848_in3 <= VN_sign_in(11091) & VN_data_in(11091);
  VN1848_in4 <= VN_sign_in(11092) & VN_data_in(11092);
  VN1848_in5 <= VN_sign_in(11093) & VN_data_in(11093);
  VN1849_in0 <= VN_sign_in(11094) & VN_data_in(11094);
  VN1849_in1 <= VN_sign_in(11095) & VN_data_in(11095);
  VN1849_in2 <= VN_sign_in(11096) & VN_data_in(11096);
  VN1849_in3 <= VN_sign_in(11097) & VN_data_in(11097);
  VN1849_in4 <= VN_sign_in(11098) & VN_data_in(11098);
  VN1849_in5 <= VN_sign_in(11099) & VN_data_in(11099);
  VN1850_in0 <= VN_sign_in(11100) & VN_data_in(11100);
  VN1850_in1 <= VN_sign_in(11101) & VN_data_in(11101);
  VN1850_in2 <= VN_sign_in(11102) & VN_data_in(11102);
  VN1850_in3 <= VN_sign_in(11103) & VN_data_in(11103);
  VN1850_in4 <= VN_sign_in(11104) & VN_data_in(11104);
  VN1850_in5 <= VN_sign_in(11105) & VN_data_in(11105);
  VN1851_in0 <= VN_sign_in(11106) & VN_data_in(11106);
  VN1851_in1 <= VN_sign_in(11107) & VN_data_in(11107);
  VN1851_in2 <= VN_sign_in(11108) & VN_data_in(11108);
  VN1851_in3 <= VN_sign_in(11109) & VN_data_in(11109);
  VN1851_in4 <= VN_sign_in(11110) & VN_data_in(11110);
  VN1851_in5 <= VN_sign_in(11111) & VN_data_in(11111);
  VN1852_in0 <= VN_sign_in(11112) & VN_data_in(11112);
  VN1852_in1 <= VN_sign_in(11113) & VN_data_in(11113);
  VN1852_in2 <= VN_sign_in(11114) & VN_data_in(11114);
  VN1852_in3 <= VN_sign_in(11115) & VN_data_in(11115);
  VN1852_in4 <= VN_sign_in(11116) & VN_data_in(11116);
  VN1852_in5 <= VN_sign_in(11117) & VN_data_in(11117);
  VN1853_in0 <= VN_sign_in(11118) & VN_data_in(11118);
  VN1853_in1 <= VN_sign_in(11119) & VN_data_in(11119);
  VN1853_in2 <= VN_sign_in(11120) & VN_data_in(11120);
  VN1853_in3 <= VN_sign_in(11121) & VN_data_in(11121);
  VN1853_in4 <= VN_sign_in(11122) & VN_data_in(11122);
  VN1853_in5 <= VN_sign_in(11123) & VN_data_in(11123);
  VN1854_in0 <= VN_sign_in(11124) & VN_data_in(11124);
  VN1854_in1 <= VN_sign_in(11125) & VN_data_in(11125);
  VN1854_in2 <= VN_sign_in(11126) & VN_data_in(11126);
  VN1854_in3 <= VN_sign_in(11127) & VN_data_in(11127);
  VN1854_in4 <= VN_sign_in(11128) & VN_data_in(11128);
  VN1854_in5 <= VN_sign_in(11129) & VN_data_in(11129);
  VN1855_in0 <= VN_sign_in(11130) & VN_data_in(11130);
  VN1855_in1 <= VN_sign_in(11131) & VN_data_in(11131);
  VN1855_in2 <= VN_sign_in(11132) & VN_data_in(11132);
  VN1855_in3 <= VN_sign_in(11133) & VN_data_in(11133);
  VN1855_in4 <= VN_sign_in(11134) & VN_data_in(11134);
  VN1855_in5 <= VN_sign_in(11135) & VN_data_in(11135);
  VN1856_in0 <= VN_sign_in(11136) & VN_data_in(11136);
  VN1856_in1 <= VN_sign_in(11137) & VN_data_in(11137);
  VN1856_in2 <= VN_sign_in(11138) & VN_data_in(11138);
  VN1856_in3 <= VN_sign_in(11139) & VN_data_in(11139);
  VN1856_in4 <= VN_sign_in(11140) & VN_data_in(11140);
  VN1856_in5 <= VN_sign_in(11141) & VN_data_in(11141);
  VN1857_in0 <= VN_sign_in(11142) & VN_data_in(11142);
  VN1857_in1 <= VN_sign_in(11143) & VN_data_in(11143);
  VN1857_in2 <= VN_sign_in(11144) & VN_data_in(11144);
  VN1857_in3 <= VN_sign_in(11145) & VN_data_in(11145);
  VN1857_in4 <= VN_sign_in(11146) & VN_data_in(11146);
  VN1857_in5 <= VN_sign_in(11147) & VN_data_in(11147);
  VN1858_in0 <= VN_sign_in(11148) & VN_data_in(11148);
  VN1858_in1 <= VN_sign_in(11149) & VN_data_in(11149);
  VN1858_in2 <= VN_sign_in(11150) & VN_data_in(11150);
  VN1858_in3 <= VN_sign_in(11151) & VN_data_in(11151);
  VN1858_in4 <= VN_sign_in(11152) & VN_data_in(11152);
  VN1858_in5 <= VN_sign_in(11153) & VN_data_in(11153);
  VN1859_in0 <= VN_sign_in(11154) & VN_data_in(11154);
  VN1859_in1 <= VN_sign_in(11155) & VN_data_in(11155);
  VN1859_in2 <= VN_sign_in(11156) & VN_data_in(11156);
  VN1859_in3 <= VN_sign_in(11157) & VN_data_in(11157);
  VN1859_in4 <= VN_sign_in(11158) & VN_data_in(11158);
  VN1859_in5 <= VN_sign_in(11159) & VN_data_in(11159);
  VN1860_in0 <= VN_sign_in(11160) & VN_data_in(11160);
  VN1860_in1 <= VN_sign_in(11161) & VN_data_in(11161);
  VN1860_in2 <= VN_sign_in(11162) & VN_data_in(11162);
  VN1860_in3 <= VN_sign_in(11163) & VN_data_in(11163);
  VN1860_in4 <= VN_sign_in(11164) & VN_data_in(11164);
  VN1860_in5 <= VN_sign_in(11165) & VN_data_in(11165);
  VN1861_in0 <= VN_sign_in(11166) & VN_data_in(11166);
  VN1861_in1 <= VN_sign_in(11167) & VN_data_in(11167);
  VN1861_in2 <= VN_sign_in(11168) & VN_data_in(11168);
  VN1861_in3 <= VN_sign_in(11169) & VN_data_in(11169);
  VN1861_in4 <= VN_sign_in(11170) & VN_data_in(11170);
  VN1861_in5 <= VN_sign_in(11171) & VN_data_in(11171);
  VN1862_in0 <= VN_sign_in(11172) & VN_data_in(11172);
  VN1862_in1 <= VN_sign_in(11173) & VN_data_in(11173);
  VN1862_in2 <= VN_sign_in(11174) & VN_data_in(11174);
  VN1862_in3 <= VN_sign_in(11175) & VN_data_in(11175);
  VN1862_in4 <= VN_sign_in(11176) & VN_data_in(11176);
  VN1862_in5 <= VN_sign_in(11177) & VN_data_in(11177);
  VN1863_in0 <= VN_sign_in(11178) & VN_data_in(11178);
  VN1863_in1 <= VN_sign_in(11179) & VN_data_in(11179);
  VN1863_in2 <= VN_sign_in(11180) & VN_data_in(11180);
  VN1863_in3 <= VN_sign_in(11181) & VN_data_in(11181);
  VN1863_in4 <= VN_sign_in(11182) & VN_data_in(11182);
  VN1863_in5 <= VN_sign_in(11183) & VN_data_in(11183);
  VN1864_in0 <= VN_sign_in(11184) & VN_data_in(11184);
  VN1864_in1 <= VN_sign_in(11185) & VN_data_in(11185);
  VN1864_in2 <= VN_sign_in(11186) & VN_data_in(11186);
  VN1864_in3 <= VN_sign_in(11187) & VN_data_in(11187);
  VN1864_in4 <= VN_sign_in(11188) & VN_data_in(11188);
  VN1864_in5 <= VN_sign_in(11189) & VN_data_in(11189);
  VN1865_in0 <= VN_sign_in(11190) & VN_data_in(11190);
  VN1865_in1 <= VN_sign_in(11191) & VN_data_in(11191);
  VN1865_in2 <= VN_sign_in(11192) & VN_data_in(11192);
  VN1865_in3 <= VN_sign_in(11193) & VN_data_in(11193);
  VN1865_in4 <= VN_sign_in(11194) & VN_data_in(11194);
  VN1865_in5 <= VN_sign_in(11195) & VN_data_in(11195);
  VN1866_in0 <= VN_sign_in(11196) & VN_data_in(11196);
  VN1866_in1 <= VN_sign_in(11197) & VN_data_in(11197);
  VN1866_in2 <= VN_sign_in(11198) & VN_data_in(11198);
  VN1866_in3 <= VN_sign_in(11199) & VN_data_in(11199);
  VN1866_in4 <= VN_sign_in(11200) & VN_data_in(11200);
  VN1866_in5 <= VN_sign_in(11201) & VN_data_in(11201);
  VN1867_in0 <= VN_sign_in(11202) & VN_data_in(11202);
  VN1867_in1 <= VN_sign_in(11203) & VN_data_in(11203);
  VN1867_in2 <= VN_sign_in(11204) & VN_data_in(11204);
  VN1867_in3 <= VN_sign_in(11205) & VN_data_in(11205);
  VN1867_in4 <= VN_sign_in(11206) & VN_data_in(11206);
  VN1867_in5 <= VN_sign_in(11207) & VN_data_in(11207);
  VN1868_in0 <= VN_sign_in(11208) & VN_data_in(11208);
  VN1868_in1 <= VN_sign_in(11209) & VN_data_in(11209);
  VN1868_in2 <= VN_sign_in(11210) & VN_data_in(11210);
  VN1868_in3 <= VN_sign_in(11211) & VN_data_in(11211);
  VN1868_in4 <= VN_sign_in(11212) & VN_data_in(11212);
  VN1868_in5 <= VN_sign_in(11213) & VN_data_in(11213);
  VN1869_in0 <= VN_sign_in(11214) & VN_data_in(11214);
  VN1869_in1 <= VN_sign_in(11215) & VN_data_in(11215);
  VN1869_in2 <= VN_sign_in(11216) & VN_data_in(11216);
  VN1869_in3 <= VN_sign_in(11217) & VN_data_in(11217);
  VN1869_in4 <= VN_sign_in(11218) & VN_data_in(11218);
  VN1869_in5 <= VN_sign_in(11219) & VN_data_in(11219);
  VN1870_in0 <= VN_sign_in(11220) & VN_data_in(11220);
  VN1870_in1 <= VN_sign_in(11221) & VN_data_in(11221);
  VN1870_in2 <= VN_sign_in(11222) & VN_data_in(11222);
  VN1870_in3 <= VN_sign_in(11223) & VN_data_in(11223);
  VN1870_in4 <= VN_sign_in(11224) & VN_data_in(11224);
  VN1870_in5 <= VN_sign_in(11225) & VN_data_in(11225);
  VN1871_in0 <= VN_sign_in(11226) & VN_data_in(11226);
  VN1871_in1 <= VN_sign_in(11227) & VN_data_in(11227);
  VN1871_in2 <= VN_sign_in(11228) & VN_data_in(11228);
  VN1871_in3 <= VN_sign_in(11229) & VN_data_in(11229);
  VN1871_in4 <= VN_sign_in(11230) & VN_data_in(11230);
  VN1871_in5 <= VN_sign_in(11231) & VN_data_in(11231);
  VN1872_in0 <= VN_sign_in(11232) & VN_data_in(11232);
  VN1872_in1 <= VN_sign_in(11233) & VN_data_in(11233);
  VN1872_in2 <= VN_sign_in(11234) & VN_data_in(11234);
  VN1872_in3 <= VN_sign_in(11235) & VN_data_in(11235);
  VN1872_in4 <= VN_sign_in(11236) & VN_data_in(11236);
  VN1872_in5 <= VN_sign_in(11237) & VN_data_in(11237);
  VN1873_in0 <= VN_sign_in(11238) & VN_data_in(11238);
  VN1873_in1 <= VN_sign_in(11239) & VN_data_in(11239);
  VN1873_in2 <= VN_sign_in(11240) & VN_data_in(11240);
  VN1873_in3 <= VN_sign_in(11241) & VN_data_in(11241);
  VN1873_in4 <= VN_sign_in(11242) & VN_data_in(11242);
  VN1873_in5 <= VN_sign_in(11243) & VN_data_in(11243);
  VN1874_in0 <= VN_sign_in(11244) & VN_data_in(11244);
  VN1874_in1 <= VN_sign_in(11245) & VN_data_in(11245);
  VN1874_in2 <= VN_sign_in(11246) & VN_data_in(11246);
  VN1874_in3 <= VN_sign_in(11247) & VN_data_in(11247);
  VN1874_in4 <= VN_sign_in(11248) & VN_data_in(11248);
  VN1874_in5 <= VN_sign_in(11249) & VN_data_in(11249);
  VN1875_in0 <= VN_sign_in(11250) & VN_data_in(11250);
  VN1875_in1 <= VN_sign_in(11251) & VN_data_in(11251);
  VN1875_in2 <= VN_sign_in(11252) & VN_data_in(11252);
  VN1875_in3 <= VN_sign_in(11253) & VN_data_in(11253);
  VN1875_in4 <= VN_sign_in(11254) & VN_data_in(11254);
  VN1875_in5 <= VN_sign_in(11255) & VN_data_in(11255);
  VN1876_in0 <= VN_sign_in(11256) & VN_data_in(11256);
  VN1876_in1 <= VN_sign_in(11257) & VN_data_in(11257);
  VN1876_in2 <= VN_sign_in(11258) & VN_data_in(11258);
  VN1876_in3 <= VN_sign_in(11259) & VN_data_in(11259);
  VN1876_in4 <= VN_sign_in(11260) & VN_data_in(11260);
  VN1876_in5 <= VN_sign_in(11261) & VN_data_in(11261);
  VN1877_in0 <= VN_sign_in(11262) & VN_data_in(11262);
  VN1877_in1 <= VN_sign_in(11263) & VN_data_in(11263);
  VN1877_in2 <= VN_sign_in(11264) & VN_data_in(11264);
  VN1877_in3 <= VN_sign_in(11265) & VN_data_in(11265);
  VN1877_in4 <= VN_sign_in(11266) & VN_data_in(11266);
  VN1877_in5 <= VN_sign_in(11267) & VN_data_in(11267);
  VN1878_in0 <= VN_sign_in(11268) & VN_data_in(11268);
  VN1878_in1 <= VN_sign_in(11269) & VN_data_in(11269);
  VN1878_in2 <= VN_sign_in(11270) & VN_data_in(11270);
  VN1878_in3 <= VN_sign_in(11271) & VN_data_in(11271);
  VN1878_in4 <= VN_sign_in(11272) & VN_data_in(11272);
  VN1878_in5 <= VN_sign_in(11273) & VN_data_in(11273);
  VN1879_in0 <= VN_sign_in(11274) & VN_data_in(11274);
  VN1879_in1 <= VN_sign_in(11275) & VN_data_in(11275);
  VN1879_in2 <= VN_sign_in(11276) & VN_data_in(11276);
  VN1879_in3 <= VN_sign_in(11277) & VN_data_in(11277);
  VN1879_in4 <= VN_sign_in(11278) & VN_data_in(11278);
  VN1879_in5 <= VN_sign_in(11279) & VN_data_in(11279);
  VN1880_in0 <= VN_sign_in(11280) & VN_data_in(11280);
  VN1880_in1 <= VN_sign_in(11281) & VN_data_in(11281);
  VN1880_in2 <= VN_sign_in(11282) & VN_data_in(11282);
  VN1880_in3 <= VN_sign_in(11283) & VN_data_in(11283);
  VN1880_in4 <= VN_sign_in(11284) & VN_data_in(11284);
  VN1880_in5 <= VN_sign_in(11285) & VN_data_in(11285);
  VN1881_in0 <= VN_sign_in(11286) & VN_data_in(11286);
  VN1881_in1 <= VN_sign_in(11287) & VN_data_in(11287);
  VN1881_in2 <= VN_sign_in(11288) & VN_data_in(11288);
  VN1881_in3 <= VN_sign_in(11289) & VN_data_in(11289);
  VN1881_in4 <= VN_sign_in(11290) & VN_data_in(11290);
  VN1881_in5 <= VN_sign_in(11291) & VN_data_in(11291);
  VN1882_in0 <= VN_sign_in(11292) & VN_data_in(11292);
  VN1882_in1 <= VN_sign_in(11293) & VN_data_in(11293);
  VN1882_in2 <= VN_sign_in(11294) & VN_data_in(11294);
  VN1882_in3 <= VN_sign_in(11295) & VN_data_in(11295);
  VN1882_in4 <= VN_sign_in(11296) & VN_data_in(11296);
  VN1882_in5 <= VN_sign_in(11297) & VN_data_in(11297);
  VN1883_in0 <= VN_sign_in(11298) & VN_data_in(11298);
  VN1883_in1 <= VN_sign_in(11299) & VN_data_in(11299);
  VN1883_in2 <= VN_sign_in(11300) & VN_data_in(11300);
  VN1883_in3 <= VN_sign_in(11301) & VN_data_in(11301);
  VN1883_in4 <= VN_sign_in(11302) & VN_data_in(11302);
  VN1883_in5 <= VN_sign_in(11303) & VN_data_in(11303);
  VN1884_in0 <= VN_sign_in(11304) & VN_data_in(11304);
  VN1884_in1 <= VN_sign_in(11305) & VN_data_in(11305);
  VN1884_in2 <= VN_sign_in(11306) & VN_data_in(11306);
  VN1884_in3 <= VN_sign_in(11307) & VN_data_in(11307);
  VN1884_in4 <= VN_sign_in(11308) & VN_data_in(11308);
  VN1884_in5 <= VN_sign_in(11309) & VN_data_in(11309);
  VN1885_in0 <= VN_sign_in(11310) & VN_data_in(11310);
  VN1885_in1 <= VN_sign_in(11311) & VN_data_in(11311);
  VN1885_in2 <= VN_sign_in(11312) & VN_data_in(11312);
  VN1885_in3 <= VN_sign_in(11313) & VN_data_in(11313);
  VN1885_in4 <= VN_sign_in(11314) & VN_data_in(11314);
  VN1885_in5 <= VN_sign_in(11315) & VN_data_in(11315);
  VN1886_in0 <= VN_sign_in(11316) & VN_data_in(11316);
  VN1886_in1 <= VN_sign_in(11317) & VN_data_in(11317);
  VN1886_in2 <= VN_sign_in(11318) & VN_data_in(11318);
  VN1886_in3 <= VN_sign_in(11319) & VN_data_in(11319);
  VN1886_in4 <= VN_sign_in(11320) & VN_data_in(11320);
  VN1886_in5 <= VN_sign_in(11321) & VN_data_in(11321);
  VN1887_in0 <= VN_sign_in(11322) & VN_data_in(11322);
  VN1887_in1 <= VN_sign_in(11323) & VN_data_in(11323);
  VN1887_in2 <= VN_sign_in(11324) & VN_data_in(11324);
  VN1887_in3 <= VN_sign_in(11325) & VN_data_in(11325);
  VN1887_in4 <= VN_sign_in(11326) & VN_data_in(11326);
  VN1887_in5 <= VN_sign_in(11327) & VN_data_in(11327);
  VN1888_in0 <= VN_sign_in(11328) & VN_data_in(11328);
  VN1888_in1 <= VN_sign_in(11329) & VN_data_in(11329);
  VN1888_in2 <= VN_sign_in(11330) & VN_data_in(11330);
  VN1888_in3 <= VN_sign_in(11331) & VN_data_in(11331);
  VN1888_in4 <= VN_sign_in(11332) & VN_data_in(11332);
  VN1888_in5 <= VN_sign_in(11333) & VN_data_in(11333);
  VN1889_in0 <= VN_sign_in(11334) & VN_data_in(11334);
  VN1889_in1 <= VN_sign_in(11335) & VN_data_in(11335);
  VN1889_in2 <= VN_sign_in(11336) & VN_data_in(11336);
  VN1889_in3 <= VN_sign_in(11337) & VN_data_in(11337);
  VN1889_in4 <= VN_sign_in(11338) & VN_data_in(11338);
  VN1889_in5 <= VN_sign_in(11339) & VN_data_in(11339);
  VN1890_in0 <= VN_sign_in(11340) & VN_data_in(11340);
  VN1890_in1 <= VN_sign_in(11341) & VN_data_in(11341);
  VN1890_in2 <= VN_sign_in(11342) & VN_data_in(11342);
  VN1890_in3 <= VN_sign_in(11343) & VN_data_in(11343);
  VN1890_in4 <= VN_sign_in(11344) & VN_data_in(11344);
  VN1890_in5 <= VN_sign_in(11345) & VN_data_in(11345);
  VN1891_in0 <= VN_sign_in(11346) & VN_data_in(11346);
  VN1891_in1 <= VN_sign_in(11347) & VN_data_in(11347);
  VN1891_in2 <= VN_sign_in(11348) & VN_data_in(11348);
  VN1891_in3 <= VN_sign_in(11349) & VN_data_in(11349);
  VN1891_in4 <= VN_sign_in(11350) & VN_data_in(11350);
  VN1891_in5 <= VN_sign_in(11351) & VN_data_in(11351);
  VN1892_in0 <= VN_sign_in(11352) & VN_data_in(11352);
  VN1892_in1 <= VN_sign_in(11353) & VN_data_in(11353);
  VN1892_in2 <= VN_sign_in(11354) & VN_data_in(11354);
  VN1892_in3 <= VN_sign_in(11355) & VN_data_in(11355);
  VN1892_in4 <= VN_sign_in(11356) & VN_data_in(11356);
  VN1892_in5 <= VN_sign_in(11357) & VN_data_in(11357);
  VN1893_in0 <= VN_sign_in(11358) & VN_data_in(11358);
  VN1893_in1 <= VN_sign_in(11359) & VN_data_in(11359);
  VN1893_in2 <= VN_sign_in(11360) & VN_data_in(11360);
  VN1893_in3 <= VN_sign_in(11361) & VN_data_in(11361);
  VN1893_in4 <= VN_sign_in(11362) & VN_data_in(11362);
  VN1893_in5 <= VN_sign_in(11363) & VN_data_in(11363);
  VN1894_in0 <= VN_sign_in(11364) & VN_data_in(11364);
  VN1894_in1 <= VN_sign_in(11365) & VN_data_in(11365);
  VN1894_in2 <= VN_sign_in(11366) & VN_data_in(11366);
  VN1894_in3 <= VN_sign_in(11367) & VN_data_in(11367);
  VN1894_in4 <= VN_sign_in(11368) & VN_data_in(11368);
  VN1894_in5 <= VN_sign_in(11369) & VN_data_in(11369);
  VN1895_in0 <= VN_sign_in(11370) & VN_data_in(11370);
  VN1895_in1 <= VN_sign_in(11371) & VN_data_in(11371);
  VN1895_in2 <= VN_sign_in(11372) & VN_data_in(11372);
  VN1895_in3 <= VN_sign_in(11373) & VN_data_in(11373);
  VN1895_in4 <= VN_sign_in(11374) & VN_data_in(11374);
  VN1895_in5 <= VN_sign_in(11375) & VN_data_in(11375);
  VN1896_in0 <= VN_sign_in(11376) & VN_data_in(11376);
  VN1896_in1 <= VN_sign_in(11377) & VN_data_in(11377);
  VN1896_in2 <= VN_sign_in(11378) & VN_data_in(11378);
  VN1896_in3 <= VN_sign_in(11379) & VN_data_in(11379);
  VN1896_in4 <= VN_sign_in(11380) & VN_data_in(11380);
  VN1896_in5 <= VN_sign_in(11381) & VN_data_in(11381);
  VN1897_in0 <= VN_sign_in(11382) & VN_data_in(11382);
  VN1897_in1 <= VN_sign_in(11383) & VN_data_in(11383);
  VN1897_in2 <= VN_sign_in(11384) & VN_data_in(11384);
  VN1897_in3 <= VN_sign_in(11385) & VN_data_in(11385);
  VN1897_in4 <= VN_sign_in(11386) & VN_data_in(11386);
  VN1897_in5 <= VN_sign_in(11387) & VN_data_in(11387);
  VN1898_in0 <= VN_sign_in(11388) & VN_data_in(11388);
  VN1898_in1 <= VN_sign_in(11389) & VN_data_in(11389);
  VN1898_in2 <= VN_sign_in(11390) & VN_data_in(11390);
  VN1898_in3 <= VN_sign_in(11391) & VN_data_in(11391);
  VN1898_in4 <= VN_sign_in(11392) & VN_data_in(11392);
  VN1898_in5 <= VN_sign_in(11393) & VN_data_in(11393);
  VN1899_in0 <= VN_sign_in(11394) & VN_data_in(11394);
  VN1899_in1 <= VN_sign_in(11395) & VN_data_in(11395);
  VN1899_in2 <= VN_sign_in(11396) & VN_data_in(11396);
  VN1899_in3 <= VN_sign_in(11397) & VN_data_in(11397);
  VN1899_in4 <= VN_sign_in(11398) & VN_data_in(11398);
  VN1899_in5 <= VN_sign_in(11399) & VN_data_in(11399);
  VN1900_in0 <= VN_sign_in(11400) & VN_data_in(11400);
  VN1900_in1 <= VN_sign_in(11401) & VN_data_in(11401);
  VN1900_in2 <= VN_sign_in(11402) & VN_data_in(11402);
  VN1900_in3 <= VN_sign_in(11403) & VN_data_in(11403);
  VN1900_in4 <= VN_sign_in(11404) & VN_data_in(11404);
  VN1900_in5 <= VN_sign_in(11405) & VN_data_in(11405);
  VN1901_in0 <= VN_sign_in(11406) & VN_data_in(11406);
  VN1901_in1 <= VN_sign_in(11407) & VN_data_in(11407);
  VN1901_in2 <= VN_sign_in(11408) & VN_data_in(11408);
  VN1901_in3 <= VN_sign_in(11409) & VN_data_in(11409);
  VN1901_in4 <= VN_sign_in(11410) & VN_data_in(11410);
  VN1901_in5 <= VN_sign_in(11411) & VN_data_in(11411);
  VN1902_in0 <= VN_sign_in(11412) & VN_data_in(11412);
  VN1902_in1 <= VN_sign_in(11413) & VN_data_in(11413);
  VN1902_in2 <= VN_sign_in(11414) & VN_data_in(11414);
  VN1902_in3 <= VN_sign_in(11415) & VN_data_in(11415);
  VN1902_in4 <= VN_sign_in(11416) & VN_data_in(11416);
  VN1902_in5 <= VN_sign_in(11417) & VN_data_in(11417);
  VN1903_in0 <= VN_sign_in(11418) & VN_data_in(11418);
  VN1903_in1 <= VN_sign_in(11419) & VN_data_in(11419);
  VN1903_in2 <= VN_sign_in(11420) & VN_data_in(11420);
  VN1903_in3 <= VN_sign_in(11421) & VN_data_in(11421);
  VN1903_in4 <= VN_sign_in(11422) & VN_data_in(11422);
  VN1903_in5 <= VN_sign_in(11423) & VN_data_in(11423);
  VN1904_in0 <= VN_sign_in(11424) & VN_data_in(11424);
  VN1904_in1 <= VN_sign_in(11425) & VN_data_in(11425);
  VN1904_in2 <= VN_sign_in(11426) & VN_data_in(11426);
  VN1904_in3 <= VN_sign_in(11427) & VN_data_in(11427);
  VN1904_in4 <= VN_sign_in(11428) & VN_data_in(11428);
  VN1904_in5 <= VN_sign_in(11429) & VN_data_in(11429);
  VN1905_in0 <= VN_sign_in(11430) & VN_data_in(11430);
  VN1905_in1 <= VN_sign_in(11431) & VN_data_in(11431);
  VN1905_in2 <= VN_sign_in(11432) & VN_data_in(11432);
  VN1905_in3 <= VN_sign_in(11433) & VN_data_in(11433);
  VN1905_in4 <= VN_sign_in(11434) & VN_data_in(11434);
  VN1905_in5 <= VN_sign_in(11435) & VN_data_in(11435);
  VN1906_in0 <= VN_sign_in(11436) & VN_data_in(11436);
  VN1906_in1 <= VN_sign_in(11437) & VN_data_in(11437);
  VN1906_in2 <= VN_sign_in(11438) & VN_data_in(11438);
  VN1906_in3 <= VN_sign_in(11439) & VN_data_in(11439);
  VN1906_in4 <= VN_sign_in(11440) & VN_data_in(11440);
  VN1906_in5 <= VN_sign_in(11441) & VN_data_in(11441);
  VN1907_in0 <= VN_sign_in(11442) & VN_data_in(11442);
  VN1907_in1 <= VN_sign_in(11443) & VN_data_in(11443);
  VN1907_in2 <= VN_sign_in(11444) & VN_data_in(11444);
  VN1907_in3 <= VN_sign_in(11445) & VN_data_in(11445);
  VN1907_in4 <= VN_sign_in(11446) & VN_data_in(11446);
  VN1907_in5 <= VN_sign_in(11447) & VN_data_in(11447);
  VN1908_in0 <= VN_sign_in(11448) & VN_data_in(11448);
  VN1908_in1 <= VN_sign_in(11449) & VN_data_in(11449);
  VN1908_in2 <= VN_sign_in(11450) & VN_data_in(11450);
  VN1908_in3 <= VN_sign_in(11451) & VN_data_in(11451);
  VN1908_in4 <= VN_sign_in(11452) & VN_data_in(11452);
  VN1908_in5 <= VN_sign_in(11453) & VN_data_in(11453);
  VN1909_in0 <= VN_sign_in(11454) & VN_data_in(11454);
  VN1909_in1 <= VN_sign_in(11455) & VN_data_in(11455);
  VN1909_in2 <= VN_sign_in(11456) & VN_data_in(11456);
  VN1909_in3 <= VN_sign_in(11457) & VN_data_in(11457);
  VN1909_in4 <= VN_sign_in(11458) & VN_data_in(11458);
  VN1909_in5 <= VN_sign_in(11459) & VN_data_in(11459);
  VN1910_in0 <= VN_sign_in(11460) & VN_data_in(11460);
  VN1910_in1 <= VN_sign_in(11461) & VN_data_in(11461);
  VN1910_in2 <= VN_sign_in(11462) & VN_data_in(11462);
  VN1910_in3 <= VN_sign_in(11463) & VN_data_in(11463);
  VN1910_in4 <= VN_sign_in(11464) & VN_data_in(11464);
  VN1910_in5 <= VN_sign_in(11465) & VN_data_in(11465);
  VN1911_in0 <= VN_sign_in(11466) & VN_data_in(11466);
  VN1911_in1 <= VN_sign_in(11467) & VN_data_in(11467);
  VN1911_in2 <= VN_sign_in(11468) & VN_data_in(11468);
  VN1911_in3 <= VN_sign_in(11469) & VN_data_in(11469);
  VN1911_in4 <= VN_sign_in(11470) & VN_data_in(11470);
  VN1911_in5 <= VN_sign_in(11471) & VN_data_in(11471);
  VN1912_in0 <= VN_sign_in(11472) & VN_data_in(11472);
  VN1912_in1 <= VN_sign_in(11473) & VN_data_in(11473);
  VN1912_in2 <= VN_sign_in(11474) & VN_data_in(11474);
  VN1912_in3 <= VN_sign_in(11475) & VN_data_in(11475);
  VN1912_in4 <= VN_sign_in(11476) & VN_data_in(11476);
  VN1912_in5 <= VN_sign_in(11477) & VN_data_in(11477);
  VN1913_in0 <= VN_sign_in(11478) & VN_data_in(11478);
  VN1913_in1 <= VN_sign_in(11479) & VN_data_in(11479);
  VN1913_in2 <= VN_sign_in(11480) & VN_data_in(11480);
  VN1913_in3 <= VN_sign_in(11481) & VN_data_in(11481);
  VN1913_in4 <= VN_sign_in(11482) & VN_data_in(11482);
  VN1913_in5 <= VN_sign_in(11483) & VN_data_in(11483);
  VN1914_in0 <= VN_sign_in(11484) & VN_data_in(11484);
  VN1914_in1 <= VN_sign_in(11485) & VN_data_in(11485);
  VN1914_in2 <= VN_sign_in(11486) & VN_data_in(11486);
  VN1914_in3 <= VN_sign_in(11487) & VN_data_in(11487);
  VN1914_in4 <= VN_sign_in(11488) & VN_data_in(11488);
  VN1914_in5 <= VN_sign_in(11489) & VN_data_in(11489);
  VN1915_in0 <= VN_sign_in(11490) & VN_data_in(11490);
  VN1915_in1 <= VN_sign_in(11491) & VN_data_in(11491);
  VN1915_in2 <= VN_sign_in(11492) & VN_data_in(11492);
  VN1915_in3 <= VN_sign_in(11493) & VN_data_in(11493);
  VN1915_in4 <= VN_sign_in(11494) & VN_data_in(11494);
  VN1915_in5 <= VN_sign_in(11495) & VN_data_in(11495);
  VN1916_in0 <= VN_sign_in(11496) & VN_data_in(11496);
  VN1916_in1 <= VN_sign_in(11497) & VN_data_in(11497);
  VN1916_in2 <= VN_sign_in(11498) & VN_data_in(11498);
  VN1916_in3 <= VN_sign_in(11499) & VN_data_in(11499);
  VN1916_in4 <= VN_sign_in(11500) & VN_data_in(11500);
  VN1916_in5 <= VN_sign_in(11501) & VN_data_in(11501);
  VN1917_in0 <= VN_sign_in(11502) & VN_data_in(11502);
  VN1917_in1 <= VN_sign_in(11503) & VN_data_in(11503);
  VN1917_in2 <= VN_sign_in(11504) & VN_data_in(11504);
  VN1917_in3 <= VN_sign_in(11505) & VN_data_in(11505);
  VN1917_in4 <= VN_sign_in(11506) & VN_data_in(11506);
  VN1917_in5 <= VN_sign_in(11507) & VN_data_in(11507);
  VN1918_in0 <= VN_sign_in(11508) & VN_data_in(11508);
  VN1918_in1 <= VN_sign_in(11509) & VN_data_in(11509);
  VN1918_in2 <= VN_sign_in(11510) & VN_data_in(11510);
  VN1918_in3 <= VN_sign_in(11511) & VN_data_in(11511);
  VN1918_in4 <= VN_sign_in(11512) & VN_data_in(11512);
  VN1918_in5 <= VN_sign_in(11513) & VN_data_in(11513);
  VN1919_in0 <= VN_sign_in(11514) & VN_data_in(11514);
  VN1919_in1 <= VN_sign_in(11515) & VN_data_in(11515);
  VN1919_in2 <= VN_sign_in(11516) & VN_data_in(11516);
  VN1919_in3 <= VN_sign_in(11517) & VN_data_in(11517);
  VN1919_in4 <= VN_sign_in(11518) & VN_data_in(11518);
  VN1919_in5 <= VN_sign_in(11519) & VN_data_in(11519);
  VN1920_in0 <= VN_sign_in(11520) & VN_data_in(11520);
  VN1920_in1 <= VN_sign_in(11521) & VN_data_in(11521);
  VN1920_in2 <= VN_sign_in(11522) & VN_data_in(11522);
  VN1920_in3 <= VN_sign_in(11523) & VN_data_in(11523);
  VN1920_in4 <= VN_sign_in(11524) & VN_data_in(11524);
  VN1920_in5 <= VN_sign_in(11525) & VN_data_in(11525);
  VN1921_in0 <= VN_sign_in(11526) & VN_data_in(11526);
  VN1921_in1 <= VN_sign_in(11527) & VN_data_in(11527);
  VN1921_in2 <= VN_sign_in(11528) & VN_data_in(11528);
  VN1921_in3 <= VN_sign_in(11529) & VN_data_in(11529);
  VN1921_in4 <= VN_sign_in(11530) & VN_data_in(11530);
  VN1921_in5 <= VN_sign_in(11531) & VN_data_in(11531);
  VN1922_in0 <= VN_sign_in(11532) & VN_data_in(11532);
  VN1922_in1 <= VN_sign_in(11533) & VN_data_in(11533);
  VN1922_in2 <= VN_sign_in(11534) & VN_data_in(11534);
  VN1922_in3 <= VN_sign_in(11535) & VN_data_in(11535);
  VN1922_in4 <= VN_sign_in(11536) & VN_data_in(11536);
  VN1922_in5 <= VN_sign_in(11537) & VN_data_in(11537);
  VN1923_in0 <= VN_sign_in(11538) & VN_data_in(11538);
  VN1923_in1 <= VN_sign_in(11539) & VN_data_in(11539);
  VN1923_in2 <= VN_sign_in(11540) & VN_data_in(11540);
  VN1923_in3 <= VN_sign_in(11541) & VN_data_in(11541);
  VN1923_in4 <= VN_sign_in(11542) & VN_data_in(11542);
  VN1923_in5 <= VN_sign_in(11543) & VN_data_in(11543);
  VN1924_in0 <= VN_sign_in(11544) & VN_data_in(11544);
  VN1924_in1 <= VN_sign_in(11545) & VN_data_in(11545);
  VN1924_in2 <= VN_sign_in(11546) & VN_data_in(11546);
  VN1924_in3 <= VN_sign_in(11547) & VN_data_in(11547);
  VN1924_in4 <= VN_sign_in(11548) & VN_data_in(11548);
  VN1924_in5 <= VN_sign_in(11549) & VN_data_in(11549);
  VN1925_in0 <= VN_sign_in(11550) & VN_data_in(11550);
  VN1925_in1 <= VN_sign_in(11551) & VN_data_in(11551);
  VN1925_in2 <= VN_sign_in(11552) & VN_data_in(11552);
  VN1925_in3 <= VN_sign_in(11553) & VN_data_in(11553);
  VN1925_in4 <= VN_sign_in(11554) & VN_data_in(11554);
  VN1925_in5 <= VN_sign_in(11555) & VN_data_in(11555);
  VN1926_in0 <= VN_sign_in(11556) & VN_data_in(11556);
  VN1926_in1 <= VN_sign_in(11557) & VN_data_in(11557);
  VN1926_in2 <= VN_sign_in(11558) & VN_data_in(11558);
  VN1926_in3 <= VN_sign_in(11559) & VN_data_in(11559);
  VN1926_in4 <= VN_sign_in(11560) & VN_data_in(11560);
  VN1926_in5 <= VN_sign_in(11561) & VN_data_in(11561);
  VN1927_in0 <= VN_sign_in(11562) & VN_data_in(11562);
  VN1927_in1 <= VN_sign_in(11563) & VN_data_in(11563);
  VN1927_in2 <= VN_sign_in(11564) & VN_data_in(11564);
  VN1927_in3 <= VN_sign_in(11565) & VN_data_in(11565);
  VN1927_in4 <= VN_sign_in(11566) & VN_data_in(11566);
  VN1927_in5 <= VN_sign_in(11567) & VN_data_in(11567);
  VN1928_in0 <= VN_sign_in(11568) & VN_data_in(11568);
  VN1928_in1 <= VN_sign_in(11569) & VN_data_in(11569);
  VN1928_in2 <= VN_sign_in(11570) & VN_data_in(11570);
  VN1928_in3 <= VN_sign_in(11571) & VN_data_in(11571);
  VN1928_in4 <= VN_sign_in(11572) & VN_data_in(11572);
  VN1928_in5 <= VN_sign_in(11573) & VN_data_in(11573);
  VN1929_in0 <= VN_sign_in(11574) & VN_data_in(11574);
  VN1929_in1 <= VN_sign_in(11575) & VN_data_in(11575);
  VN1929_in2 <= VN_sign_in(11576) & VN_data_in(11576);
  VN1929_in3 <= VN_sign_in(11577) & VN_data_in(11577);
  VN1929_in4 <= VN_sign_in(11578) & VN_data_in(11578);
  VN1929_in5 <= VN_sign_in(11579) & VN_data_in(11579);
  VN1930_in0 <= VN_sign_in(11580) & VN_data_in(11580);
  VN1930_in1 <= VN_sign_in(11581) & VN_data_in(11581);
  VN1930_in2 <= VN_sign_in(11582) & VN_data_in(11582);
  VN1930_in3 <= VN_sign_in(11583) & VN_data_in(11583);
  VN1930_in4 <= VN_sign_in(11584) & VN_data_in(11584);
  VN1930_in5 <= VN_sign_in(11585) & VN_data_in(11585);
  VN1931_in0 <= VN_sign_in(11586) & VN_data_in(11586);
  VN1931_in1 <= VN_sign_in(11587) & VN_data_in(11587);
  VN1931_in2 <= VN_sign_in(11588) & VN_data_in(11588);
  VN1931_in3 <= VN_sign_in(11589) & VN_data_in(11589);
  VN1931_in4 <= VN_sign_in(11590) & VN_data_in(11590);
  VN1931_in5 <= VN_sign_in(11591) & VN_data_in(11591);
  VN1932_in0 <= VN_sign_in(11592) & VN_data_in(11592);
  VN1932_in1 <= VN_sign_in(11593) & VN_data_in(11593);
  VN1932_in2 <= VN_sign_in(11594) & VN_data_in(11594);
  VN1932_in3 <= VN_sign_in(11595) & VN_data_in(11595);
  VN1932_in4 <= VN_sign_in(11596) & VN_data_in(11596);
  VN1932_in5 <= VN_sign_in(11597) & VN_data_in(11597);
  VN1933_in0 <= VN_sign_in(11598) & VN_data_in(11598);
  VN1933_in1 <= VN_sign_in(11599) & VN_data_in(11599);
  VN1933_in2 <= VN_sign_in(11600) & VN_data_in(11600);
  VN1933_in3 <= VN_sign_in(11601) & VN_data_in(11601);
  VN1933_in4 <= VN_sign_in(11602) & VN_data_in(11602);
  VN1933_in5 <= VN_sign_in(11603) & VN_data_in(11603);
  VN1934_in0 <= VN_sign_in(11604) & VN_data_in(11604);
  VN1934_in1 <= VN_sign_in(11605) & VN_data_in(11605);
  VN1934_in2 <= VN_sign_in(11606) & VN_data_in(11606);
  VN1934_in3 <= VN_sign_in(11607) & VN_data_in(11607);
  VN1934_in4 <= VN_sign_in(11608) & VN_data_in(11608);
  VN1934_in5 <= VN_sign_in(11609) & VN_data_in(11609);
  VN1935_in0 <= VN_sign_in(11610) & VN_data_in(11610);
  VN1935_in1 <= VN_sign_in(11611) & VN_data_in(11611);
  VN1935_in2 <= VN_sign_in(11612) & VN_data_in(11612);
  VN1935_in3 <= VN_sign_in(11613) & VN_data_in(11613);
  VN1935_in4 <= VN_sign_in(11614) & VN_data_in(11614);
  VN1935_in5 <= VN_sign_in(11615) & VN_data_in(11615);
  VN1936_in0 <= VN_sign_in(11616) & VN_data_in(11616);
  VN1936_in1 <= VN_sign_in(11617) & VN_data_in(11617);
  VN1936_in2 <= VN_sign_in(11618) & VN_data_in(11618);
  VN1936_in3 <= VN_sign_in(11619) & VN_data_in(11619);
  VN1936_in4 <= VN_sign_in(11620) & VN_data_in(11620);
  VN1936_in5 <= VN_sign_in(11621) & VN_data_in(11621);
  VN1937_in0 <= VN_sign_in(11622) & VN_data_in(11622);
  VN1937_in1 <= VN_sign_in(11623) & VN_data_in(11623);
  VN1937_in2 <= VN_sign_in(11624) & VN_data_in(11624);
  VN1937_in3 <= VN_sign_in(11625) & VN_data_in(11625);
  VN1937_in4 <= VN_sign_in(11626) & VN_data_in(11626);
  VN1937_in5 <= VN_sign_in(11627) & VN_data_in(11627);
  VN1938_in0 <= VN_sign_in(11628) & VN_data_in(11628);
  VN1938_in1 <= VN_sign_in(11629) & VN_data_in(11629);
  VN1938_in2 <= VN_sign_in(11630) & VN_data_in(11630);
  VN1938_in3 <= VN_sign_in(11631) & VN_data_in(11631);
  VN1938_in4 <= VN_sign_in(11632) & VN_data_in(11632);
  VN1938_in5 <= VN_sign_in(11633) & VN_data_in(11633);
  VN1939_in0 <= VN_sign_in(11634) & VN_data_in(11634);
  VN1939_in1 <= VN_sign_in(11635) & VN_data_in(11635);
  VN1939_in2 <= VN_sign_in(11636) & VN_data_in(11636);
  VN1939_in3 <= VN_sign_in(11637) & VN_data_in(11637);
  VN1939_in4 <= VN_sign_in(11638) & VN_data_in(11638);
  VN1939_in5 <= VN_sign_in(11639) & VN_data_in(11639);
  VN1940_in0 <= VN_sign_in(11640) & VN_data_in(11640);
  VN1940_in1 <= VN_sign_in(11641) & VN_data_in(11641);
  VN1940_in2 <= VN_sign_in(11642) & VN_data_in(11642);
  VN1940_in3 <= VN_sign_in(11643) & VN_data_in(11643);
  VN1940_in4 <= VN_sign_in(11644) & VN_data_in(11644);
  VN1940_in5 <= VN_sign_in(11645) & VN_data_in(11645);
  VN1941_in0 <= VN_sign_in(11646) & VN_data_in(11646);
  VN1941_in1 <= VN_sign_in(11647) & VN_data_in(11647);
  VN1941_in2 <= VN_sign_in(11648) & VN_data_in(11648);
  VN1941_in3 <= VN_sign_in(11649) & VN_data_in(11649);
  VN1941_in4 <= VN_sign_in(11650) & VN_data_in(11650);
  VN1941_in5 <= VN_sign_in(11651) & VN_data_in(11651);
  VN1942_in0 <= VN_sign_in(11652) & VN_data_in(11652);
  VN1942_in1 <= VN_sign_in(11653) & VN_data_in(11653);
  VN1942_in2 <= VN_sign_in(11654) & VN_data_in(11654);
  VN1942_in3 <= VN_sign_in(11655) & VN_data_in(11655);
  VN1942_in4 <= VN_sign_in(11656) & VN_data_in(11656);
  VN1942_in5 <= VN_sign_in(11657) & VN_data_in(11657);
  VN1943_in0 <= VN_sign_in(11658) & VN_data_in(11658);
  VN1943_in1 <= VN_sign_in(11659) & VN_data_in(11659);
  VN1943_in2 <= VN_sign_in(11660) & VN_data_in(11660);
  VN1943_in3 <= VN_sign_in(11661) & VN_data_in(11661);
  VN1943_in4 <= VN_sign_in(11662) & VN_data_in(11662);
  VN1943_in5 <= VN_sign_in(11663) & VN_data_in(11663);
  VN1944_in0 <= VN_sign_in(11664) & VN_data_in(11664);
  VN1944_in1 <= VN_sign_in(11665) & VN_data_in(11665);
  VN1944_in2 <= VN_sign_in(11666) & VN_data_in(11666);
  VN1944_in3 <= VN_sign_in(11667) & VN_data_in(11667);
  VN1944_in4 <= VN_sign_in(11668) & VN_data_in(11668);
  VN1944_in5 <= VN_sign_in(11669) & VN_data_in(11669);
  VN1945_in0 <= VN_sign_in(11670) & VN_data_in(11670);
  VN1945_in1 <= VN_sign_in(11671) & VN_data_in(11671);
  VN1945_in2 <= VN_sign_in(11672) & VN_data_in(11672);
  VN1945_in3 <= VN_sign_in(11673) & VN_data_in(11673);
  VN1945_in4 <= VN_sign_in(11674) & VN_data_in(11674);
  VN1945_in5 <= VN_sign_in(11675) & VN_data_in(11675);
  VN1946_in0 <= VN_sign_in(11676) & VN_data_in(11676);
  VN1946_in1 <= VN_sign_in(11677) & VN_data_in(11677);
  VN1946_in2 <= VN_sign_in(11678) & VN_data_in(11678);
  VN1946_in3 <= VN_sign_in(11679) & VN_data_in(11679);
  VN1946_in4 <= VN_sign_in(11680) & VN_data_in(11680);
  VN1946_in5 <= VN_sign_in(11681) & VN_data_in(11681);
  VN1947_in0 <= VN_sign_in(11682) & VN_data_in(11682);
  VN1947_in1 <= VN_sign_in(11683) & VN_data_in(11683);
  VN1947_in2 <= VN_sign_in(11684) & VN_data_in(11684);
  VN1947_in3 <= VN_sign_in(11685) & VN_data_in(11685);
  VN1947_in4 <= VN_sign_in(11686) & VN_data_in(11686);
  VN1947_in5 <= VN_sign_in(11687) & VN_data_in(11687);
  VN1948_in0 <= VN_sign_in(11688) & VN_data_in(11688);
  VN1948_in1 <= VN_sign_in(11689) & VN_data_in(11689);
  VN1948_in2 <= VN_sign_in(11690) & VN_data_in(11690);
  VN1948_in3 <= VN_sign_in(11691) & VN_data_in(11691);
  VN1948_in4 <= VN_sign_in(11692) & VN_data_in(11692);
  VN1948_in5 <= VN_sign_in(11693) & VN_data_in(11693);
  VN1949_in0 <= VN_sign_in(11694) & VN_data_in(11694);
  VN1949_in1 <= VN_sign_in(11695) & VN_data_in(11695);
  VN1949_in2 <= VN_sign_in(11696) & VN_data_in(11696);
  VN1949_in3 <= VN_sign_in(11697) & VN_data_in(11697);
  VN1949_in4 <= VN_sign_in(11698) & VN_data_in(11698);
  VN1949_in5 <= VN_sign_in(11699) & VN_data_in(11699);
  VN1950_in0 <= VN_sign_in(11700) & VN_data_in(11700);
  VN1950_in1 <= VN_sign_in(11701) & VN_data_in(11701);
  VN1950_in2 <= VN_sign_in(11702) & VN_data_in(11702);
  VN1950_in3 <= VN_sign_in(11703) & VN_data_in(11703);
  VN1950_in4 <= VN_sign_in(11704) & VN_data_in(11704);
  VN1950_in5 <= VN_sign_in(11705) & VN_data_in(11705);
  VN1951_in0 <= VN_sign_in(11706) & VN_data_in(11706);
  VN1951_in1 <= VN_sign_in(11707) & VN_data_in(11707);
  VN1951_in2 <= VN_sign_in(11708) & VN_data_in(11708);
  VN1951_in3 <= VN_sign_in(11709) & VN_data_in(11709);
  VN1951_in4 <= VN_sign_in(11710) & VN_data_in(11710);
  VN1951_in5 <= VN_sign_in(11711) & VN_data_in(11711);
  VN1952_in0 <= VN_sign_in(11712) & VN_data_in(11712);
  VN1952_in1 <= VN_sign_in(11713) & VN_data_in(11713);
  VN1952_in2 <= VN_sign_in(11714) & VN_data_in(11714);
  VN1952_in3 <= VN_sign_in(11715) & VN_data_in(11715);
  VN1952_in4 <= VN_sign_in(11716) & VN_data_in(11716);
  VN1952_in5 <= VN_sign_in(11717) & VN_data_in(11717);
  VN1953_in0 <= VN_sign_in(11718) & VN_data_in(11718);
  VN1953_in1 <= VN_sign_in(11719) & VN_data_in(11719);
  VN1953_in2 <= VN_sign_in(11720) & VN_data_in(11720);
  VN1953_in3 <= VN_sign_in(11721) & VN_data_in(11721);
  VN1953_in4 <= VN_sign_in(11722) & VN_data_in(11722);
  VN1953_in5 <= VN_sign_in(11723) & VN_data_in(11723);
  VN1954_in0 <= VN_sign_in(11724) & VN_data_in(11724);
  VN1954_in1 <= VN_sign_in(11725) & VN_data_in(11725);
  VN1954_in2 <= VN_sign_in(11726) & VN_data_in(11726);
  VN1954_in3 <= VN_sign_in(11727) & VN_data_in(11727);
  VN1954_in4 <= VN_sign_in(11728) & VN_data_in(11728);
  VN1954_in5 <= VN_sign_in(11729) & VN_data_in(11729);
  VN1955_in0 <= VN_sign_in(11730) & VN_data_in(11730);
  VN1955_in1 <= VN_sign_in(11731) & VN_data_in(11731);
  VN1955_in2 <= VN_sign_in(11732) & VN_data_in(11732);
  VN1955_in3 <= VN_sign_in(11733) & VN_data_in(11733);
  VN1955_in4 <= VN_sign_in(11734) & VN_data_in(11734);
  VN1955_in5 <= VN_sign_in(11735) & VN_data_in(11735);
  VN1956_in0 <= VN_sign_in(11736) & VN_data_in(11736);
  VN1956_in1 <= VN_sign_in(11737) & VN_data_in(11737);
  VN1956_in2 <= VN_sign_in(11738) & VN_data_in(11738);
  VN1956_in3 <= VN_sign_in(11739) & VN_data_in(11739);
  VN1956_in4 <= VN_sign_in(11740) & VN_data_in(11740);
  VN1956_in5 <= VN_sign_in(11741) & VN_data_in(11741);
  VN1957_in0 <= VN_sign_in(11742) & VN_data_in(11742);
  VN1957_in1 <= VN_sign_in(11743) & VN_data_in(11743);
  VN1957_in2 <= VN_sign_in(11744) & VN_data_in(11744);
  VN1957_in3 <= VN_sign_in(11745) & VN_data_in(11745);
  VN1957_in4 <= VN_sign_in(11746) & VN_data_in(11746);
  VN1957_in5 <= VN_sign_in(11747) & VN_data_in(11747);
  VN1958_in0 <= VN_sign_in(11748) & VN_data_in(11748);
  VN1958_in1 <= VN_sign_in(11749) & VN_data_in(11749);
  VN1958_in2 <= VN_sign_in(11750) & VN_data_in(11750);
  VN1958_in3 <= VN_sign_in(11751) & VN_data_in(11751);
  VN1958_in4 <= VN_sign_in(11752) & VN_data_in(11752);
  VN1958_in5 <= VN_sign_in(11753) & VN_data_in(11753);
  VN1959_in0 <= VN_sign_in(11754) & VN_data_in(11754);
  VN1959_in1 <= VN_sign_in(11755) & VN_data_in(11755);
  VN1959_in2 <= VN_sign_in(11756) & VN_data_in(11756);
  VN1959_in3 <= VN_sign_in(11757) & VN_data_in(11757);
  VN1959_in4 <= VN_sign_in(11758) & VN_data_in(11758);
  VN1959_in5 <= VN_sign_in(11759) & VN_data_in(11759);
  VN1960_in0 <= VN_sign_in(11760) & VN_data_in(11760);
  VN1960_in1 <= VN_sign_in(11761) & VN_data_in(11761);
  VN1960_in2 <= VN_sign_in(11762) & VN_data_in(11762);
  VN1960_in3 <= VN_sign_in(11763) & VN_data_in(11763);
  VN1960_in4 <= VN_sign_in(11764) & VN_data_in(11764);
  VN1960_in5 <= VN_sign_in(11765) & VN_data_in(11765);
  VN1961_in0 <= VN_sign_in(11766) & VN_data_in(11766);
  VN1961_in1 <= VN_sign_in(11767) & VN_data_in(11767);
  VN1961_in2 <= VN_sign_in(11768) & VN_data_in(11768);
  VN1961_in3 <= VN_sign_in(11769) & VN_data_in(11769);
  VN1961_in4 <= VN_sign_in(11770) & VN_data_in(11770);
  VN1961_in5 <= VN_sign_in(11771) & VN_data_in(11771);
  VN1962_in0 <= VN_sign_in(11772) & VN_data_in(11772);
  VN1962_in1 <= VN_sign_in(11773) & VN_data_in(11773);
  VN1962_in2 <= VN_sign_in(11774) & VN_data_in(11774);
  VN1962_in3 <= VN_sign_in(11775) & VN_data_in(11775);
  VN1962_in4 <= VN_sign_in(11776) & VN_data_in(11776);
  VN1962_in5 <= VN_sign_in(11777) & VN_data_in(11777);
  VN1963_in0 <= VN_sign_in(11778) & VN_data_in(11778);
  VN1963_in1 <= VN_sign_in(11779) & VN_data_in(11779);
  VN1963_in2 <= VN_sign_in(11780) & VN_data_in(11780);
  VN1963_in3 <= VN_sign_in(11781) & VN_data_in(11781);
  VN1963_in4 <= VN_sign_in(11782) & VN_data_in(11782);
  VN1963_in5 <= VN_sign_in(11783) & VN_data_in(11783);
  VN1964_in0 <= VN_sign_in(11784) & VN_data_in(11784);
  VN1964_in1 <= VN_sign_in(11785) & VN_data_in(11785);
  VN1964_in2 <= VN_sign_in(11786) & VN_data_in(11786);
  VN1964_in3 <= VN_sign_in(11787) & VN_data_in(11787);
  VN1964_in4 <= VN_sign_in(11788) & VN_data_in(11788);
  VN1964_in5 <= VN_sign_in(11789) & VN_data_in(11789);
  VN1965_in0 <= VN_sign_in(11790) & VN_data_in(11790);
  VN1965_in1 <= VN_sign_in(11791) & VN_data_in(11791);
  VN1965_in2 <= VN_sign_in(11792) & VN_data_in(11792);
  VN1965_in3 <= VN_sign_in(11793) & VN_data_in(11793);
  VN1965_in4 <= VN_sign_in(11794) & VN_data_in(11794);
  VN1965_in5 <= VN_sign_in(11795) & VN_data_in(11795);
  VN1966_in0 <= VN_sign_in(11796) & VN_data_in(11796);
  VN1966_in1 <= VN_sign_in(11797) & VN_data_in(11797);
  VN1966_in2 <= VN_sign_in(11798) & VN_data_in(11798);
  VN1966_in3 <= VN_sign_in(11799) & VN_data_in(11799);
  VN1966_in4 <= VN_sign_in(11800) & VN_data_in(11800);
  VN1966_in5 <= VN_sign_in(11801) & VN_data_in(11801);
  VN1967_in0 <= VN_sign_in(11802) & VN_data_in(11802);
  VN1967_in1 <= VN_sign_in(11803) & VN_data_in(11803);
  VN1967_in2 <= VN_sign_in(11804) & VN_data_in(11804);
  VN1967_in3 <= VN_sign_in(11805) & VN_data_in(11805);
  VN1967_in4 <= VN_sign_in(11806) & VN_data_in(11806);
  VN1967_in5 <= VN_sign_in(11807) & VN_data_in(11807);
  VN1968_in0 <= VN_sign_in(11808) & VN_data_in(11808);
  VN1968_in1 <= VN_sign_in(11809) & VN_data_in(11809);
  VN1968_in2 <= VN_sign_in(11810) & VN_data_in(11810);
  VN1968_in3 <= VN_sign_in(11811) & VN_data_in(11811);
  VN1968_in4 <= VN_sign_in(11812) & VN_data_in(11812);
  VN1968_in5 <= VN_sign_in(11813) & VN_data_in(11813);
  VN1969_in0 <= VN_sign_in(11814) & VN_data_in(11814);
  VN1969_in1 <= VN_sign_in(11815) & VN_data_in(11815);
  VN1969_in2 <= VN_sign_in(11816) & VN_data_in(11816);
  VN1969_in3 <= VN_sign_in(11817) & VN_data_in(11817);
  VN1969_in4 <= VN_sign_in(11818) & VN_data_in(11818);
  VN1969_in5 <= VN_sign_in(11819) & VN_data_in(11819);
  VN1970_in0 <= VN_sign_in(11820) & VN_data_in(11820);
  VN1970_in1 <= VN_sign_in(11821) & VN_data_in(11821);
  VN1970_in2 <= VN_sign_in(11822) & VN_data_in(11822);
  VN1970_in3 <= VN_sign_in(11823) & VN_data_in(11823);
  VN1970_in4 <= VN_sign_in(11824) & VN_data_in(11824);
  VN1970_in5 <= VN_sign_in(11825) & VN_data_in(11825);
  VN1971_in0 <= VN_sign_in(11826) & VN_data_in(11826);
  VN1971_in1 <= VN_sign_in(11827) & VN_data_in(11827);
  VN1971_in2 <= VN_sign_in(11828) & VN_data_in(11828);
  VN1971_in3 <= VN_sign_in(11829) & VN_data_in(11829);
  VN1971_in4 <= VN_sign_in(11830) & VN_data_in(11830);
  VN1971_in5 <= VN_sign_in(11831) & VN_data_in(11831);
  VN1972_in0 <= VN_sign_in(11832) & VN_data_in(11832);
  VN1972_in1 <= VN_sign_in(11833) & VN_data_in(11833);
  VN1972_in2 <= VN_sign_in(11834) & VN_data_in(11834);
  VN1972_in3 <= VN_sign_in(11835) & VN_data_in(11835);
  VN1972_in4 <= VN_sign_in(11836) & VN_data_in(11836);
  VN1972_in5 <= VN_sign_in(11837) & VN_data_in(11837);
  VN1973_in0 <= VN_sign_in(11838) & VN_data_in(11838);
  VN1973_in1 <= VN_sign_in(11839) & VN_data_in(11839);
  VN1973_in2 <= VN_sign_in(11840) & VN_data_in(11840);
  VN1973_in3 <= VN_sign_in(11841) & VN_data_in(11841);
  VN1973_in4 <= VN_sign_in(11842) & VN_data_in(11842);
  VN1973_in5 <= VN_sign_in(11843) & VN_data_in(11843);
  VN1974_in0 <= VN_sign_in(11844) & VN_data_in(11844);
  VN1974_in1 <= VN_sign_in(11845) & VN_data_in(11845);
  VN1974_in2 <= VN_sign_in(11846) & VN_data_in(11846);
  VN1974_in3 <= VN_sign_in(11847) & VN_data_in(11847);
  VN1974_in4 <= VN_sign_in(11848) & VN_data_in(11848);
  VN1974_in5 <= VN_sign_in(11849) & VN_data_in(11849);
  VN1975_in0 <= VN_sign_in(11850) & VN_data_in(11850);
  VN1975_in1 <= VN_sign_in(11851) & VN_data_in(11851);
  VN1975_in2 <= VN_sign_in(11852) & VN_data_in(11852);
  VN1975_in3 <= VN_sign_in(11853) & VN_data_in(11853);
  VN1975_in4 <= VN_sign_in(11854) & VN_data_in(11854);
  VN1975_in5 <= VN_sign_in(11855) & VN_data_in(11855);
  VN1976_in0 <= VN_sign_in(11856) & VN_data_in(11856);
  VN1976_in1 <= VN_sign_in(11857) & VN_data_in(11857);
  VN1976_in2 <= VN_sign_in(11858) & VN_data_in(11858);
  VN1976_in3 <= VN_sign_in(11859) & VN_data_in(11859);
  VN1976_in4 <= VN_sign_in(11860) & VN_data_in(11860);
  VN1976_in5 <= VN_sign_in(11861) & VN_data_in(11861);
  VN1977_in0 <= VN_sign_in(11862) & VN_data_in(11862);
  VN1977_in1 <= VN_sign_in(11863) & VN_data_in(11863);
  VN1977_in2 <= VN_sign_in(11864) & VN_data_in(11864);
  VN1977_in3 <= VN_sign_in(11865) & VN_data_in(11865);
  VN1977_in4 <= VN_sign_in(11866) & VN_data_in(11866);
  VN1977_in5 <= VN_sign_in(11867) & VN_data_in(11867);
  VN1978_in0 <= VN_sign_in(11868) & VN_data_in(11868);
  VN1978_in1 <= VN_sign_in(11869) & VN_data_in(11869);
  VN1978_in2 <= VN_sign_in(11870) & VN_data_in(11870);
  VN1978_in3 <= VN_sign_in(11871) & VN_data_in(11871);
  VN1978_in4 <= VN_sign_in(11872) & VN_data_in(11872);
  VN1978_in5 <= VN_sign_in(11873) & VN_data_in(11873);
  VN1979_in0 <= VN_sign_in(11874) & VN_data_in(11874);
  VN1979_in1 <= VN_sign_in(11875) & VN_data_in(11875);
  VN1979_in2 <= VN_sign_in(11876) & VN_data_in(11876);
  VN1979_in3 <= VN_sign_in(11877) & VN_data_in(11877);
  VN1979_in4 <= VN_sign_in(11878) & VN_data_in(11878);
  VN1979_in5 <= VN_sign_in(11879) & VN_data_in(11879);
  VN1980_in0 <= VN_sign_in(11880) & VN_data_in(11880);
  VN1980_in1 <= VN_sign_in(11881) & VN_data_in(11881);
  VN1980_in2 <= VN_sign_in(11882) & VN_data_in(11882);
  VN1980_in3 <= VN_sign_in(11883) & VN_data_in(11883);
  VN1980_in4 <= VN_sign_in(11884) & VN_data_in(11884);
  VN1980_in5 <= VN_sign_in(11885) & VN_data_in(11885);
  VN1981_in0 <= VN_sign_in(11886) & VN_data_in(11886);
  VN1981_in1 <= VN_sign_in(11887) & VN_data_in(11887);
  VN1981_in2 <= VN_sign_in(11888) & VN_data_in(11888);
  VN1981_in3 <= VN_sign_in(11889) & VN_data_in(11889);
  VN1981_in4 <= VN_sign_in(11890) & VN_data_in(11890);
  VN1981_in5 <= VN_sign_in(11891) & VN_data_in(11891);
  VN1982_in0 <= VN_sign_in(11892) & VN_data_in(11892);
  VN1982_in1 <= VN_sign_in(11893) & VN_data_in(11893);
  VN1982_in2 <= VN_sign_in(11894) & VN_data_in(11894);
  VN1982_in3 <= VN_sign_in(11895) & VN_data_in(11895);
  VN1982_in4 <= VN_sign_in(11896) & VN_data_in(11896);
  VN1982_in5 <= VN_sign_in(11897) & VN_data_in(11897);
  VN1983_in0 <= VN_sign_in(11898) & VN_data_in(11898);
  VN1983_in1 <= VN_sign_in(11899) & VN_data_in(11899);
  VN1983_in2 <= VN_sign_in(11900) & VN_data_in(11900);
  VN1983_in3 <= VN_sign_in(11901) & VN_data_in(11901);
  VN1983_in4 <= VN_sign_in(11902) & VN_data_in(11902);
  VN1983_in5 <= VN_sign_in(11903) & VN_data_in(11903);
  VN1984_in0 <= VN_sign_in(11904) & VN_data_in(11904);
  VN1984_in1 <= VN_sign_in(11905) & VN_data_in(11905);
  VN1984_in2 <= VN_sign_in(11906) & VN_data_in(11906);
  VN1984_in3 <= VN_sign_in(11907) & VN_data_in(11907);
  VN1984_in4 <= VN_sign_in(11908) & VN_data_in(11908);
  VN1984_in5 <= VN_sign_in(11909) & VN_data_in(11909);
  VN1985_in0 <= VN_sign_in(11910) & VN_data_in(11910);
  VN1985_in1 <= VN_sign_in(11911) & VN_data_in(11911);
  VN1985_in2 <= VN_sign_in(11912) & VN_data_in(11912);
  VN1985_in3 <= VN_sign_in(11913) & VN_data_in(11913);
  VN1985_in4 <= VN_sign_in(11914) & VN_data_in(11914);
  VN1985_in5 <= VN_sign_in(11915) & VN_data_in(11915);
  VN1986_in0 <= VN_sign_in(11916) & VN_data_in(11916);
  VN1986_in1 <= VN_sign_in(11917) & VN_data_in(11917);
  VN1986_in2 <= VN_sign_in(11918) & VN_data_in(11918);
  VN1986_in3 <= VN_sign_in(11919) & VN_data_in(11919);
  VN1986_in4 <= VN_sign_in(11920) & VN_data_in(11920);
  VN1986_in5 <= VN_sign_in(11921) & VN_data_in(11921);
  VN1987_in0 <= VN_sign_in(11922) & VN_data_in(11922);
  VN1987_in1 <= VN_sign_in(11923) & VN_data_in(11923);
  VN1987_in2 <= VN_sign_in(11924) & VN_data_in(11924);
  VN1987_in3 <= VN_sign_in(11925) & VN_data_in(11925);
  VN1987_in4 <= VN_sign_in(11926) & VN_data_in(11926);
  VN1987_in5 <= VN_sign_in(11927) & VN_data_in(11927);
  VN1988_in0 <= VN_sign_in(11928) & VN_data_in(11928);
  VN1988_in1 <= VN_sign_in(11929) & VN_data_in(11929);
  VN1988_in2 <= VN_sign_in(11930) & VN_data_in(11930);
  VN1988_in3 <= VN_sign_in(11931) & VN_data_in(11931);
  VN1988_in4 <= VN_sign_in(11932) & VN_data_in(11932);
  VN1988_in5 <= VN_sign_in(11933) & VN_data_in(11933);
  VN1989_in0 <= VN_sign_in(11934) & VN_data_in(11934);
  VN1989_in1 <= VN_sign_in(11935) & VN_data_in(11935);
  VN1989_in2 <= VN_sign_in(11936) & VN_data_in(11936);
  VN1989_in3 <= VN_sign_in(11937) & VN_data_in(11937);
  VN1989_in4 <= VN_sign_in(11938) & VN_data_in(11938);
  VN1989_in5 <= VN_sign_in(11939) & VN_data_in(11939);
  VN1990_in0 <= VN_sign_in(11940) & VN_data_in(11940);
  VN1990_in1 <= VN_sign_in(11941) & VN_data_in(11941);
  VN1990_in2 <= VN_sign_in(11942) & VN_data_in(11942);
  VN1990_in3 <= VN_sign_in(11943) & VN_data_in(11943);
  VN1990_in4 <= VN_sign_in(11944) & VN_data_in(11944);
  VN1990_in5 <= VN_sign_in(11945) & VN_data_in(11945);
  VN1991_in0 <= VN_sign_in(11946) & VN_data_in(11946);
  VN1991_in1 <= VN_sign_in(11947) & VN_data_in(11947);
  VN1991_in2 <= VN_sign_in(11948) & VN_data_in(11948);
  VN1991_in3 <= VN_sign_in(11949) & VN_data_in(11949);
  VN1991_in4 <= VN_sign_in(11950) & VN_data_in(11950);
  VN1991_in5 <= VN_sign_in(11951) & VN_data_in(11951);
  VN1992_in0 <= VN_sign_in(11952) & VN_data_in(11952);
  VN1992_in1 <= VN_sign_in(11953) & VN_data_in(11953);
  VN1992_in2 <= VN_sign_in(11954) & VN_data_in(11954);
  VN1992_in3 <= VN_sign_in(11955) & VN_data_in(11955);
  VN1992_in4 <= VN_sign_in(11956) & VN_data_in(11956);
  VN1992_in5 <= VN_sign_in(11957) & VN_data_in(11957);
  VN1993_in0 <= VN_sign_in(11958) & VN_data_in(11958);
  VN1993_in1 <= VN_sign_in(11959) & VN_data_in(11959);
  VN1993_in2 <= VN_sign_in(11960) & VN_data_in(11960);
  VN1993_in3 <= VN_sign_in(11961) & VN_data_in(11961);
  VN1993_in4 <= VN_sign_in(11962) & VN_data_in(11962);
  VN1993_in5 <= VN_sign_in(11963) & VN_data_in(11963);
  VN1994_in0 <= VN_sign_in(11964) & VN_data_in(11964);
  VN1994_in1 <= VN_sign_in(11965) & VN_data_in(11965);
  VN1994_in2 <= VN_sign_in(11966) & VN_data_in(11966);
  VN1994_in3 <= VN_sign_in(11967) & VN_data_in(11967);
  VN1994_in4 <= VN_sign_in(11968) & VN_data_in(11968);
  VN1994_in5 <= VN_sign_in(11969) & VN_data_in(11969);
  VN1995_in0 <= VN_sign_in(11970) & VN_data_in(11970);
  VN1995_in1 <= VN_sign_in(11971) & VN_data_in(11971);
  VN1995_in2 <= VN_sign_in(11972) & VN_data_in(11972);
  VN1995_in3 <= VN_sign_in(11973) & VN_data_in(11973);
  VN1995_in4 <= VN_sign_in(11974) & VN_data_in(11974);
  VN1995_in5 <= VN_sign_in(11975) & VN_data_in(11975);
  VN1996_in0 <= VN_sign_in(11976) & VN_data_in(11976);
  VN1996_in1 <= VN_sign_in(11977) & VN_data_in(11977);
  VN1996_in2 <= VN_sign_in(11978) & VN_data_in(11978);
  VN1996_in3 <= VN_sign_in(11979) & VN_data_in(11979);
  VN1996_in4 <= VN_sign_in(11980) & VN_data_in(11980);
  VN1996_in5 <= VN_sign_in(11981) & VN_data_in(11981);
  VN1997_in0 <= VN_sign_in(11982) & VN_data_in(11982);
  VN1997_in1 <= VN_sign_in(11983) & VN_data_in(11983);
  VN1997_in2 <= VN_sign_in(11984) & VN_data_in(11984);
  VN1997_in3 <= VN_sign_in(11985) & VN_data_in(11985);
  VN1997_in4 <= VN_sign_in(11986) & VN_data_in(11986);
  VN1997_in5 <= VN_sign_in(11987) & VN_data_in(11987);
  VN1998_in0 <= VN_sign_in(11988) & VN_data_in(11988);
  VN1998_in1 <= VN_sign_in(11989) & VN_data_in(11989);
  VN1998_in2 <= VN_sign_in(11990) & VN_data_in(11990);
  VN1998_in3 <= VN_sign_in(11991) & VN_data_in(11991);
  VN1998_in4 <= VN_sign_in(11992) & VN_data_in(11992);
  VN1998_in5 <= VN_sign_in(11993) & VN_data_in(11993);
  VN1999_in0 <= VN_sign_in(11994) & VN_data_in(11994);
  VN1999_in1 <= VN_sign_in(11995) & VN_data_in(11995);
  VN1999_in2 <= VN_sign_in(11996) & VN_data_in(11996);
  VN1999_in3 <= VN_sign_in(11997) & VN_data_in(11997);
  VN1999_in4 <= VN_sign_in(11998) & VN_data_in(11998);
  VN1999_in5 <= VN_sign_in(11999) & VN_data_in(11999);
  VN2000_in0 <= VN_sign_in(12000) & VN_data_in(12000);
  VN2000_in1 <= VN_sign_in(12001) & VN_data_in(12001);
  VN2000_in2 <= VN_sign_in(12002) & VN_data_in(12002);
  VN2000_in3 <= VN_sign_in(12003) & VN_data_in(12003);
  VN2000_in4 <= VN_sign_in(12004) & VN_data_in(12004);
  VN2000_in5 <= VN_sign_in(12005) & VN_data_in(12005);
  VN2001_in0 <= VN_sign_in(12006) & VN_data_in(12006);
  VN2001_in1 <= VN_sign_in(12007) & VN_data_in(12007);
  VN2001_in2 <= VN_sign_in(12008) & VN_data_in(12008);
  VN2001_in3 <= VN_sign_in(12009) & VN_data_in(12009);
  VN2001_in4 <= VN_sign_in(12010) & VN_data_in(12010);
  VN2001_in5 <= VN_sign_in(12011) & VN_data_in(12011);
  VN2002_in0 <= VN_sign_in(12012) & VN_data_in(12012);
  VN2002_in1 <= VN_sign_in(12013) & VN_data_in(12013);
  VN2002_in2 <= VN_sign_in(12014) & VN_data_in(12014);
  VN2002_in3 <= VN_sign_in(12015) & VN_data_in(12015);
  VN2002_in4 <= VN_sign_in(12016) & VN_data_in(12016);
  VN2002_in5 <= VN_sign_in(12017) & VN_data_in(12017);
  VN2003_in0 <= VN_sign_in(12018) & VN_data_in(12018);
  VN2003_in1 <= VN_sign_in(12019) & VN_data_in(12019);
  VN2003_in2 <= VN_sign_in(12020) & VN_data_in(12020);
  VN2003_in3 <= VN_sign_in(12021) & VN_data_in(12021);
  VN2003_in4 <= VN_sign_in(12022) & VN_data_in(12022);
  VN2003_in5 <= VN_sign_in(12023) & VN_data_in(12023);
  VN2004_in0 <= VN_sign_in(12024) & VN_data_in(12024);
  VN2004_in1 <= VN_sign_in(12025) & VN_data_in(12025);
  VN2004_in2 <= VN_sign_in(12026) & VN_data_in(12026);
  VN2004_in3 <= VN_sign_in(12027) & VN_data_in(12027);
  VN2004_in4 <= VN_sign_in(12028) & VN_data_in(12028);
  VN2004_in5 <= VN_sign_in(12029) & VN_data_in(12029);
  VN2005_in0 <= VN_sign_in(12030) & VN_data_in(12030);
  VN2005_in1 <= VN_sign_in(12031) & VN_data_in(12031);
  VN2005_in2 <= VN_sign_in(12032) & VN_data_in(12032);
  VN2005_in3 <= VN_sign_in(12033) & VN_data_in(12033);
  VN2005_in4 <= VN_sign_in(12034) & VN_data_in(12034);
  VN2005_in5 <= VN_sign_in(12035) & VN_data_in(12035);
  VN2006_in0 <= VN_sign_in(12036) & VN_data_in(12036);
  VN2006_in1 <= VN_sign_in(12037) & VN_data_in(12037);
  VN2006_in2 <= VN_sign_in(12038) & VN_data_in(12038);
  VN2006_in3 <= VN_sign_in(12039) & VN_data_in(12039);
  VN2006_in4 <= VN_sign_in(12040) & VN_data_in(12040);
  VN2006_in5 <= VN_sign_in(12041) & VN_data_in(12041);
  VN2007_in0 <= VN_sign_in(12042) & VN_data_in(12042);
  VN2007_in1 <= VN_sign_in(12043) & VN_data_in(12043);
  VN2007_in2 <= VN_sign_in(12044) & VN_data_in(12044);
  VN2007_in3 <= VN_sign_in(12045) & VN_data_in(12045);
  VN2007_in4 <= VN_sign_in(12046) & VN_data_in(12046);
  VN2007_in5 <= VN_sign_in(12047) & VN_data_in(12047);
  VN2008_in0 <= VN_sign_in(12048) & VN_data_in(12048);
  VN2008_in1 <= VN_sign_in(12049) & VN_data_in(12049);
  VN2008_in2 <= VN_sign_in(12050) & VN_data_in(12050);
  VN2008_in3 <= VN_sign_in(12051) & VN_data_in(12051);
  VN2008_in4 <= VN_sign_in(12052) & VN_data_in(12052);
  VN2008_in5 <= VN_sign_in(12053) & VN_data_in(12053);
  VN2009_in0 <= VN_sign_in(12054) & VN_data_in(12054);
  VN2009_in1 <= VN_sign_in(12055) & VN_data_in(12055);
  VN2009_in2 <= VN_sign_in(12056) & VN_data_in(12056);
  VN2009_in3 <= VN_sign_in(12057) & VN_data_in(12057);
  VN2009_in4 <= VN_sign_in(12058) & VN_data_in(12058);
  VN2009_in5 <= VN_sign_in(12059) & VN_data_in(12059);
  VN2010_in0 <= VN_sign_in(12060) & VN_data_in(12060);
  VN2010_in1 <= VN_sign_in(12061) & VN_data_in(12061);
  VN2010_in2 <= VN_sign_in(12062) & VN_data_in(12062);
  VN2010_in3 <= VN_sign_in(12063) & VN_data_in(12063);
  VN2010_in4 <= VN_sign_in(12064) & VN_data_in(12064);
  VN2010_in5 <= VN_sign_in(12065) & VN_data_in(12065);
  VN2011_in0 <= VN_sign_in(12066) & VN_data_in(12066);
  VN2011_in1 <= VN_sign_in(12067) & VN_data_in(12067);
  VN2011_in2 <= VN_sign_in(12068) & VN_data_in(12068);
  VN2011_in3 <= VN_sign_in(12069) & VN_data_in(12069);
  VN2011_in4 <= VN_sign_in(12070) & VN_data_in(12070);
  VN2011_in5 <= VN_sign_in(12071) & VN_data_in(12071);
  VN2012_in0 <= VN_sign_in(12072) & VN_data_in(12072);
  VN2012_in1 <= VN_sign_in(12073) & VN_data_in(12073);
  VN2012_in2 <= VN_sign_in(12074) & VN_data_in(12074);
  VN2012_in3 <= VN_sign_in(12075) & VN_data_in(12075);
  VN2012_in4 <= VN_sign_in(12076) & VN_data_in(12076);
  VN2012_in5 <= VN_sign_in(12077) & VN_data_in(12077);
  VN2013_in0 <= VN_sign_in(12078) & VN_data_in(12078);
  VN2013_in1 <= VN_sign_in(12079) & VN_data_in(12079);
  VN2013_in2 <= VN_sign_in(12080) & VN_data_in(12080);
  VN2013_in3 <= VN_sign_in(12081) & VN_data_in(12081);
  VN2013_in4 <= VN_sign_in(12082) & VN_data_in(12082);
  VN2013_in5 <= VN_sign_in(12083) & VN_data_in(12083);
  VN2014_in0 <= VN_sign_in(12084) & VN_data_in(12084);
  VN2014_in1 <= VN_sign_in(12085) & VN_data_in(12085);
  VN2014_in2 <= VN_sign_in(12086) & VN_data_in(12086);
  VN2014_in3 <= VN_sign_in(12087) & VN_data_in(12087);
  VN2014_in4 <= VN_sign_in(12088) & VN_data_in(12088);
  VN2014_in5 <= VN_sign_in(12089) & VN_data_in(12089);
  VN2015_in0 <= VN_sign_in(12090) & VN_data_in(12090);
  VN2015_in1 <= VN_sign_in(12091) & VN_data_in(12091);
  VN2015_in2 <= VN_sign_in(12092) & VN_data_in(12092);
  VN2015_in3 <= VN_sign_in(12093) & VN_data_in(12093);
  VN2015_in4 <= VN_sign_in(12094) & VN_data_in(12094);
  VN2015_in5 <= VN_sign_in(12095) & VN_data_in(12095);
  VN2016_in0 <= VN_sign_in(12096) & VN_data_in(12096);
  VN2016_in1 <= VN_sign_in(12097) & VN_data_in(12097);
  VN2016_in2 <= VN_sign_in(12098) & VN_data_in(12098);
  VN2016_in3 <= VN_sign_in(12099) & VN_data_in(12099);
  VN2016_in4 <= VN_sign_in(12100) & VN_data_in(12100);
  VN2016_in5 <= VN_sign_in(12101) & VN_data_in(12101);
  VN2017_in0 <= VN_sign_in(12102) & VN_data_in(12102);
  VN2017_in1 <= VN_sign_in(12103) & VN_data_in(12103);
  VN2017_in2 <= VN_sign_in(12104) & VN_data_in(12104);
  VN2017_in3 <= VN_sign_in(12105) & VN_data_in(12105);
  VN2017_in4 <= VN_sign_in(12106) & VN_data_in(12106);
  VN2017_in5 <= VN_sign_in(12107) & VN_data_in(12107);
  VN2018_in0 <= VN_sign_in(12108) & VN_data_in(12108);
  VN2018_in1 <= VN_sign_in(12109) & VN_data_in(12109);
  VN2018_in2 <= VN_sign_in(12110) & VN_data_in(12110);
  VN2018_in3 <= VN_sign_in(12111) & VN_data_in(12111);
  VN2018_in4 <= VN_sign_in(12112) & VN_data_in(12112);
  VN2018_in5 <= VN_sign_in(12113) & VN_data_in(12113);
  VN2019_in0 <= VN_sign_in(12114) & VN_data_in(12114);
  VN2019_in1 <= VN_sign_in(12115) & VN_data_in(12115);
  VN2019_in2 <= VN_sign_in(12116) & VN_data_in(12116);
  VN2019_in3 <= VN_sign_in(12117) & VN_data_in(12117);
  VN2019_in4 <= VN_sign_in(12118) & VN_data_in(12118);
  VN2019_in5 <= VN_sign_in(12119) & VN_data_in(12119);
  VN2020_in0 <= VN_sign_in(12120) & VN_data_in(12120);
  VN2020_in1 <= VN_sign_in(12121) & VN_data_in(12121);
  VN2020_in2 <= VN_sign_in(12122) & VN_data_in(12122);
  VN2020_in3 <= VN_sign_in(12123) & VN_data_in(12123);
  VN2020_in4 <= VN_sign_in(12124) & VN_data_in(12124);
  VN2020_in5 <= VN_sign_in(12125) & VN_data_in(12125);
  VN2021_in0 <= VN_sign_in(12126) & VN_data_in(12126);
  VN2021_in1 <= VN_sign_in(12127) & VN_data_in(12127);
  VN2021_in2 <= VN_sign_in(12128) & VN_data_in(12128);
  VN2021_in3 <= VN_sign_in(12129) & VN_data_in(12129);
  VN2021_in4 <= VN_sign_in(12130) & VN_data_in(12130);
  VN2021_in5 <= VN_sign_in(12131) & VN_data_in(12131);
  VN2022_in0 <= VN_sign_in(12132) & VN_data_in(12132);
  VN2022_in1 <= VN_sign_in(12133) & VN_data_in(12133);
  VN2022_in2 <= VN_sign_in(12134) & VN_data_in(12134);
  VN2022_in3 <= VN_sign_in(12135) & VN_data_in(12135);
  VN2022_in4 <= VN_sign_in(12136) & VN_data_in(12136);
  VN2022_in5 <= VN_sign_in(12137) & VN_data_in(12137);
  VN2023_in0 <= VN_sign_in(12138) & VN_data_in(12138);
  VN2023_in1 <= VN_sign_in(12139) & VN_data_in(12139);
  VN2023_in2 <= VN_sign_in(12140) & VN_data_in(12140);
  VN2023_in3 <= VN_sign_in(12141) & VN_data_in(12141);
  VN2023_in4 <= VN_sign_in(12142) & VN_data_in(12142);
  VN2023_in5 <= VN_sign_in(12143) & VN_data_in(12143);
  VN2024_in0 <= VN_sign_in(12144) & VN_data_in(12144);
  VN2024_in1 <= VN_sign_in(12145) & VN_data_in(12145);
  VN2024_in2 <= VN_sign_in(12146) & VN_data_in(12146);
  VN2024_in3 <= VN_sign_in(12147) & VN_data_in(12147);
  VN2024_in4 <= VN_sign_in(12148) & VN_data_in(12148);
  VN2024_in5 <= VN_sign_in(12149) & VN_data_in(12149);
  VN2025_in0 <= VN_sign_in(12150) & VN_data_in(12150);
  VN2025_in1 <= VN_sign_in(12151) & VN_data_in(12151);
  VN2025_in2 <= VN_sign_in(12152) & VN_data_in(12152);
  VN2025_in3 <= VN_sign_in(12153) & VN_data_in(12153);
  VN2025_in4 <= VN_sign_in(12154) & VN_data_in(12154);
  VN2025_in5 <= VN_sign_in(12155) & VN_data_in(12155);
  VN2026_in0 <= VN_sign_in(12156) & VN_data_in(12156);
  VN2026_in1 <= VN_sign_in(12157) & VN_data_in(12157);
  VN2026_in2 <= VN_sign_in(12158) & VN_data_in(12158);
  VN2026_in3 <= VN_sign_in(12159) & VN_data_in(12159);
  VN2026_in4 <= VN_sign_in(12160) & VN_data_in(12160);
  VN2026_in5 <= VN_sign_in(12161) & VN_data_in(12161);
  VN2027_in0 <= VN_sign_in(12162) & VN_data_in(12162);
  VN2027_in1 <= VN_sign_in(12163) & VN_data_in(12163);
  VN2027_in2 <= VN_sign_in(12164) & VN_data_in(12164);
  VN2027_in3 <= VN_sign_in(12165) & VN_data_in(12165);
  VN2027_in4 <= VN_sign_in(12166) & VN_data_in(12166);
  VN2027_in5 <= VN_sign_in(12167) & VN_data_in(12167);
  VN2028_in0 <= VN_sign_in(12168) & VN_data_in(12168);
  VN2028_in1 <= VN_sign_in(12169) & VN_data_in(12169);
  VN2028_in2 <= VN_sign_in(12170) & VN_data_in(12170);
  VN2028_in3 <= VN_sign_in(12171) & VN_data_in(12171);
  VN2028_in4 <= VN_sign_in(12172) & VN_data_in(12172);
  VN2028_in5 <= VN_sign_in(12173) & VN_data_in(12173);
  VN2029_in0 <= VN_sign_in(12174) & VN_data_in(12174);
  VN2029_in1 <= VN_sign_in(12175) & VN_data_in(12175);
  VN2029_in2 <= VN_sign_in(12176) & VN_data_in(12176);
  VN2029_in3 <= VN_sign_in(12177) & VN_data_in(12177);
  VN2029_in4 <= VN_sign_in(12178) & VN_data_in(12178);
  VN2029_in5 <= VN_sign_in(12179) & VN_data_in(12179);
  VN2030_in0 <= VN_sign_in(12180) & VN_data_in(12180);
  VN2030_in1 <= VN_sign_in(12181) & VN_data_in(12181);
  VN2030_in2 <= VN_sign_in(12182) & VN_data_in(12182);
  VN2030_in3 <= VN_sign_in(12183) & VN_data_in(12183);
  VN2030_in4 <= VN_sign_in(12184) & VN_data_in(12184);
  VN2030_in5 <= VN_sign_in(12185) & VN_data_in(12185);
  VN2031_in0 <= VN_sign_in(12186) & VN_data_in(12186);
  VN2031_in1 <= VN_sign_in(12187) & VN_data_in(12187);
  VN2031_in2 <= VN_sign_in(12188) & VN_data_in(12188);
  VN2031_in3 <= VN_sign_in(12189) & VN_data_in(12189);
  VN2031_in4 <= VN_sign_in(12190) & VN_data_in(12190);
  VN2031_in5 <= VN_sign_in(12191) & VN_data_in(12191);
  VN2032_in0 <= VN_sign_in(12192) & VN_data_in(12192);
  VN2032_in1 <= VN_sign_in(12193) & VN_data_in(12193);
  VN2032_in2 <= VN_sign_in(12194) & VN_data_in(12194);
  VN2032_in3 <= VN_sign_in(12195) & VN_data_in(12195);
  VN2032_in4 <= VN_sign_in(12196) & VN_data_in(12196);
  VN2032_in5 <= VN_sign_in(12197) & VN_data_in(12197);
  VN2033_in0 <= VN_sign_in(12198) & VN_data_in(12198);
  VN2033_in1 <= VN_sign_in(12199) & VN_data_in(12199);
  VN2033_in2 <= VN_sign_in(12200) & VN_data_in(12200);
  VN2033_in3 <= VN_sign_in(12201) & VN_data_in(12201);
  VN2033_in4 <= VN_sign_in(12202) & VN_data_in(12202);
  VN2033_in5 <= VN_sign_in(12203) & VN_data_in(12203);
  VN2034_in0 <= VN_sign_in(12204) & VN_data_in(12204);
  VN2034_in1 <= VN_sign_in(12205) & VN_data_in(12205);
  VN2034_in2 <= VN_sign_in(12206) & VN_data_in(12206);
  VN2034_in3 <= VN_sign_in(12207) & VN_data_in(12207);
  VN2034_in4 <= VN_sign_in(12208) & VN_data_in(12208);
  VN2034_in5 <= VN_sign_in(12209) & VN_data_in(12209);
  VN2035_in0 <= VN_sign_in(12210) & VN_data_in(12210);
  VN2035_in1 <= VN_sign_in(12211) & VN_data_in(12211);
  VN2035_in2 <= VN_sign_in(12212) & VN_data_in(12212);
  VN2035_in3 <= VN_sign_in(12213) & VN_data_in(12213);
  VN2035_in4 <= VN_sign_in(12214) & VN_data_in(12214);
  VN2035_in5 <= VN_sign_in(12215) & VN_data_in(12215);
  VN2036_in0 <= VN_sign_in(12216) & VN_data_in(12216);
  VN2036_in1 <= VN_sign_in(12217) & VN_data_in(12217);
  VN2036_in2 <= VN_sign_in(12218) & VN_data_in(12218);
  VN2036_in3 <= VN_sign_in(12219) & VN_data_in(12219);
  VN2036_in4 <= VN_sign_in(12220) & VN_data_in(12220);
  VN2036_in5 <= VN_sign_in(12221) & VN_data_in(12221);
  VN2037_in0 <= VN_sign_in(12222) & VN_data_in(12222);
  VN2037_in1 <= VN_sign_in(12223) & VN_data_in(12223);
  VN2037_in2 <= VN_sign_in(12224) & VN_data_in(12224);
  VN2037_in3 <= VN_sign_in(12225) & VN_data_in(12225);
  VN2037_in4 <= VN_sign_in(12226) & VN_data_in(12226);
  VN2037_in5 <= VN_sign_in(12227) & VN_data_in(12227);
  VN2038_in0 <= VN_sign_in(12228) & VN_data_in(12228);
  VN2038_in1 <= VN_sign_in(12229) & VN_data_in(12229);
  VN2038_in2 <= VN_sign_in(12230) & VN_data_in(12230);
  VN2038_in3 <= VN_sign_in(12231) & VN_data_in(12231);
  VN2038_in4 <= VN_sign_in(12232) & VN_data_in(12232);
  VN2038_in5 <= VN_sign_in(12233) & VN_data_in(12233);
  VN2039_in0 <= VN_sign_in(12234) & VN_data_in(12234);
  VN2039_in1 <= VN_sign_in(12235) & VN_data_in(12235);
  VN2039_in2 <= VN_sign_in(12236) & VN_data_in(12236);
  VN2039_in3 <= VN_sign_in(12237) & VN_data_in(12237);
  VN2039_in4 <= VN_sign_in(12238) & VN_data_in(12238);
  VN2039_in5 <= VN_sign_in(12239) & VN_data_in(12239);
  VN2040_in0 <= VN_sign_in(12240) & VN_data_in(12240);
  VN2040_in1 <= VN_sign_in(12241) & VN_data_in(12241);
  VN2040_in2 <= VN_sign_in(12242) & VN_data_in(12242);
  VN2040_in3 <= VN_sign_in(12243) & VN_data_in(12243);
  VN2040_in4 <= VN_sign_in(12244) & VN_data_in(12244);
  VN2040_in5 <= VN_sign_in(12245) & VN_data_in(12245);
  VN2041_in0 <= VN_sign_in(12246) & VN_data_in(12246);
  VN2041_in1 <= VN_sign_in(12247) & VN_data_in(12247);
  VN2041_in2 <= VN_sign_in(12248) & VN_data_in(12248);
  VN2041_in3 <= VN_sign_in(12249) & VN_data_in(12249);
  VN2041_in4 <= VN_sign_in(12250) & VN_data_in(12250);
  VN2041_in5 <= VN_sign_in(12251) & VN_data_in(12251);
  VN2042_in0 <= VN_sign_in(12252) & VN_data_in(12252);
  VN2042_in1 <= VN_sign_in(12253) & VN_data_in(12253);
  VN2042_in2 <= VN_sign_in(12254) & VN_data_in(12254);
  VN2042_in3 <= VN_sign_in(12255) & VN_data_in(12255);
  VN2042_in4 <= VN_sign_in(12256) & VN_data_in(12256);
  VN2042_in5 <= VN_sign_in(12257) & VN_data_in(12257);
  VN2043_in0 <= VN_sign_in(12258) & VN_data_in(12258);
  VN2043_in1 <= VN_sign_in(12259) & VN_data_in(12259);
  VN2043_in2 <= VN_sign_in(12260) & VN_data_in(12260);
  VN2043_in3 <= VN_sign_in(12261) & VN_data_in(12261);
  VN2043_in4 <= VN_sign_in(12262) & VN_data_in(12262);
  VN2043_in5 <= VN_sign_in(12263) & VN_data_in(12263);
  VN2044_in0 <= VN_sign_in(12264) & VN_data_in(12264);
  VN2044_in1 <= VN_sign_in(12265) & VN_data_in(12265);
  VN2044_in2 <= VN_sign_in(12266) & VN_data_in(12266);
  VN2044_in3 <= VN_sign_in(12267) & VN_data_in(12267);
  VN2044_in4 <= VN_sign_in(12268) & VN_data_in(12268);
  VN2044_in5 <= VN_sign_in(12269) & VN_data_in(12269);
  VN2045_in0 <= VN_sign_in(12270) & VN_data_in(12270);
  VN2045_in1 <= VN_sign_in(12271) & VN_data_in(12271);
  VN2045_in2 <= VN_sign_in(12272) & VN_data_in(12272);
  VN2045_in3 <= VN_sign_in(12273) & VN_data_in(12273);
  VN2045_in4 <= VN_sign_in(12274) & VN_data_in(12274);
  VN2045_in5 <= VN_sign_in(12275) & VN_data_in(12275);
  VN2046_in0 <= VN_sign_in(12276) & VN_data_in(12276);
  VN2046_in1 <= VN_sign_in(12277) & VN_data_in(12277);
  VN2046_in2 <= VN_sign_in(12278) & VN_data_in(12278);
  VN2046_in3 <= VN_sign_in(12279) & VN_data_in(12279);
  VN2046_in4 <= VN_sign_in(12280) & VN_data_in(12280);
  VN2046_in5 <= VN_sign_in(12281) & VN_data_in(12281);
  VN2047_in0 <= VN_sign_in(12282) & VN_data_in(12282);
  VN2047_in1 <= VN_sign_in(12283) & VN_data_in(12283);
  VN2047_in2 <= VN_sign_in(12284) & VN_data_in(12284);
  VN2047_in3 <= VN_sign_in(12285) & VN_data_in(12285);
  VN2047_in4 <= VN_sign_in(12286) & VN_data_in(12286);
  VN2047_in5 <= VN_sign_in(12287) & VN_data_in(12287);


    --VN0 : VN_Dv6 port map(
    --    clk => clk,
    --    rst_n => rst_n,
    --    DV_in => DV_in,
    --    RandomNum => RandomNum,
    --    LLR(5 downto 0) => LLLR,
    --    VN0_in0 => Din0,
    --    VN0_in1 => Din1,
    --    VN0_in2 => Din2,
    --    VN0_in3 => Din3,
    --    VN0_in4 => Din4,
    --    VN0_in5 => Din5,
    --    VN_data_out(0) => VN2CN0_bit,
    --    VN_data_out(1) => VN2CN1_bit,
    --    VN_data_out(2) => VN2CN2_bit,
    --    VN_data_out(3) => VN2CN3_bit,
    --    VN_data_out(4) => VN2CN4_bit,
    --    VN_data_out(5) => VN2CN5_bit,
    --    VN_sign_out(0) => VN2CN0_sign,
    --    VN_sign_out(1) => VN2CN1_sign,
    --    VN_sign_out(2) => VN2CN2_sign,
    --    VN_sign_out(3) => VN2CN3_sign,
    --    VN_sign_out(4) => VN2CN4_sign,
    --    VN_sign_out(5) => VN2CN5_sign,
    --    codeword(0) => codeword,
    --    Iterations => Iterations,
    --    DV_out => DV_out
    --);

--end architecture; --arch

    VN0 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5 downto 0),
        Din0 => VN0_in0,
        Din1 => VN0_in1,
        Din2 => VN0_in2,
        Din3 => VN0_in3,
        Din4 => VN0_in4,
        Din5 => VN0_in5,
        VN2CN0_bit => VN_data_out(0),
        VN2CN1_bit => VN_data_out(1),
        VN2CN2_bit => VN_data_out(2),
        VN2CN3_bit => VN_data_out(3),
        VN2CN4_bit => VN_data_out(4),
        VN2CN5_bit => VN_data_out(5),
        VN2CN0_sign => VN_sign_out(0),
        VN2CN1_sign => VN_sign_out(1),
        VN2CN2_sign => VN_sign_out(2),
        VN2CN3_sign => VN_sign_out(3),
        VN2CN4_sign => VN_sign_out(4),
        VN2CN5_sign => VN_sign_out(5),
        codeword => codeword(0),
        Iterations => Iterations,
        DV_out => DV_out,
        DecodeState => DecodeState
    );
    VN1 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11 downto 6),
        Din0 => VN1_in0,
        Din1 => VN1_in1,
        Din2 => VN1_in2,
        Din3 => VN1_in3,
        Din4 => VN1_in4,
        Din5 => VN1_in5,
        VN2CN0_bit => VN_data_out(6),
        VN2CN1_bit => VN_data_out(7),
        VN2CN2_bit => VN_data_out(8),
        VN2CN3_bit => VN_data_out(9),
        VN2CN4_bit => VN_data_out(10),
        VN2CN5_bit => VN_data_out(11),
        VN2CN0_sign => VN_sign_out(6),
        VN2CN1_sign => VN_sign_out(7),
        VN2CN2_sign => VN_sign_out(8),
        VN2CN3_sign => VN_sign_out(9),
        VN2CN4_sign => VN_sign_out(10),
        VN2CN5_sign => VN_sign_out(11),
        codeword => codeword(1),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(17 downto 12),
        Din0 => VN2_in0,
        Din1 => VN2_in1,
        Din2 => VN2_in2,
        Din3 => VN2_in3,
        Din4 => VN2_in4,
        Din5 => VN2_in5,
        VN2CN0_bit => VN_data_out(12),
        VN2CN1_bit => VN_data_out(13),
        VN2CN2_bit => VN_data_out(14),
        VN2CN3_bit => VN_data_out(15),
        VN2CN4_bit => VN_data_out(16),
        VN2CN5_bit => VN_data_out(17),
        VN2CN0_sign => VN_sign_out(12),
        VN2CN1_sign => VN_sign_out(13),
        VN2CN2_sign => VN_sign_out(14),
        VN2CN3_sign => VN_sign_out(15),
        VN2CN4_sign => VN_sign_out(16),
        VN2CN5_sign => VN_sign_out(17),
        codeword => codeword(2),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN3 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(23 downto 18),
        Din0 => VN3_in0,
        Din1 => VN3_in1,
        Din2 => VN3_in2,
        Din3 => VN3_in3,
        Din4 => VN3_in4,
        Din5 => VN3_in5,
        VN2CN0_bit => VN_data_out(18),
        VN2CN1_bit => VN_data_out(19),
        VN2CN2_bit => VN_data_out(20),
        VN2CN3_bit => VN_data_out(21),
        VN2CN4_bit => VN_data_out(22),
        VN2CN5_bit => VN_data_out(23),
        VN2CN0_sign => VN_sign_out(18),
        VN2CN1_sign => VN_sign_out(19),
        VN2CN2_sign => VN_sign_out(20),
        VN2CN3_sign => VN_sign_out(21),
        VN2CN4_sign => VN_sign_out(22),
        VN2CN5_sign => VN_sign_out(23),
        codeword => codeword(3),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN4 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(29 downto 24),
        Din0 => VN4_in0,
        Din1 => VN4_in1,
        Din2 => VN4_in2,
        Din3 => VN4_in3,
        Din4 => VN4_in4,
        Din5 => VN4_in5,
        VN2CN0_bit => VN_data_out(24),
        VN2CN1_bit => VN_data_out(25),
        VN2CN2_bit => VN_data_out(26),
        VN2CN3_bit => VN_data_out(27),
        VN2CN4_bit => VN_data_out(28),
        VN2CN5_bit => VN_data_out(29),
        VN2CN0_sign => VN_sign_out(24),
        VN2CN1_sign => VN_sign_out(25),
        VN2CN2_sign => VN_sign_out(26),
        VN2CN3_sign => VN_sign_out(27),
        VN2CN4_sign => VN_sign_out(28),
        VN2CN5_sign => VN_sign_out(29),
        codeword => codeword(4),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN5 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(35 downto 30),
        Din0 => VN5_in0,
        Din1 => VN5_in1,
        Din2 => VN5_in2,
        Din3 => VN5_in3,
        Din4 => VN5_in4,
        Din5 => VN5_in5,
        VN2CN0_bit => VN_data_out(30),
        VN2CN1_bit => VN_data_out(31),
        VN2CN2_bit => VN_data_out(32),
        VN2CN3_bit => VN_data_out(33),
        VN2CN4_bit => VN_data_out(34),
        VN2CN5_bit => VN_data_out(35),
        VN2CN0_sign => VN_sign_out(30),
        VN2CN1_sign => VN_sign_out(31),
        VN2CN2_sign => VN_sign_out(32),
        VN2CN3_sign => VN_sign_out(33),
        VN2CN4_sign => VN_sign_out(34),
        VN2CN5_sign => VN_sign_out(35),
        codeword => codeword(5),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN6 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(41 downto 36),
        Din0 => VN6_in0,
        Din1 => VN6_in1,
        Din2 => VN6_in2,
        Din3 => VN6_in3,
        Din4 => VN6_in4,
        Din5 => VN6_in5,
        VN2CN0_bit => VN_data_out(36),
        VN2CN1_bit => VN_data_out(37),
        VN2CN2_bit => VN_data_out(38),
        VN2CN3_bit => VN_data_out(39),
        VN2CN4_bit => VN_data_out(40),
        VN2CN5_bit => VN_data_out(41),
        VN2CN0_sign => VN_sign_out(36),
        VN2CN1_sign => VN_sign_out(37),
        VN2CN2_sign => VN_sign_out(38),
        VN2CN3_sign => VN_sign_out(39),
        VN2CN4_sign => VN_sign_out(40),
        VN2CN5_sign => VN_sign_out(41),
        codeword => codeword(6),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN7 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(47 downto 42),
        Din0 => VN7_in0,
        Din1 => VN7_in1,
        Din2 => VN7_in2,
        Din3 => VN7_in3,
        Din4 => VN7_in4,
        Din5 => VN7_in5,
        VN2CN0_bit => VN_data_out(42),
        VN2CN1_bit => VN_data_out(43),
        VN2CN2_bit => VN_data_out(44),
        VN2CN3_bit => VN_data_out(45),
        VN2CN4_bit => VN_data_out(46),
        VN2CN5_bit => VN_data_out(47),
        VN2CN0_sign => VN_sign_out(42),
        VN2CN1_sign => VN_sign_out(43),
        VN2CN2_sign => VN_sign_out(44),
        VN2CN3_sign => VN_sign_out(45),
        VN2CN4_sign => VN_sign_out(46),
        VN2CN5_sign => VN_sign_out(47),
        codeword => codeword(7),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN8 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(53 downto 48),
        Din0 => VN8_in0,
        Din1 => VN8_in1,
        Din2 => VN8_in2,
        Din3 => VN8_in3,
        Din4 => VN8_in4,
        Din5 => VN8_in5,
        VN2CN0_bit => VN_data_out(48),
        VN2CN1_bit => VN_data_out(49),
        VN2CN2_bit => VN_data_out(50),
        VN2CN3_bit => VN_data_out(51),
        VN2CN4_bit => VN_data_out(52),
        VN2CN5_bit => VN_data_out(53),
        VN2CN0_sign => VN_sign_out(48),
        VN2CN1_sign => VN_sign_out(49),
        VN2CN2_sign => VN_sign_out(50),
        VN2CN3_sign => VN_sign_out(51),
        VN2CN4_sign => VN_sign_out(52),
        VN2CN5_sign => VN_sign_out(53),
        codeword => codeword(8),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN9 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(59 downto 54),
        Din0 => VN9_in0,
        Din1 => VN9_in1,
        Din2 => VN9_in2,
        Din3 => VN9_in3,
        Din4 => VN9_in4,
        Din5 => VN9_in5,
        VN2CN0_bit => VN_data_out(54),
        VN2CN1_bit => VN_data_out(55),
        VN2CN2_bit => VN_data_out(56),
        VN2CN3_bit => VN_data_out(57),
        VN2CN4_bit => VN_data_out(58),
        VN2CN5_bit => VN_data_out(59),
        VN2CN0_sign => VN_sign_out(54),
        VN2CN1_sign => VN_sign_out(55),
        VN2CN2_sign => VN_sign_out(56),
        VN2CN3_sign => VN_sign_out(57),
        VN2CN4_sign => VN_sign_out(58),
        VN2CN5_sign => VN_sign_out(59),
        codeword => codeword(9),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN10 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(65 downto 60),
        Din0 => VN10_in0,
        Din1 => VN10_in1,
        Din2 => VN10_in2,
        Din3 => VN10_in3,
        Din4 => VN10_in4,
        Din5 => VN10_in5,
        VN2CN0_bit => VN_data_out(60),
        VN2CN1_bit => VN_data_out(61),
        VN2CN2_bit => VN_data_out(62),
        VN2CN3_bit => VN_data_out(63),
        VN2CN4_bit => VN_data_out(64),
        VN2CN5_bit => VN_data_out(65),
        VN2CN0_sign => VN_sign_out(60),
        VN2CN1_sign => VN_sign_out(61),
        VN2CN2_sign => VN_sign_out(62),
        VN2CN3_sign => VN_sign_out(63),
        VN2CN4_sign => VN_sign_out(64),
        VN2CN5_sign => VN_sign_out(65),
        codeword => codeword(10),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN11 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(71 downto 66),
        Din0 => VN11_in0,
        Din1 => VN11_in1,
        Din2 => VN11_in2,
        Din3 => VN11_in3,
        Din4 => VN11_in4,
        Din5 => VN11_in5,
        VN2CN0_bit => VN_data_out(66),
        VN2CN1_bit => VN_data_out(67),
        VN2CN2_bit => VN_data_out(68),
        VN2CN3_bit => VN_data_out(69),
        VN2CN4_bit => VN_data_out(70),
        VN2CN5_bit => VN_data_out(71),
        VN2CN0_sign => VN_sign_out(66),
        VN2CN1_sign => VN_sign_out(67),
        VN2CN2_sign => VN_sign_out(68),
        VN2CN3_sign => VN_sign_out(69),
        VN2CN4_sign => VN_sign_out(70),
        VN2CN5_sign => VN_sign_out(71),
        codeword => codeword(11),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN12 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(77 downto 72),
        Din0 => VN12_in0,
        Din1 => VN12_in1,
        Din2 => VN12_in2,
        Din3 => VN12_in3,
        Din4 => VN12_in4,
        Din5 => VN12_in5,
        VN2CN0_bit => VN_data_out(72),
        VN2CN1_bit => VN_data_out(73),
        VN2CN2_bit => VN_data_out(74),
        VN2CN3_bit => VN_data_out(75),
        VN2CN4_bit => VN_data_out(76),
        VN2CN5_bit => VN_data_out(77),
        VN2CN0_sign => VN_sign_out(72),
        VN2CN1_sign => VN_sign_out(73),
        VN2CN2_sign => VN_sign_out(74),
        VN2CN3_sign => VN_sign_out(75),
        VN2CN4_sign => VN_sign_out(76),
        VN2CN5_sign => VN_sign_out(77),
        codeword => codeword(12),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN13 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(83 downto 78),
        Din0 => VN13_in0,
        Din1 => VN13_in1,
        Din2 => VN13_in2,
        Din3 => VN13_in3,
        Din4 => VN13_in4,
        Din5 => VN13_in5,
        VN2CN0_bit => VN_data_out(78),
        VN2CN1_bit => VN_data_out(79),
        VN2CN2_bit => VN_data_out(80),
        VN2CN3_bit => VN_data_out(81),
        VN2CN4_bit => VN_data_out(82),
        VN2CN5_bit => VN_data_out(83),
        VN2CN0_sign => VN_sign_out(78),
        VN2CN1_sign => VN_sign_out(79),
        VN2CN2_sign => VN_sign_out(80),
        VN2CN3_sign => VN_sign_out(81),
        VN2CN4_sign => VN_sign_out(82),
        VN2CN5_sign => VN_sign_out(83),
        codeword => codeword(13),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN14 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(89 downto 84),
        Din0 => VN14_in0,
        Din1 => VN14_in1,
        Din2 => VN14_in2,
        Din3 => VN14_in3,
        Din4 => VN14_in4,
        Din5 => VN14_in5,
        VN2CN0_bit => VN_data_out(84),
        VN2CN1_bit => VN_data_out(85),
        VN2CN2_bit => VN_data_out(86),
        VN2CN3_bit => VN_data_out(87),
        VN2CN4_bit => VN_data_out(88),
        VN2CN5_bit => VN_data_out(89),
        VN2CN0_sign => VN_sign_out(84),
        VN2CN1_sign => VN_sign_out(85),
        VN2CN2_sign => VN_sign_out(86),
        VN2CN3_sign => VN_sign_out(87),
        VN2CN4_sign => VN_sign_out(88),
        VN2CN5_sign => VN_sign_out(89),
        codeword => codeword(14),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN15 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(95 downto 90),
        Din0 => VN15_in0,
        Din1 => VN15_in1,
        Din2 => VN15_in2,
        Din3 => VN15_in3,
        Din4 => VN15_in4,
        Din5 => VN15_in5,
        VN2CN0_bit => VN_data_out(90),
        VN2CN1_bit => VN_data_out(91),
        VN2CN2_bit => VN_data_out(92),
        VN2CN3_bit => VN_data_out(93),
        VN2CN4_bit => VN_data_out(94),
        VN2CN5_bit => VN_data_out(95),
        VN2CN0_sign => VN_sign_out(90),
        VN2CN1_sign => VN_sign_out(91),
        VN2CN2_sign => VN_sign_out(92),
        VN2CN3_sign => VN_sign_out(93),
        VN2CN4_sign => VN_sign_out(94),
        VN2CN5_sign => VN_sign_out(95),
        codeword => codeword(15),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN16 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(101 downto 96),
        Din0 => VN16_in0,
        Din1 => VN16_in1,
        Din2 => VN16_in2,
        Din3 => VN16_in3,
        Din4 => VN16_in4,
        Din5 => VN16_in5,
        VN2CN0_bit => VN_data_out(96),
        VN2CN1_bit => VN_data_out(97),
        VN2CN2_bit => VN_data_out(98),
        VN2CN3_bit => VN_data_out(99),
        VN2CN4_bit => VN_data_out(100),
        VN2CN5_bit => VN_data_out(101),
        VN2CN0_sign => VN_sign_out(96),
        VN2CN1_sign => VN_sign_out(97),
        VN2CN2_sign => VN_sign_out(98),
        VN2CN3_sign => VN_sign_out(99),
        VN2CN4_sign => VN_sign_out(100),
        VN2CN5_sign => VN_sign_out(101),
        codeword => codeword(16),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN17 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(107 downto 102),
        Din0 => VN17_in0,
        Din1 => VN17_in1,
        Din2 => VN17_in2,
        Din3 => VN17_in3,
        Din4 => VN17_in4,
        Din5 => VN17_in5,
        VN2CN0_bit => VN_data_out(102),
        VN2CN1_bit => VN_data_out(103),
        VN2CN2_bit => VN_data_out(104),
        VN2CN3_bit => VN_data_out(105),
        VN2CN4_bit => VN_data_out(106),
        VN2CN5_bit => VN_data_out(107),
        VN2CN0_sign => VN_sign_out(102),
        VN2CN1_sign => VN_sign_out(103),
        VN2CN2_sign => VN_sign_out(104),
        VN2CN3_sign => VN_sign_out(105),
        VN2CN4_sign => VN_sign_out(106),
        VN2CN5_sign => VN_sign_out(107),
        codeword => codeword(17),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN18 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(113 downto 108),
        Din0 => VN18_in0,
        Din1 => VN18_in1,
        Din2 => VN18_in2,
        Din3 => VN18_in3,
        Din4 => VN18_in4,
        Din5 => VN18_in5,
        VN2CN0_bit => VN_data_out(108),
        VN2CN1_bit => VN_data_out(109),
        VN2CN2_bit => VN_data_out(110),
        VN2CN3_bit => VN_data_out(111),
        VN2CN4_bit => VN_data_out(112),
        VN2CN5_bit => VN_data_out(113),
        VN2CN0_sign => VN_sign_out(108),
        VN2CN1_sign => VN_sign_out(109),
        VN2CN2_sign => VN_sign_out(110),
        VN2CN3_sign => VN_sign_out(111),
        VN2CN4_sign => VN_sign_out(112),
        VN2CN5_sign => VN_sign_out(113),
        codeword => codeword(18),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN19 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(119 downto 114),
        Din0 => VN19_in0,
        Din1 => VN19_in1,
        Din2 => VN19_in2,
        Din3 => VN19_in3,
        Din4 => VN19_in4,
        Din5 => VN19_in5,
        VN2CN0_bit => VN_data_out(114),
        VN2CN1_bit => VN_data_out(115),
        VN2CN2_bit => VN_data_out(116),
        VN2CN3_bit => VN_data_out(117),
        VN2CN4_bit => VN_data_out(118),
        VN2CN5_bit => VN_data_out(119),
        VN2CN0_sign => VN_sign_out(114),
        VN2CN1_sign => VN_sign_out(115),
        VN2CN2_sign => VN_sign_out(116),
        VN2CN3_sign => VN_sign_out(117),
        VN2CN4_sign => VN_sign_out(118),
        VN2CN5_sign => VN_sign_out(119),
        codeword => codeword(19),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN20 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(125 downto 120),
        Din0 => VN20_in0,
        Din1 => VN20_in1,
        Din2 => VN20_in2,
        Din3 => VN20_in3,
        Din4 => VN20_in4,
        Din5 => VN20_in5,
        VN2CN0_bit => VN_data_out(120),
        VN2CN1_bit => VN_data_out(121),
        VN2CN2_bit => VN_data_out(122),
        VN2CN3_bit => VN_data_out(123),
        VN2CN4_bit => VN_data_out(124),
        VN2CN5_bit => VN_data_out(125),
        VN2CN0_sign => VN_sign_out(120),
        VN2CN1_sign => VN_sign_out(121),
        VN2CN2_sign => VN_sign_out(122),
        VN2CN3_sign => VN_sign_out(123),
        VN2CN4_sign => VN_sign_out(124),
        VN2CN5_sign => VN_sign_out(125),
        codeword => codeword(20),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN21 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(131 downto 126),
        Din0 => VN21_in0,
        Din1 => VN21_in1,
        Din2 => VN21_in2,
        Din3 => VN21_in3,
        Din4 => VN21_in4,
        Din5 => VN21_in5,
        VN2CN0_bit => VN_data_out(126),
        VN2CN1_bit => VN_data_out(127),
        VN2CN2_bit => VN_data_out(128),
        VN2CN3_bit => VN_data_out(129),
        VN2CN4_bit => VN_data_out(130),
        VN2CN5_bit => VN_data_out(131),
        VN2CN0_sign => VN_sign_out(126),
        VN2CN1_sign => VN_sign_out(127),
        VN2CN2_sign => VN_sign_out(128),
        VN2CN3_sign => VN_sign_out(129),
        VN2CN4_sign => VN_sign_out(130),
        VN2CN5_sign => VN_sign_out(131),
        codeword => codeword(21),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN22 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(137 downto 132),
        Din0 => VN22_in0,
        Din1 => VN22_in1,
        Din2 => VN22_in2,
        Din3 => VN22_in3,
        Din4 => VN22_in4,
        Din5 => VN22_in5,
        VN2CN0_bit => VN_data_out(132),
        VN2CN1_bit => VN_data_out(133),
        VN2CN2_bit => VN_data_out(134),
        VN2CN3_bit => VN_data_out(135),
        VN2CN4_bit => VN_data_out(136),
        VN2CN5_bit => VN_data_out(137),
        VN2CN0_sign => VN_sign_out(132),
        VN2CN1_sign => VN_sign_out(133),
        VN2CN2_sign => VN_sign_out(134),
        VN2CN3_sign => VN_sign_out(135),
        VN2CN4_sign => VN_sign_out(136),
        VN2CN5_sign => VN_sign_out(137),
        codeword => codeword(22),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN23 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(143 downto 138),
        Din0 => VN23_in0,
        Din1 => VN23_in1,
        Din2 => VN23_in2,
        Din3 => VN23_in3,
        Din4 => VN23_in4,
        Din5 => VN23_in5,
        VN2CN0_bit => VN_data_out(138),
        VN2CN1_bit => VN_data_out(139),
        VN2CN2_bit => VN_data_out(140),
        VN2CN3_bit => VN_data_out(141),
        VN2CN4_bit => VN_data_out(142),
        VN2CN5_bit => VN_data_out(143),
        VN2CN0_sign => VN_sign_out(138),
        VN2CN1_sign => VN_sign_out(139),
        VN2CN2_sign => VN_sign_out(140),
        VN2CN3_sign => VN_sign_out(141),
        VN2CN4_sign => VN_sign_out(142),
        VN2CN5_sign => VN_sign_out(143),
        codeword => codeword(23),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN24 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(149 downto 144),
        Din0 => VN24_in0,
        Din1 => VN24_in1,
        Din2 => VN24_in2,
        Din3 => VN24_in3,
        Din4 => VN24_in4,
        Din5 => VN24_in5,
        VN2CN0_bit => VN_data_out(144),
        VN2CN1_bit => VN_data_out(145),
        VN2CN2_bit => VN_data_out(146),
        VN2CN3_bit => VN_data_out(147),
        VN2CN4_bit => VN_data_out(148),
        VN2CN5_bit => VN_data_out(149),
        VN2CN0_sign => VN_sign_out(144),
        VN2CN1_sign => VN_sign_out(145),
        VN2CN2_sign => VN_sign_out(146),
        VN2CN3_sign => VN_sign_out(147),
        VN2CN4_sign => VN_sign_out(148),
        VN2CN5_sign => VN_sign_out(149),
        codeword => codeword(24),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN25 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(155 downto 150),
        Din0 => VN25_in0,
        Din1 => VN25_in1,
        Din2 => VN25_in2,
        Din3 => VN25_in3,
        Din4 => VN25_in4,
        Din5 => VN25_in5,
        VN2CN0_bit => VN_data_out(150),
        VN2CN1_bit => VN_data_out(151),
        VN2CN2_bit => VN_data_out(152),
        VN2CN3_bit => VN_data_out(153),
        VN2CN4_bit => VN_data_out(154),
        VN2CN5_bit => VN_data_out(155),
        VN2CN0_sign => VN_sign_out(150),
        VN2CN1_sign => VN_sign_out(151),
        VN2CN2_sign => VN_sign_out(152),
        VN2CN3_sign => VN_sign_out(153),
        VN2CN4_sign => VN_sign_out(154),
        VN2CN5_sign => VN_sign_out(155),
        codeword => codeword(25),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN26 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(161 downto 156),
        Din0 => VN26_in0,
        Din1 => VN26_in1,
        Din2 => VN26_in2,
        Din3 => VN26_in3,
        Din4 => VN26_in4,
        Din5 => VN26_in5,
        VN2CN0_bit => VN_data_out(156),
        VN2CN1_bit => VN_data_out(157),
        VN2CN2_bit => VN_data_out(158),
        VN2CN3_bit => VN_data_out(159),
        VN2CN4_bit => VN_data_out(160),
        VN2CN5_bit => VN_data_out(161),
        VN2CN0_sign => VN_sign_out(156),
        VN2CN1_sign => VN_sign_out(157),
        VN2CN2_sign => VN_sign_out(158),
        VN2CN3_sign => VN_sign_out(159),
        VN2CN4_sign => VN_sign_out(160),
        VN2CN5_sign => VN_sign_out(161),
        codeword => codeword(26),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN27 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(167 downto 162),
        Din0 => VN27_in0,
        Din1 => VN27_in1,
        Din2 => VN27_in2,
        Din3 => VN27_in3,
        Din4 => VN27_in4,
        Din5 => VN27_in5,
        VN2CN0_bit => VN_data_out(162),
        VN2CN1_bit => VN_data_out(163),
        VN2CN2_bit => VN_data_out(164),
        VN2CN3_bit => VN_data_out(165),
        VN2CN4_bit => VN_data_out(166),
        VN2CN5_bit => VN_data_out(167),
        VN2CN0_sign => VN_sign_out(162),
        VN2CN1_sign => VN_sign_out(163),
        VN2CN2_sign => VN_sign_out(164),
        VN2CN3_sign => VN_sign_out(165),
        VN2CN4_sign => VN_sign_out(166),
        VN2CN5_sign => VN_sign_out(167),
        codeword => codeword(27),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN28 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(173 downto 168),
        Din0 => VN28_in0,
        Din1 => VN28_in1,
        Din2 => VN28_in2,
        Din3 => VN28_in3,
        Din4 => VN28_in4,
        Din5 => VN28_in5,
        VN2CN0_bit => VN_data_out(168),
        VN2CN1_bit => VN_data_out(169),
        VN2CN2_bit => VN_data_out(170),
        VN2CN3_bit => VN_data_out(171),
        VN2CN4_bit => VN_data_out(172),
        VN2CN5_bit => VN_data_out(173),
        VN2CN0_sign => VN_sign_out(168),
        VN2CN1_sign => VN_sign_out(169),
        VN2CN2_sign => VN_sign_out(170),
        VN2CN3_sign => VN_sign_out(171),
        VN2CN4_sign => VN_sign_out(172),
        VN2CN5_sign => VN_sign_out(173),
        codeword => codeword(28),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN29 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(179 downto 174),
        Din0 => VN29_in0,
        Din1 => VN29_in1,
        Din2 => VN29_in2,
        Din3 => VN29_in3,
        Din4 => VN29_in4,
        Din5 => VN29_in5,
        VN2CN0_bit => VN_data_out(174),
        VN2CN1_bit => VN_data_out(175),
        VN2CN2_bit => VN_data_out(176),
        VN2CN3_bit => VN_data_out(177),
        VN2CN4_bit => VN_data_out(178),
        VN2CN5_bit => VN_data_out(179),
        VN2CN0_sign => VN_sign_out(174),
        VN2CN1_sign => VN_sign_out(175),
        VN2CN2_sign => VN_sign_out(176),
        VN2CN3_sign => VN_sign_out(177),
        VN2CN4_sign => VN_sign_out(178),
        VN2CN5_sign => VN_sign_out(179),
        codeword => codeword(29),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN30 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(185 downto 180),
        Din0 => VN30_in0,
        Din1 => VN30_in1,
        Din2 => VN30_in2,
        Din3 => VN30_in3,
        Din4 => VN30_in4,
        Din5 => VN30_in5,
        VN2CN0_bit => VN_data_out(180),
        VN2CN1_bit => VN_data_out(181),
        VN2CN2_bit => VN_data_out(182),
        VN2CN3_bit => VN_data_out(183),
        VN2CN4_bit => VN_data_out(184),
        VN2CN5_bit => VN_data_out(185),
        VN2CN0_sign => VN_sign_out(180),
        VN2CN1_sign => VN_sign_out(181),
        VN2CN2_sign => VN_sign_out(182),
        VN2CN3_sign => VN_sign_out(183),
        VN2CN4_sign => VN_sign_out(184),
        VN2CN5_sign => VN_sign_out(185),
        codeword => codeword(30),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN31 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(191 downto 186),
        Din0 => VN31_in0,
        Din1 => VN31_in1,
        Din2 => VN31_in2,
        Din3 => VN31_in3,
        Din4 => VN31_in4,
        Din5 => VN31_in5,
        VN2CN0_bit => VN_data_out(186),
        VN2CN1_bit => VN_data_out(187),
        VN2CN2_bit => VN_data_out(188),
        VN2CN3_bit => VN_data_out(189),
        VN2CN4_bit => VN_data_out(190),
        VN2CN5_bit => VN_data_out(191),
        VN2CN0_sign => VN_sign_out(186),
        VN2CN1_sign => VN_sign_out(187),
        VN2CN2_sign => VN_sign_out(188),
        VN2CN3_sign => VN_sign_out(189),
        VN2CN4_sign => VN_sign_out(190),
        VN2CN5_sign => VN_sign_out(191),
        codeword => codeword(31),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN32 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(197 downto 192),
        Din0 => VN32_in0,
        Din1 => VN32_in1,
        Din2 => VN32_in2,
        Din3 => VN32_in3,
        Din4 => VN32_in4,
        Din5 => VN32_in5,
        VN2CN0_bit => VN_data_out(192),
        VN2CN1_bit => VN_data_out(193),
        VN2CN2_bit => VN_data_out(194),
        VN2CN3_bit => VN_data_out(195),
        VN2CN4_bit => VN_data_out(196),
        VN2CN5_bit => VN_data_out(197),
        VN2CN0_sign => VN_sign_out(192),
        VN2CN1_sign => VN_sign_out(193),
        VN2CN2_sign => VN_sign_out(194),
        VN2CN3_sign => VN_sign_out(195),
        VN2CN4_sign => VN_sign_out(196),
        VN2CN5_sign => VN_sign_out(197),
        codeword => codeword(32),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN33 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(203 downto 198),
        Din0 => VN33_in0,
        Din1 => VN33_in1,
        Din2 => VN33_in2,
        Din3 => VN33_in3,
        Din4 => VN33_in4,
        Din5 => VN33_in5,
        VN2CN0_bit => VN_data_out(198),
        VN2CN1_bit => VN_data_out(199),
        VN2CN2_bit => VN_data_out(200),
        VN2CN3_bit => VN_data_out(201),
        VN2CN4_bit => VN_data_out(202),
        VN2CN5_bit => VN_data_out(203),
        VN2CN0_sign => VN_sign_out(198),
        VN2CN1_sign => VN_sign_out(199),
        VN2CN2_sign => VN_sign_out(200),
        VN2CN3_sign => VN_sign_out(201),
        VN2CN4_sign => VN_sign_out(202),
        VN2CN5_sign => VN_sign_out(203),
        codeword => codeword(33),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN34 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(209 downto 204),
        Din0 => VN34_in0,
        Din1 => VN34_in1,
        Din2 => VN34_in2,
        Din3 => VN34_in3,
        Din4 => VN34_in4,
        Din5 => VN34_in5,
        VN2CN0_bit => VN_data_out(204),
        VN2CN1_bit => VN_data_out(205),
        VN2CN2_bit => VN_data_out(206),
        VN2CN3_bit => VN_data_out(207),
        VN2CN4_bit => VN_data_out(208),
        VN2CN5_bit => VN_data_out(209),
        VN2CN0_sign => VN_sign_out(204),
        VN2CN1_sign => VN_sign_out(205),
        VN2CN2_sign => VN_sign_out(206),
        VN2CN3_sign => VN_sign_out(207),
        VN2CN4_sign => VN_sign_out(208),
        VN2CN5_sign => VN_sign_out(209),
        codeword => codeword(34),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN35 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(215 downto 210),
        Din0 => VN35_in0,
        Din1 => VN35_in1,
        Din2 => VN35_in2,
        Din3 => VN35_in3,
        Din4 => VN35_in4,
        Din5 => VN35_in5,
        VN2CN0_bit => VN_data_out(210),
        VN2CN1_bit => VN_data_out(211),
        VN2CN2_bit => VN_data_out(212),
        VN2CN3_bit => VN_data_out(213),
        VN2CN4_bit => VN_data_out(214),
        VN2CN5_bit => VN_data_out(215),
        VN2CN0_sign => VN_sign_out(210),
        VN2CN1_sign => VN_sign_out(211),
        VN2CN2_sign => VN_sign_out(212),
        VN2CN3_sign => VN_sign_out(213),
        VN2CN4_sign => VN_sign_out(214),
        VN2CN5_sign => VN_sign_out(215),
        codeword => codeword(35),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN36 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(221 downto 216),
        Din0 => VN36_in0,
        Din1 => VN36_in1,
        Din2 => VN36_in2,
        Din3 => VN36_in3,
        Din4 => VN36_in4,
        Din5 => VN36_in5,
        VN2CN0_bit => VN_data_out(216),
        VN2CN1_bit => VN_data_out(217),
        VN2CN2_bit => VN_data_out(218),
        VN2CN3_bit => VN_data_out(219),
        VN2CN4_bit => VN_data_out(220),
        VN2CN5_bit => VN_data_out(221),
        VN2CN0_sign => VN_sign_out(216),
        VN2CN1_sign => VN_sign_out(217),
        VN2CN2_sign => VN_sign_out(218),
        VN2CN3_sign => VN_sign_out(219),
        VN2CN4_sign => VN_sign_out(220),
        VN2CN5_sign => VN_sign_out(221),
        codeword => codeword(36),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN37 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(227 downto 222),
        Din0 => VN37_in0,
        Din1 => VN37_in1,
        Din2 => VN37_in2,
        Din3 => VN37_in3,
        Din4 => VN37_in4,
        Din5 => VN37_in5,
        VN2CN0_bit => VN_data_out(222),
        VN2CN1_bit => VN_data_out(223),
        VN2CN2_bit => VN_data_out(224),
        VN2CN3_bit => VN_data_out(225),
        VN2CN4_bit => VN_data_out(226),
        VN2CN5_bit => VN_data_out(227),
        VN2CN0_sign => VN_sign_out(222),
        VN2CN1_sign => VN_sign_out(223),
        VN2CN2_sign => VN_sign_out(224),
        VN2CN3_sign => VN_sign_out(225),
        VN2CN4_sign => VN_sign_out(226),
        VN2CN5_sign => VN_sign_out(227),
        codeword => codeword(37),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN38 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(233 downto 228),
        Din0 => VN38_in0,
        Din1 => VN38_in1,
        Din2 => VN38_in2,
        Din3 => VN38_in3,
        Din4 => VN38_in4,
        Din5 => VN38_in5,
        VN2CN0_bit => VN_data_out(228),
        VN2CN1_bit => VN_data_out(229),
        VN2CN2_bit => VN_data_out(230),
        VN2CN3_bit => VN_data_out(231),
        VN2CN4_bit => VN_data_out(232),
        VN2CN5_bit => VN_data_out(233),
        VN2CN0_sign => VN_sign_out(228),
        VN2CN1_sign => VN_sign_out(229),
        VN2CN2_sign => VN_sign_out(230),
        VN2CN3_sign => VN_sign_out(231),
        VN2CN4_sign => VN_sign_out(232),
        VN2CN5_sign => VN_sign_out(233),
        codeword => codeword(38),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN39 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(239 downto 234),
        Din0 => VN39_in0,
        Din1 => VN39_in1,
        Din2 => VN39_in2,
        Din3 => VN39_in3,
        Din4 => VN39_in4,
        Din5 => VN39_in5,
        VN2CN0_bit => VN_data_out(234),
        VN2CN1_bit => VN_data_out(235),
        VN2CN2_bit => VN_data_out(236),
        VN2CN3_bit => VN_data_out(237),
        VN2CN4_bit => VN_data_out(238),
        VN2CN5_bit => VN_data_out(239),
        VN2CN0_sign => VN_sign_out(234),
        VN2CN1_sign => VN_sign_out(235),
        VN2CN2_sign => VN_sign_out(236),
        VN2CN3_sign => VN_sign_out(237),
        VN2CN4_sign => VN_sign_out(238),
        VN2CN5_sign => VN_sign_out(239),
        codeword => codeword(39),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN40 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(245 downto 240),
        Din0 => VN40_in0,
        Din1 => VN40_in1,
        Din2 => VN40_in2,
        Din3 => VN40_in3,
        Din4 => VN40_in4,
        Din5 => VN40_in5,
        VN2CN0_bit => VN_data_out(240),
        VN2CN1_bit => VN_data_out(241),
        VN2CN2_bit => VN_data_out(242),
        VN2CN3_bit => VN_data_out(243),
        VN2CN4_bit => VN_data_out(244),
        VN2CN5_bit => VN_data_out(245),
        VN2CN0_sign => VN_sign_out(240),
        VN2CN1_sign => VN_sign_out(241),
        VN2CN2_sign => VN_sign_out(242),
        VN2CN3_sign => VN_sign_out(243),
        VN2CN4_sign => VN_sign_out(244),
        VN2CN5_sign => VN_sign_out(245),
        codeword => codeword(40),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN41 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(251 downto 246),
        Din0 => VN41_in0,
        Din1 => VN41_in1,
        Din2 => VN41_in2,
        Din3 => VN41_in3,
        Din4 => VN41_in4,
        Din5 => VN41_in5,
        VN2CN0_bit => VN_data_out(246),
        VN2CN1_bit => VN_data_out(247),
        VN2CN2_bit => VN_data_out(248),
        VN2CN3_bit => VN_data_out(249),
        VN2CN4_bit => VN_data_out(250),
        VN2CN5_bit => VN_data_out(251),
        VN2CN0_sign => VN_sign_out(246),
        VN2CN1_sign => VN_sign_out(247),
        VN2CN2_sign => VN_sign_out(248),
        VN2CN3_sign => VN_sign_out(249),
        VN2CN4_sign => VN_sign_out(250),
        VN2CN5_sign => VN_sign_out(251),
        codeword => codeword(41),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN42 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(257 downto 252),
        Din0 => VN42_in0,
        Din1 => VN42_in1,
        Din2 => VN42_in2,
        Din3 => VN42_in3,
        Din4 => VN42_in4,
        Din5 => VN42_in5,
        VN2CN0_bit => VN_data_out(252),
        VN2CN1_bit => VN_data_out(253),
        VN2CN2_bit => VN_data_out(254),
        VN2CN3_bit => VN_data_out(255),
        VN2CN4_bit => VN_data_out(256),
        VN2CN5_bit => VN_data_out(257),
        VN2CN0_sign => VN_sign_out(252),
        VN2CN1_sign => VN_sign_out(253),
        VN2CN2_sign => VN_sign_out(254),
        VN2CN3_sign => VN_sign_out(255),
        VN2CN4_sign => VN_sign_out(256),
        VN2CN5_sign => VN_sign_out(257),
        codeword => codeword(42),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN43 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(263 downto 258),
        Din0 => VN43_in0,
        Din1 => VN43_in1,
        Din2 => VN43_in2,
        Din3 => VN43_in3,
        Din4 => VN43_in4,
        Din5 => VN43_in5,
        VN2CN0_bit => VN_data_out(258),
        VN2CN1_bit => VN_data_out(259),
        VN2CN2_bit => VN_data_out(260),
        VN2CN3_bit => VN_data_out(261),
        VN2CN4_bit => VN_data_out(262),
        VN2CN5_bit => VN_data_out(263),
        VN2CN0_sign => VN_sign_out(258),
        VN2CN1_sign => VN_sign_out(259),
        VN2CN2_sign => VN_sign_out(260),
        VN2CN3_sign => VN_sign_out(261),
        VN2CN4_sign => VN_sign_out(262),
        VN2CN5_sign => VN_sign_out(263),
        codeword => codeword(43),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN44 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(269 downto 264),
        Din0 => VN44_in0,
        Din1 => VN44_in1,
        Din2 => VN44_in2,
        Din3 => VN44_in3,
        Din4 => VN44_in4,
        Din5 => VN44_in5,
        VN2CN0_bit => VN_data_out(264),
        VN2CN1_bit => VN_data_out(265),
        VN2CN2_bit => VN_data_out(266),
        VN2CN3_bit => VN_data_out(267),
        VN2CN4_bit => VN_data_out(268),
        VN2CN5_bit => VN_data_out(269),
        VN2CN0_sign => VN_sign_out(264),
        VN2CN1_sign => VN_sign_out(265),
        VN2CN2_sign => VN_sign_out(266),
        VN2CN3_sign => VN_sign_out(267),
        VN2CN4_sign => VN_sign_out(268),
        VN2CN5_sign => VN_sign_out(269),
        codeword => codeword(44),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN45 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(275 downto 270),
        Din0 => VN45_in0,
        Din1 => VN45_in1,
        Din2 => VN45_in2,
        Din3 => VN45_in3,
        Din4 => VN45_in4,
        Din5 => VN45_in5,
        VN2CN0_bit => VN_data_out(270),
        VN2CN1_bit => VN_data_out(271),
        VN2CN2_bit => VN_data_out(272),
        VN2CN3_bit => VN_data_out(273),
        VN2CN4_bit => VN_data_out(274),
        VN2CN5_bit => VN_data_out(275),
        VN2CN0_sign => VN_sign_out(270),
        VN2CN1_sign => VN_sign_out(271),
        VN2CN2_sign => VN_sign_out(272),
        VN2CN3_sign => VN_sign_out(273),
        VN2CN4_sign => VN_sign_out(274),
        VN2CN5_sign => VN_sign_out(275),
        codeword => codeword(45),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN46 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(281 downto 276),
        Din0 => VN46_in0,
        Din1 => VN46_in1,
        Din2 => VN46_in2,
        Din3 => VN46_in3,
        Din4 => VN46_in4,
        Din5 => VN46_in5,
        VN2CN0_bit => VN_data_out(276),
        VN2CN1_bit => VN_data_out(277),
        VN2CN2_bit => VN_data_out(278),
        VN2CN3_bit => VN_data_out(279),
        VN2CN4_bit => VN_data_out(280),
        VN2CN5_bit => VN_data_out(281),
        VN2CN0_sign => VN_sign_out(276),
        VN2CN1_sign => VN_sign_out(277),
        VN2CN2_sign => VN_sign_out(278),
        VN2CN3_sign => VN_sign_out(279),
        VN2CN4_sign => VN_sign_out(280),
        VN2CN5_sign => VN_sign_out(281),
        codeword => codeword(46),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN47 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(287 downto 282),
        Din0 => VN47_in0,
        Din1 => VN47_in1,
        Din2 => VN47_in2,
        Din3 => VN47_in3,
        Din4 => VN47_in4,
        Din5 => VN47_in5,
        VN2CN0_bit => VN_data_out(282),
        VN2CN1_bit => VN_data_out(283),
        VN2CN2_bit => VN_data_out(284),
        VN2CN3_bit => VN_data_out(285),
        VN2CN4_bit => VN_data_out(286),
        VN2CN5_bit => VN_data_out(287),
        VN2CN0_sign => VN_sign_out(282),
        VN2CN1_sign => VN_sign_out(283),
        VN2CN2_sign => VN_sign_out(284),
        VN2CN3_sign => VN_sign_out(285),
        VN2CN4_sign => VN_sign_out(286),
        VN2CN5_sign => VN_sign_out(287),
        codeword => codeword(47),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN48 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(293 downto 288),
        Din0 => VN48_in0,
        Din1 => VN48_in1,
        Din2 => VN48_in2,
        Din3 => VN48_in3,
        Din4 => VN48_in4,
        Din5 => VN48_in5,
        VN2CN0_bit => VN_data_out(288),
        VN2CN1_bit => VN_data_out(289),
        VN2CN2_bit => VN_data_out(290),
        VN2CN3_bit => VN_data_out(291),
        VN2CN4_bit => VN_data_out(292),
        VN2CN5_bit => VN_data_out(293),
        VN2CN0_sign => VN_sign_out(288),
        VN2CN1_sign => VN_sign_out(289),
        VN2CN2_sign => VN_sign_out(290),
        VN2CN3_sign => VN_sign_out(291),
        VN2CN4_sign => VN_sign_out(292),
        VN2CN5_sign => VN_sign_out(293),
        codeword => codeword(48),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN49 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(299 downto 294),
        Din0 => VN49_in0,
        Din1 => VN49_in1,
        Din2 => VN49_in2,
        Din3 => VN49_in3,
        Din4 => VN49_in4,
        Din5 => VN49_in5,
        VN2CN0_bit => VN_data_out(294),
        VN2CN1_bit => VN_data_out(295),
        VN2CN2_bit => VN_data_out(296),
        VN2CN3_bit => VN_data_out(297),
        VN2CN4_bit => VN_data_out(298),
        VN2CN5_bit => VN_data_out(299),
        VN2CN0_sign => VN_sign_out(294),
        VN2CN1_sign => VN_sign_out(295),
        VN2CN2_sign => VN_sign_out(296),
        VN2CN3_sign => VN_sign_out(297),
        VN2CN4_sign => VN_sign_out(298),
        VN2CN5_sign => VN_sign_out(299),
        codeword => codeword(49),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN50 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(305 downto 300),
        Din0 => VN50_in0,
        Din1 => VN50_in1,
        Din2 => VN50_in2,
        Din3 => VN50_in3,
        Din4 => VN50_in4,
        Din5 => VN50_in5,
        VN2CN0_bit => VN_data_out(300),
        VN2CN1_bit => VN_data_out(301),
        VN2CN2_bit => VN_data_out(302),
        VN2CN3_bit => VN_data_out(303),
        VN2CN4_bit => VN_data_out(304),
        VN2CN5_bit => VN_data_out(305),
        VN2CN0_sign => VN_sign_out(300),
        VN2CN1_sign => VN_sign_out(301),
        VN2CN2_sign => VN_sign_out(302),
        VN2CN3_sign => VN_sign_out(303),
        VN2CN4_sign => VN_sign_out(304),
        VN2CN5_sign => VN_sign_out(305),
        codeword => codeword(50),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN51 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(311 downto 306),
        Din0 => VN51_in0,
        Din1 => VN51_in1,
        Din2 => VN51_in2,
        Din3 => VN51_in3,
        Din4 => VN51_in4,
        Din5 => VN51_in5,
        VN2CN0_bit => VN_data_out(306),
        VN2CN1_bit => VN_data_out(307),
        VN2CN2_bit => VN_data_out(308),
        VN2CN3_bit => VN_data_out(309),
        VN2CN4_bit => VN_data_out(310),
        VN2CN5_bit => VN_data_out(311),
        VN2CN0_sign => VN_sign_out(306),
        VN2CN1_sign => VN_sign_out(307),
        VN2CN2_sign => VN_sign_out(308),
        VN2CN3_sign => VN_sign_out(309),
        VN2CN4_sign => VN_sign_out(310),
        VN2CN5_sign => VN_sign_out(311),
        codeword => codeword(51),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN52 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(317 downto 312),
        Din0 => VN52_in0,
        Din1 => VN52_in1,
        Din2 => VN52_in2,
        Din3 => VN52_in3,
        Din4 => VN52_in4,
        Din5 => VN52_in5,
        VN2CN0_bit => VN_data_out(312),
        VN2CN1_bit => VN_data_out(313),
        VN2CN2_bit => VN_data_out(314),
        VN2CN3_bit => VN_data_out(315),
        VN2CN4_bit => VN_data_out(316),
        VN2CN5_bit => VN_data_out(317),
        VN2CN0_sign => VN_sign_out(312),
        VN2CN1_sign => VN_sign_out(313),
        VN2CN2_sign => VN_sign_out(314),
        VN2CN3_sign => VN_sign_out(315),
        VN2CN4_sign => VN_sign_out(316),
        VN2CN5_sign => VN_sign_out(317),
        codeword => codeword(52),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN53 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(323 downto 318),
        Din0 => VN53_in0,
        Din1 => VN53_in1,
        Din2 => VN53_in2,
        Din3 => VN53_in3,
        Din4 => VN53_in4,
        Din5 => VN53_in5,
        VN2CN0_bit => VN_data_out(318),
        VN2CN1_bit => VN_data_out(319),
        VN2CN2_bit => VN_data_out(320),
        VN2CN3_bit => VN_data_out(321),
        VN2CN4_bit => VN_data_out(322),
        VN2CN5_bit => VN_data_out(323),
        VN2CN0_sign => VN_sign_out(318),
        VN2CN1_sign => VN_sign_out(319),
        VN2CN2_sign => VN_sign_out(320),
        VN2CN3_sign => VN_sign_out(321),
        VN2CN4_sign => VN_sign_out(322),
        VN2CN5_sign => VN_sign_out(323),
        codeword => codeword(53),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN54 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(329 downto 324),
        Din0 => VN54_in0,
        Din1 => VN54_in1,
        Din2 => VN54_in2,
        Din3 => VN54_in3,
        Din4 => VN54_in4,
        Din5 => VN54_in5,
        VN2CN0_bit => VN_data_out(324),
        VN2CN1_bit => VN_data_out(325),
        VN2CN2_bit => VN_data_out(326),
        VN2CN3_bit => VN_data_out(327),
        VN2CN4_bit => VN_data_out(328),
        VN2CN5_bit => VN_data_out(329),
        VN2CN0_sign => VN_sign_out(324),
        VN2CN1_sign => VN_sign_out(325),
        VN2CN2_sign => VN_sign_out(326),
        VN2CN3_sign => VN_sign_out(327),
        VN2CN4_sign => VN_sign_out(328),
        VN2CN5_sign => VN_sign_out(329),
        codeword => codeword(54),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN55 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(335 downto 330),
        Din0 => VN55_in0,
        Din1 => VN55_in1,
        Din2 => VN55_in2,
        Din3 => VN55_in3,
        Din4 => VN55_in4,
        Din5 => VN55_in5,
        VN2CN0_bit => VN_data_out(330),
        VN2CN1_bit => VN_data_out(331),
        VN2CN2_bit => VN_data_out(332),
        VN2CN3_bit => VN_data_out(333),
        VN2CN4_bit => VN_data_out(334),
        VN2CN5_bit => VN_data_out(335),
        VN2CN0_sign => VN_sign_out(330),
        VN2CN1_sign => VN_sign_out(331),
        VN2CN2_sign => VN_sign_out(332),
        VN2CN3_sign => VN_sign_out(333),
        VN2CN4_sign => VN_sign_out(334),
        VN2CN5_sign => VN_sign_out(335),
        codeword => codeword(55),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN56 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(341 downto 336),
        Din0 => VN56_in0,
        Din1 => VN56_in1,
        Din2 => VN56_in2,
        Din3 => VN56_in3,
        Din4 => VN56_in4,
        Din5 => VN56_in5,
        VN2CN0_bit => VN_data_out(336),
        VN2CN1_bit => VN_data_out(337),
        VN2CN2_bit => VN_data_out(338),
        VN2CN3_bit => VN_data_out(339),
        VN2CN4_bit => VN_data_out(340),
        VN2CN5_bit => VN_data_out(341),
        VN2CN0_sign => VN_sign_out(336),
        VN2CN1_sign => VN_sign_out(337),
        VN2CN2_sign => VN_sign_out(338),
        VN2CN3_sign => VN_sign_out(339),
        VN2CN4_sign => VN_sign_out(340),
        VN2CN5_sign => VN_sign_out(341),
        codeword => codeword(56),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN57 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(347 downto 342),
        Din0 => VN57_in0,
        Din1 => VN57_in1,
        Din2 => VN57_in2,
        Din3 => VN57_in3,
        Din4 => VN57_in4,
        Din5 => VN57_in5,
        VN2CN0_bit => VN_data_out(342),
        VN2CN1_bit => VN_data_out(343),
        VN2CN2_bit => VN_data_out(344),
        VN2CN3_bit => VN_data_out(345),
        VN2CN4_bit => VN_data_out(346),
        VN2CN5_bit => VN_data_out(347),
        VN2CN0_sign => VN_sign_out(342),
        VN2CN1_sign => VN_sign_out(343),
        VN2CN2_sign => VN_sign_out(344),
        VN2CN3_sign => VN_sign_out(345),
        VN2CN4_sign => VN_sign_out(346),
        VN2CN5_sign => VN_sign_out(347),
        codeword => codeword(57),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN58 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(353 downto 348),
        Din0 => VN58_in0,
        Din1 => VN58_in1,
        Din2 => VN58_in2,
        Din3 => VN58_in3,
        Din4 => VN58_in4,
        Din5 => VN58_in5,
        VN2CN0_bit => VN_data_out(348),
        VN2CN1_bit => VN_data_out(349),
        VN2CN2_bit => VN_data_out(350),
        VN2CN3_bit => VN_data_out(351),
        VN2CN4_bit => VN_data_out(352),
        VN2CN5_bit => VN_data_out(353),
        VN2CN0_sign => VN_sign_out(348),
        VN2CN1_sign => VN_sign_out(349),
        VN2CN2_sign => VN_sign_out(350),
        VN2CN3_sign => VN_sign_out(351),
        VN2CN4_sign => VN_sign_out(352),
        VN2CN5_sign => VN_sign_out(353),
        codeword => codeword(58),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN59 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(359 downto 354),
        Din0 => VN59_in0,
        Din1 => VN59_in1,
        Din2 => VN59_in2,
        Din3 => VN59_in3,
        Din4 => VN59_in4,
        Din5 => VN59_in5,
        VN2CN0_bit => VN_data_out(354),
        VN2CN1_bit => VN_data_out(355),
        VN2CN2_bit => VN_data_out(356),
        VN2CN3_bit => VN_data_out(357),
        VN2CN4_bit => VN_data_out(358),
        VN2CN5_bit => VN_data_out(359),
        VN2CN0_sign => VN_sign_out(354),
        VN2CN1_sign => VN_sign_out(355),
        VN2CN2_sign => VN_sign_out(356),
        VN2CN3_sign => VN_sign_out(357),
        VN2CN4_sign => VN_sign_out(358),
        VN2CN5_sign => VN_sign_out(359),
        codeword => codeword(59),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN60 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(365 downto 360),
        Din0 => VN60_in0,
        Din1 => VN60_in1,
        Din2 => VN60_in2,
        Din3 => VN60_in3,
        Din4 => VN60_in4,
        Din5 => VN60_in5,
        VN2CN0_bit => VN_data_out(360),
        VN2CN1_bit => VN_data_out(361),
        VN2CN2_bit => VN_data_out(362),
        VN2CN3_bit => VN_data_out(363),
        VN2CN4_bit => VN_data_out(364),
        VN2CN5_bit => VN_data_out(365),
        VN2CN0_sign => VN_sign_out(360),
        VN2CN1_sign => VN_sign_out(361),
        VN2CN2_sign => VN_sign_out(362),
        VN2CN3_sign => VN_sign_out(363),
        VN2CN4_sign => VN_sign_out(364),
        VN2CN5_sign => VN_sign_out(365),
        codeword => codeword(60),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN61 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(371 downto 366),
        Din0 => VN61_in0,
        Din1 => VN61_in1,
        Din2 => VN61_in2,
        Din3 => VN61_in3,
        Din4 => VN61_in4,
        Din5 => VN61_in5,
        VN2CN0_bit => VN_data_out(366),
        VN2CN1_bit => VN_data_out(367),
        VN2CN2_bit => VN_data_out(368),
        VN2CN3_bit => VN_data_out(369),
        VN2CN4_bit => VN_data_out(370),
        VN2CN5_bit => VN_data_out(371),
        VN2CN0_sign => VN_sign_out(366),
        VN2CN1_sign => VN_sign_out(367),
        VN2CN2_sign => VN_sign_out(368),
        VN2CN3_sign => VN_sign_out(369),
        VN2CN4_sign => VN_sign_out(370),
        VN2CN5_sign => VN_sign_out(371),
        codeword => codeword(61),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN62 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(377 downto 372),
        Din0 => VN62_in0,
        Din1 => VN62_in1,
        Din2 => VN62_in2,
        Din3 => VN62_in3,
        Din4 => VN62_in4,
        Din5 => VN62_in5,
        VN2CN0_bit => VN_data_out(372),
        VN2CN1_bit => VN_data_out(373),
        VN2CN2_bit => VN_data_out(374),
        VN2CN3_bit => VN_data_out(375),
        VN2CN4_bit => VN_data_out(376),
        VN2CN5_bit => VN_data_out(377),
        VN2CN0_sign => VN_sign_out(372),
        VN2CN1_sign => VN_sign_out(373),
        VN2CN2_sign => VN_sign_out(374),
        VN2CN3_sign => VN_sign_out(375),
        VN2CN4_sign => VN_sign_out(376),
        VN2CN5_sign => VN_sign_out(377),
        codeword => codeword(62),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN63 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(383 downto 378),
        Din0 => VN63_in0,
        Din1 => VN63_in1,
        Din2 => VN63_in2,
        Din3 => VN63_in3,
        Din4 => VN63_in4,
        Din5 => VN63_in5,
        VN2CN0_bit => VN_data_out(378),
        VN2CN1_bit => VN_data_out(379),
        VN2CN2_bit => VN_data_out(380),
        VN2CN3_bit => VN_data_out(381),
        VN2CN4_bit => VN_data_out(382),
        VN2CN5_bit => VN_data_out(383),
        VN2CN0_sign => VN_sign_out(378),
        VN2CN1_sign => VN_sign_out(379),
        VN2CN2_sign => VN_sign_out(380),
        VN2CN3_sign => VN_sign_out(381),
        VN2CN4_sign => VN_sign_out(382),
        VN2CN5_sign => VN_sign_out(383),
        codeword => codeword(63),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN64 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(389 downto 384),
        Din0 => VN64_in0,
        Din1 => VN64_in1,
        Din2 => VN64_in2,
        Din3 => VN64_in3,
        Din4 => VN64_in4,
        Din5 => VN64_in5,
        VN2CN0_bit => VN_data_out(384),
        VN2CN1_bit => VN_data_out(385),
        VN2CN2_bit => VN_data_out(386),
        VN2CN3_bit => VN_data_out(387),
        VN2CN4_bit => VN_data_out(388),
        VN2CN5_bit => VN_data_out(389),
        VN2CN0_sign => VN_sign_out(384),
        VN2CN1_sign => VN_sign_out(385),
        VN2CN2_sign => VN_sign_out(386),
        VN2CN3_sign => VN_sign_out(387),
        VN2CN4_sign => VN_sign_out(388),
        VN2CN5_sign => VN_sign_out(389),
        codeword => codeword(64),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN65 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(395 downto 390),
        Din0 => VN65_in0,
        Din1 => VN65_in1,
        Din2 => VN65_in2,
        Din3 => VN65_in3,
        Din4 => VN65_in4,
        Din5 => VN65_in5,
        VN2CN0_bit => VN_data_out(390),
        VN2CN1_bit => VN_data_out(391),
        VN2CN2_bit => VN_data_out(392),
        VN2CN3_bit => VN_data_out(393),
        VN2CN4_bit => VN_data_out(394),
        VN2CN5_bit => VN_data_out(395),
        VN2CN0_sign => VN_sign_out(390),
        VN2CN1_sign => VN_sign_out(391),
        VN2CN2_sign => VN_sign_out(392),
        VN2CN3_sign => VN_sign_out(393),
        VN2CN4_sign => VN_sign_out(394),
        VN2CN5_sign => VN_sign_out(395),
        codeword => codeword(65),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN66 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(401 downto 396),
        Din0 => VN66_in0,
        Din1 => VN66_in1,
        Din2 => VN66_in2,
        Din3 => VN66_in3,
        Din4 => VN66_in4,
        Din5 => VN66_in5,
        VN2CN0_bit => VN_data_out(396),
        VN2CN1_bit => VN_data_out(397),
        VN2CN2_bit => VN_data_out(398),
        VN2CN3_bit => VN_data_out(399),
        VN2CN4_bit => VN_data_out(400),
        VN2CN5_bit => VN_data_out(401),
        VN2CN0_sign => VN_sign_out(396),
        VN2CN1_sign => VN_sign_out(397),
        VN2CN2_sign => VN_sign_out(398),
        VN2CN3_sign => VN_sign_out(399),
        VN2CN4_sign => VN_sign_out(400),
        VN2CN5_sign => VN_sign_out(401),
        codeword => codeword(66),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN67 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(407 downto 402),
        Din0 => VN67_in0,
        Din1 => VN67_in1,
        Din2 => VN67_in2,
        Din3 => VN67_in3,
        Din4 => VN67_in4,
        Din5 => VN67_in5,
        VN2CN0_bit => VN_data_out(402),
        VN2CN1_bit => VN_data_out(403),
        VN2CN2_bit => VN_data_out(404),
        VN2CN3_bit => VN_data_out(405),
        VN2CN4_bit => VN_data_out(406),
        VN2CN5_bit => VN_data_out(407),
        VN2CN0_sign => VN_sign_out(402),
        VN2CN1_sign => VN_sign_out(403),
        VN2CN2_sign => VN_sign_out(404),
        VN2CN3_sign => VN_sign_out(405),
        VN2CN4_sign => VN_sign_out(406),
        VN2CN5_sign => VN_sign_out(407),
        codeword => codeword(67),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN68 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(413 downto 408),
        Din0 => VN68_in0,
        Din1 => VN68_in1,
        Din2 => VN68_in2,
        Din3 => VN68_in3,
        Din4 => VN68_in4,
        Din5 => VN68_in5,
        VN2CN0_bit => VN_data_out(408),
        VN2CN1_bit => VN_data_out(409),
        VN2CN2_bit => VN_data_out(410),
        VN2CN3_bit => VN_data_out(411),
        VN2CN4_bit => VN_data_out(412),
        VN2CN5_bit => VN_data_out(413),
        VN2CN0_sign => VN_sign_out(408),
        VN2CN1_sign => VN_sign_out(409),
        VN2CN2_sign => VN_sign_out(410),
        VN2CN3_sign => VN_sign_out(411),
        VN2CN4_sign => VN_sign_out(412),
        VN2CN5_sign => VN_sign_out(413),
        codeword => codeword(68),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN69 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(419 downto 414),
        Din0 => VN69_in0,
        Din1 => VN69_in1,
        Din2 => VN69_in2,
        Din3 => VN69_in3,
        Din4 => VN69_in4,
        Din5 => VN69_in5,
        VN2CN0_bit => VN_data_out(414),
        VN2CN1_bit => VN_data_out(415),
        VN2CN2_bit => VN_data_out(416),
        VN2CN3_bit => VN_data_out(417),
        VN2CN4_bit => VN_data_out(418),
        VN2CN5_bit => VN_data_out(419),
        VN2CN0_sign => VN_sign_out(414),
        VN2CN1_sign => VN_sign_out(415),
        VN2CN2_sign => VN_sign_out(416),
        VN2CN3_sign => VN_sign_out(417),
        VN2CN4_sign => VN_sign_out(418),
        VN2CN5_sign => VN_sign_out(419),
        codeword => codeword(69),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN70 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(425 downto 420),
        Din0 => VN70_in0,
        Din1 => VN70_in1,
        Din2 => VN70_in2,
        Din3 => VN70_in3,
        Din4 => VN70_in4,
        Din5 => VN70_in5,
        VN2CN0_bit => VN_data_out(420),
        VN2CN1_bit => VN_data_out(421),
        VN2CN2_bit => VN_data_out(422),
        VN2CN3_bit => VN_data_out(423),
        VN2CN4_bit => VN_data_out(424),
        VN2CN5_bit => VN_data_out(425),
        VN2CN0_sign => VN_sign_out(420),
        VN2CN1_sign => VN_sign_out(421),
        VN2CN2_sign => VN_sign_out(422),
        VN2CN3_sign => VN_sign_out(423),
        VN2CN4_sign => VN_sign_out(424),
        VN2CN5_sign => VN_sign_out(425),
        codeword => codeword(70),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN71 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(431 downto 426),
        Din0 => VN71_in0,
        Din1 => VN71_in1,
        Din2 => VN71_in2,
        Din3 => VN71_in3,
        Din4 => VN71_in4,
        Din5 => VN71_in5,
        VN2CN0_bit => VN_data_out(426),
        VN2CN1_bit => VN_data_out(427),
        VN2CN2_bit => VN_data_out(428),
        VN2CN3_bit => VN_data_out(429),
        VN2CN4_bit => VN_data_out(430),
        VN2CN5_bit => VN_data_out(431),
        VN2CN0_sign => VN_sign_out(426),
        VN2CN1_sign => VN_sign_out(427),
        VN2CN2_sign => VN_sign_out(428),
        VN2CN3_sign => VN_sign_out(429),
        VN2CN4_sign => VN_sign_out(430),
        VN2CN5_sign => VN_sign_out(431),
        codeword => codeword(71),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN72 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(437 downto 432),
        Din0 => VN72_in0,
        Din1 => VN72_in1,
        Din2 => VN72_in2,
        Din3 => VN72_in3,
        Din4 => VN72_in4,
        Din5 => VN72_in5,
        VN2CN0_bit => VN_data_out(432),
        VN2CN1_bit => VN_data_out(433),
        VN2CN2_bit => VN_data_out(434),
        VN2CN3_bit => VN_data_out(435),
        VN2CN4_bit => VN_data_out(436),
        VN2CN5_bit => VN_data_out(437),
        VN2CN0_sign => VN_sign_out(432),
        VN2CN1_sign => VN_sign_out(433),
        VN2CN2_sign => VN_sign_out(434),
        VN2CN3_sign => VN_sign_out(435),
        VN2CN4_sign => VN_sign_out(436),
        VN2CN5_sign => VN_sign_out(437),
        codeword => codeword(72),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN73 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(443 downto 438),
        Din0 => VN73_in0,
        Din1 => VN73_in1,
        Din2 => VN73_in2,
        Din3 => VN73_in3,
        Din4 => VN73_in4,
        Din5 => VN73_in5,
        VN2CN0_bit => VN_data_out(438),
        VN2CN1_bit => VN_data_out(439),
        VN2CN2_bit => VN_data_out(440),
        VN2CN3_bit => VN_data_out(441),
        VN2CN4_bit => VN_data_out(442),
        VN2CN5_bit => VN_data_out(443),
        VN2CN0_sign => VN_sign_out(438),
        VN2CN1_sign => VN_sign_out(439),
        VN2CN2_sign => VN_sign_out(440),
        VN2CN3_sign => VN_sign_out(441),
        VN2CN4_sign => VN_sign_out(442),
        VN2CN5_sign => VN_sign_out(443),
        codeword => codeword(73),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN74 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(449 downto 444),
        Din0 => VN74_in0,
        Din1 => VN74_in1,
        Din2 => VN74_in2,
        Din3 => VN74_in3,
        Din4 => VN74_in4,
        Din5 => VN74_in5,
        VN2CN0_bit => VN_data_out(444),
        VN2CN1_bit => VN_data_out(445),
        VN2CN2_bit => VN_data_out(446),
        VN2CN3_bit => VN_data_out(447),
        VN2CN4_bit => VN_data_out(448),
        VN2CN5_bit => VN_data_out(449),
        VN2CN0_sign => VN_sign_out(444),
        VN2CN1_sign => VN_sign_out(445),
        VN2CN2_sign => VN_sign_out(446),
        VN2CN3_sign => VN_sign_out(447),
        VN2CN4_sign => VN_sign_out(448),
        VN2CN5_sign => VN_sign_out(449),
        codeword => codeword(74),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN75 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(455 downto 450),
        Din0 => VN75_in0,
        Din1 => VN75_in1,
        Din2 => VN75_in2,
        Din3 => VN75_in3,
        Din4 => VN75_in4,
        Din5 => VN75_in5,
        VN2CN0_bit => VN_data_out(450),
        VN2CN1_bit => VN_data_out(451),
        VN2CN2_bit => VN_data_out(452),
        VN2CN3_bit => VN_data_out(453),
        VN2CN4_bit => VN_data_out(454),
        VN2CN5_bit => VN_data_out(455),
        VN2CN0_sign => VN_sign_out(450),
        VN2CN1_sign => VN_sign_out(451),
        VN2CN2_sign => VN_sign_out(452),
        VN2CN3_sign => VN_sign_out(453),
        VN2CN4_sign => VN_sign_out(454),
        VN2CN5_sign => VN_sign_out(455),
        codeword => codeword(75),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN76 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(461 downto 456),
        Din0 => VN76_in0,
        Din1 => VN76_in1,
        Din2 => VN76_in2,
        Din3 => VN76_in3,
        Din4 => VN76_in4,
        Din5 => VN76_in5,
        VN2CN0_bit => VN_data_out(456),
        VN2CN1_bit => VN_data_out(457),
        VN2CN2_bit => VN_data_out(458),
        VN2CN3_bit => VN_data_out(459),
        VN2CN4_bit => VN_data_out(460),
        VN2CN5_bit => VN_data_out(461),
        VN2CN0_sign => VN_sign_out(456),
        VN2CN1_sign => VN_sign_out(457),
        VN2CN2_sign => VN_sign_out(458),
        VN2CN3_sign => VN_sign_out(459),
        VN2CN4_sign => VN_sign_out(460),
        VN2CN5_sign => VN_sign_out(461),
        codeword => codeword(76),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN77 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(467 downto 462),
        Din0 => VN77_in0,
        Din1 => VN77_in1,
        Din2 => VN77_in2,
        Din3 => VN77_in3,
        Din4 => VN77_in4,
        Din5 => VN77_in5,
        VN2CN0_bit => VN_data_out(462),
        VN2CN1_bit => VN_data_out(463),
        VN2CN2_bit => VN_data_out(464),
        VN2CN3_bit => VN_data_out(465),
        VN2CN4_bit => VN_data_out(466),
        VN2CN5_bit => VN_data_out(467),
        VN2CN0_sign => VN_sign_out(462),
        VN2CN1_sign => VN_sign_out(463),
        VN2CN2_sign => VN_sign_out(464),
        VN2CN3_sign => VN_sign_out(465),
        VN2CN4_sign => VN_sign_out(466),
        VN2CN5_sign => VN_sign_out(467),
        codeword => codeword(77),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN78 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(473 downto 468),
        Din0 => VN78_in0,
        Din1 => VN78_in1,
        Din2 => VN78_in2,
        Din3 => VN78_in3,
        Din4 => VN78_in4,
        Din5 => VN78_in5,
        VN2CN0_bit => VN_data_out(468),
        VN2CN1_bit => VN_data_out(469),
        VN2CN2_bit => VN_data_out(470),
        VN2CN3_bit => VN_data_out(471),
        VN2CN4_bit => VN_data_out(472),
        VN2CN5_bit => VN_data_out(473),
        VN2CN0_sign => VN_sign_out(468),
        VN2CN1_sign => VN_sign_out(469),
        VN2CN2_sign => VN_sign_out(470),
        VN2CN3_sign => VN_sign_out(471),
        VN2CN4_sign => VN_sign_out(472),
        VN2CN5_sign => VN_sign_out(473),
        codeword => codeword(78),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN79 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(479 downto 474),
        Din0 => VN79_in0,
        Din1 => VN79_in1,
        Din2 => VN79_in2,
        Din3 => VN79_in3,
        Din4 => VN79_in4,
        Din5 => VN79_in5,
        VN2CN0_bit => VN_data_out(474),
        VN2CN1_bit => VN_data_out(475),
        VN2CN2_bit => VN_data_out(476),
        VN2CN3_bit => VN_data_out(477),
        VN2CN4_bit => VN_data_out(478),
        VN2CN5_bit => VN_data_out(479),
        VN2CN0_sign => VN_sign_out(474),
        VN2CN1_sign => VN_sign_out(475),
        VN2CN2_sign => VN_sign_out(476),
        VN2CN3_sign => VN_sign_out(477),
        VN2CN4_sign => VN_sign_out(478),
        VN2CN5_sign => VN_sign_out(479),
        codeword => codeword(79),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN80 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(485 downto 480),
        Din0 => VN80_in0,
        Din1 => VN80_in1,
        Din2 => VN80_in2,
        Din3 => VN80_in3,
        Din4 => VN80_in4,
        Din5 => VN80_in5,
        VN2CN0_bit => VN_data_out(480),
        VN2CN1_bit => VN_data_out(481),
        VN2CN2_bit => VN_data_out(482),
        VN2CN3_bit => VN_data_out(483),
        VN2CN4_bit => VN_data_out(484),
        VN2CN5_bit => VN_data_out(485),
        VN2CN0_sign => VN_sign_out(480),
        VN2CN1_sign => VN_sign_out(481),
        VN2CN2_sign => VN_sign_out(482),
        VN2CN3_sign => VN_sign_out(483),
        VN2CN4_sign => VN_sign_out(484),
        VN2CN5_sign => VN_sign_out(485),
        codeword => codeword(80),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN81 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(491 downto 486),
        Din0 => VN81_in0,
        Din1 => VN81_in1,
        Din2 => VN81_in2,
        Din3 => VN81_in3,
        Din4 => VN81_in4,
        Din5 => VN81_in5,
        VN2CN0_bit => VN_data_out(486),
        VN2CN1_bit => VN_data_out(487),
        VN2CN2_bit => VN_data_out(488),
        VN2CN3_bit => VN_data_out(489),
        VN2CN4_bit => VN_data_out(490),
        VN2CN5_bit => VN_data_out(491),
        VN2CN0_sign => VN_sign_out(486),
        VN2CN1_sign => VN_sign_out(487),
        VN2CN2_sign => VN_sign_out(488),
        VN2CN3_sign => VN_sign_out(489),
        VN2CN4_sign => VN_sign_out(490),
        VN2CN5_sign => VN_sign_out(491),
        codeword => codeword(81),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN82 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(497 downto 492),
        Din0 => VN82_in0,
        Din1 => VN82_in1,
        Din2 => VN82_in2,
        Din3 => VN82_in3,
        Din4 => VN82_in4,
        Din5 => VN82_in5,
        VN2CN0_bit => VN_data_out(492),
        VN2CN1_bit => VN_data_out(493),
        VN2CN2_bit => VN_data_out(494),
        VN2CN3_bit => VN_data_out(495),
        VN2CN4_bit => VN_data_out(496),
        VN2CN5_bit => VN_data_out(497),
        VN2CN0_sign => VN_sign_out(492),
        VN2CN1_sign => VN_sign_out(493),
        VN2CN2_sign => VN_sign_out(494),
        VN2CN3_sign => VN_sign_out(495),
        VN2CN4_sign => VN_sign_out(496),
        VN2CN5_sign => VN_sign_out(497),
        codeword => codeword(82),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN83 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(503 downto 498),
        Din0 => VN83_in0,
        Din1 => VN83_in1,
        Din2 => VN83_in2,
        Din3 => VN83_in3,
        Din4 => VN83_in4,
        Din5 => VN83_in5,
        VN2CN0_bit => VN_data_out(498),
        VN2CN1_bit => VN_data_out(499),
        VN2CN2_bit => VN_data_out(500),
        VN2CN3_bit => VN_data_out(501),
        VN2CN4_bit => VN_data_out(502),
        VN2CN5_bit => VN_data_out(503),
        VN2CN0_sign => VN_sign_out(498),
        VN2CN1_sign => VN_sign_out(499),
        VN2CN2_sign => VN_sign_out(500),
        VN2CN3_sign => VN_sign_out(501),
        VN2CN4_sign => VN_sign_out(502),
        VN2CN5_sign => VN_sign_out(503),
        codeword => codeword(83),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN84 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(509 downto 504),
        Din0 => VN84_in0,
        Din1 => VN84_in1,
        Din2 => VN84_in2,
        Din3 => VN84_in3,
        Din4 => VN84_in4,
        Din5 => VN84_in5,
        VN2CN0_bit => VN_data_out(504),
        VN2CN1_bit => VN_data_out(505),
        VN2CN2_bit => VN_data_out(506),
        VN2CN3_bit => VN_data_out(507),
        VN2CN4_bit => VN_data_out(508),
        VN2CN5_bit => VN_data_out(509),
        VN2CN0_sign => VN_sign_out(504),
        VN2CN1_sign => VN_sign_out(505),
        VN2CN2_sign => VN_sign_out(506),
        VN2CN3_sign => VN_sign_out(507),
        VN2CN4_sign => VN_sign_out(508),
        VN2CN5_sign => VN_sign_out(509),
        codeword => codeword(84),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN85 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(515 downto 510),
        Din0 => VN85_in0,
        Din1 => VN85_in1,
        Din2 => VN85_in2,
        Din3 => VN85_in3,
        Din4 => VN85_in4,
        Din5 => VN85_in5,
        VN2CN0_bit => VN_data_out(510),
        VN2CN1_bit => VN_data_out(511),
        VN2CN2_bit => VN_data_out(512),
        VN2CN3_bit => VN_data_out(513),
        VN2CN4_bit => VN_data_out(514),
        VN2CN5_bit => VN_data_out(515),
        VN2CN0_sign => VN_sign_out(510),
        VN2CN1_sign => VN_sign_out(511),
        VN2CN2_sign => VN_sign_out(512),
        VN2CN3_sign => VN_sign_out(513),
        VN2CN4_sign => VN_sign_out(514),
        VN2CN5_sign => VN_sign_out(515),
        codeword => codeword(85),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN86 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(521 downto 516),
        Din0 => VN86_in0,
        Din1 => VN86_in1,
        Din2 => VN86_in2,
        Din3 => VN86_in3,
        Din4 => VN86_in4,
        Din5 => VN86_in5,
        VN2CN0_bit => VN_data_out(516),
        VN2CN1_bit => VN_data_out(517),
        VN2CN2_bit => VN_data_out(518),
        VN2CN3_bit => VN_data_out(519),
        VN2CN4_bit => VN_data_out(520),
        VN2CN5_bit => VN_data_out(521),
        VN2CN0_sign => VN_sign_out(516),
        VN2CN1_sign => VN_sign_out(517),
        VN2CN2_sign => VN_sign_out(518),
        VN2CN3_sign => VN_sign_out(519),
        VN2CN4_sign => VN_sign_out(520),
        VN2CN5_sign => VN_sign_out(521),
        codeword => codeword(86),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN87 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(527 downto 522),
        Din0 => VN87_in0,
        Din1 => VN87_in1,
        Din2 => VN87_in2,
        Din3 => VN87_in3,
        Din4 => VN87_in4,
        Din5 => VN87_in5,
        VN2CN0_bit => VN_data_out(522),
        VN2CN1_bit => VN_data_out(523),
        VN2CN2_bit => VN_data_out(524),
        VN2CN3_bit => VN_data_out(525),
        VN2CN4_bit => VN_data_out(526),
        VN2CN5_bit => VN_data_out(527),
        VN2CN0_sign => VN_sign_out(522),
        VN2CN1_sign => VN_sign_out(523),
        VN2CN2_sign => VN_sign_out(524),
        VN2CN3_sign => VN_sign_out(525),
        VN2CN4_sign => VN_sign_out(526),
        VN2CN5_sign => VN_sign_out(527),
        codeword => codeword(87),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN88 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(533 downto 528),
        Din0 => VN88_in0,
        Din1 => VN88_in1,
        Din2 => VN88_in2,
        Din3 => VN88_in3,
        Din4 => VN88_in4,
        Din5 => VN88_in5,
        VN2CN0_bit => VN_data_out(528),
        VN2CN1_bit => VN_data_out(529),
        VN2CN2_bit => VN_data_out(530),
        VN2CN3_bit => VN_data_out(531),
        VN2CN4_bit => VN_data_out(532),
        VN2CN5_bit => VN_data_out(533),
        VN2CN0_sign => VN_sign_out(528),
        VN2CN1_sign => VN_sign_out(529),
        VN2CN2_sign => VN_sign_out(530),
        VN2CN3_sign => VN_sign_out(531),
        VN2CN4_sign => VN_sign_out(532),
        VN2CN5_sign => VN_sign_out(533),
        codeword => codeword(88),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN89 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(539 downto 534),
        Din0 => VN89_in0,
        Din1 => VN89_in1,
        Din2 => VN89_in2,
        Din3 => VN89_in3,
        Din4 => VN89_in4,
        Din5 => VN89_in5,
        VN2CN0_bit => VN_data_out(534),
        VN2CN1_bit => VN_data_out(535),
        VN2CN2_bit => VN_data_out(536),
        VN2CN3_bit => VN_data_out(537),
        VN2CN4_bit => VN_data_out(538),
        VN2CN5_bit => VN_data_out(539),
        VN2CN0_sign => VN_sign_out(534),
        VN2CN1_sign => VN_sign_out(535),
        VN2CN2_sign => VN_sign_out(536),
        VN2CN3_sign => VN_sign_out(537),
        VN2CN4_sign => VN_sign_out(538),
        VN2CN5_sign => VN_sign_out(539),
        codeword => codeword(89),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN90 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(545 downto 540),
        Din0 => VN90_in0,
        Din1 => VN90_in1,
        Din2 => VN90_in2,
        Din3 => VN90_in3,
        Din4 => VN90_in4,
        Din5 => VN90_in5,
        VN2CN0_bit => VN_data_out(540),
        VN2CN1_bit => VN_data_out(541),
        VN2CN2_bit => VN_data_out(542),
        VN2CN3_bit => VN_data_out(543),
        VN2CN4_bit => VN_data_out(544),
        VN2CN5_bit => VN_data_out(545),
        VN2CN0_sign => VN_sign_out(540),
        VN2CN1_sign => VN_sign_out(541),
        VN2CN2_sign => VN_sign_out(542),
        VN2CN3_sign => VN_sign_out(543),
        VN2CN4_sign => VN_sign_out(544),
        VN2CN5_sign => VN_sign_out(545),
        codeword => codeword(90),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN91 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(551 downto 546),
        Din0 => VN91_in0,
        Din1 => VN91_in1,
        Din2 => VN91_in2,
        Din3 => VN91_in3,
        Din4 => VN91_in4,
        Din5 => VN91_in5,
        VN2CN0_bit => VN_data_out(546),
        VN2CN1_bit => VN_data_out(547),
        VN2CN2_bit => VN_data_out(548),
        VN2CN3_bit => VN_data_out(549),
        VN2CN4_bit => VN_data_out(550),
        VN2CN5_bit => VN_data_out(551),
        VN2CN0_sign => VN_sign_out(546),
        VN2CN1_sign => VN_sign_out(547),
        VN2CN2_sign => VN_sign_out(548),
        VN2CN3_sign => VN_sign_out(549),
        VN2CN4_sign => VN_sign_out(550),
        VN2CN5_sign => VN_sign_out(551),
        codeword => codeword(91),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN92 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(557 downto 552),
        Din0 => VN92_in0,
        Din1 => VN92_in1,
        Din2 => VN92_in2,
        Din3 => VN92_in3,
        Din4 => VN92_in4,
        Din5 => VN92_in5,
        VN2CN0_bit => VN_data_out(552),
        VN2CN1_bit => VN_data_out(553),
        VN2CN2_bit => VN_data_out(554),
        VN2CN3_bit => VN_data_out(555),
        VN2CN4_bit => VN_data_out(556),
        VN2CN5_bit => VN_data_out(557),
        VN2CN0_sign => VN_sign_out(552),
        VN2CN1_sign => VN_sign_out(553),
        VN2CN2_sign => VN_sign_out(554),
        VN2CN3_sign => VN_sign_out(555),
        VN2CN4_sign => VN_sign_out(556),
        VN2CN5_sign => VN_sign_out(557),
        codeword => codeword(92),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN93 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(563 downto 558),
        Din0 => VN93_in0,
        Din1 => VN93_in1,
        Din2 => VN93_in2,
        Din3 => VN93_in3,
        Din4 => VN93_in4,
        Din5 => VN93_in5,
        VN2CN0_bit => VN_data_out(558),
        VN2CN1_bit => VN_data_out(559),
        VN2CN2_bit => VN_data_out(560),
        VN2CN3_bit => VN_data_out(561),
        VN2CN4_bit => VN_data_out(562),
        VN2CN5_bit => VN_data_out(563),
        VN2CN0_sign => VN_sign_out(558),
        VN2CN1_sign => VN_sign_out(559),
        VN2CN2_sign => VN_sign_out(560),
        VN2CN3_sign => VN_sign_out(561),
        VN2CN4_sign => VN_sign_out(562),
        VN2CN5_sign => VN_sign_out(563),
        codeword => codeword(93),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN94 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(569 downto 564),
        Din0 => VN94_in0,
        Din1 => VN94_in1,
        Din2 => VN94_in2,
        Din3 => VN94_in3,
        Din4 => VN94_in4,
        Din5 => VN94_in5,
        VN2CN0_bit => VN_data_out(564),
        VN2CN1_bit => VN_data_out(565),
        VN2CN2_bit => VN_data_out(566),
        VN2CN3_bit => VN_data_out(567),
        VN2CN4_bit => VN_data_out(568),
        VN2CN5_bit => VN_data_out(569),
        VN2CN0_sign => VN_sign_out(564),
        VN2CN1_sign => VN_sign_out(565),
        VN2CN2_sign => VN_sign_out(566),
        VN2CN3_sign => VN_sign_out(567),
        VN2CN4_sign => VN_sign_out(568),
        VN2CN5_sign => VN_sign_out(569),
        codeword => codeword(94),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN95 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(575 downto 570),
        Din0 => VN95_in0,
        Din1 => VN95_in1,
        Din2 => VN95_in2,
        Din3 => VN95_in3,
        Din4 => VN95_in4,
        Din5 => VN95_in5,
        VN2CN0_bit => VN_data_out(570),
        VN2CN1_bit => VN_data_out(571),
        VN2CN2_bit => VN_data_out(572),
        VN2CN3_bit => VN_data_out(573),
        VN2CN4_bit => VN_data_out(574),
        VN2CN5_bit => VN_data_out(575),
        VN2CN0_sign => VN_sign_out(570),
        VN2CN1_sign => VN_sign_out(571),
        VN2CN2_sign => VN_sign_out(572),
        VN2CN3_sign => VN_sign_out(573),
        VN2CN4_sign => VN_sign_out(574),
        VN2CN5_sign => VN_sign_out(575),
        codeword => codeword(95),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN96 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(581 downto 576),
        Din0 => VN96_in0,
        Din1 => VN96_in1,
        Din2 => VN96_in2,
        Din3 => VN96_in3,
        Din4 => VN96_in4,
        Din5 => VN96_in5,
        VN2CN0_bit => VN_data_out(576),
        VN2CN1_bit => VN_data_out(577),
        VN2CN2_bit => VN_data_out(578),
        VN2CN3_bit => VN_data_out(579),
        VN2CN4_bit => VN_data_out(580),
        VN2CN5_bit => VN_data_out(581),
        VN2CN0_sign => VN_sign_out(576),
        VN2CN1_sign => VN_sign_out(577),
        VN2CN2_sign => VN_sign_out(578),
        VN2CN3_sign => VN_sign_out(579),
        VN2CN4_sign => VN_sign_out(580),
        VN2CN5_sign => VN_sign_out(581),
        codeword => codeword(96),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN97 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(587 downto 582),
        Din0 => VN97_in0,
        Din1 => VN97_in1,
        Din2 => VN97_in2,
        Din3 => VN97_in3,
        Din4 => VN97_in4,
        Din5 => VN97_in5,
        VN2CN0_bit => VN_data_out(582),
        VN2CN1_bit => VN_data_out(583),
        VN2CN2_bit => VN_data_out(584),
        VN2CN3_bit => VN_data_out(585),
        VN2CN4_bit => VN_data_out(586),
        VN2CN5_bit => VN_data_out(587),
        VN2CN0_sign => VN_sign_out(582),
        VN2CN1_sign => VN_sign_out(583),
        VN2CN2_sign => VN_sign_out(584),
        VN2CN3_sign => VN_sign_out(585),
        VN2CN4_sign => VN_sign_out(586),
        VN2CN5_sign => VN_sign_out(587),
        codeword => codeword(97),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN98 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(593 downto 588),
        Din0 => VN98_in0,
        Din1 => VN98_in1,
        Din2 => VN98_in2,
        Din3 => VN98_in3,
        Din4 => VN98_in4,
        Din5 => VN98_in5,
        VN2CN0_bit => VN_data_out(588),
        VN2CN1_bit => VN_data_out(589),
        VN2CN2_bit => VN_data_out(590),
        VN2CN3_bit => VN_data_out(591),
        VN2CN4_bit => VN_data_out(592),
        VN2CN5_bit => VN_data_out(593),
        VN2CN0_sign => VN_sign_out(588),
        VN2CN1_sign => VN_sign_out(589),
        VN2CN2_sign => VN_sign_out(590),
        VN2CN3_sign => VN_sign_out(591),
        VN2CN4_sign => VN_sign_out(592),
        VN2CN5_sign => VN_sign_out(593),
        codeword => codeword(98),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN99 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(599 downto 594),
        Din0 => VN99_in0,
        Din1 => VN99_in1,
        Din2 => VN99_in2,
        Din3 => VN99_in3,
        Din4 => VN99_in4,
        Din5 => VN99_in5,
        VN2CN0_bit => VN_data_out(594),
        VN2CN1_bit => VN_data_out(595),
        VN2CN2_bit => VN_data_out(596),
        VN2CN3_bit => VN_data_out(597),
        VN2CN4_bit => VN_data_out(598),
        VN2CN5_bit => VN_data_out(599),
        VN2CN0_sign => VN_sign_out(594),
        VN2CN1_sign => VN_sign_out(595),
        VN2CN2_sign => VN_sign_out(596),
        VN2CN3_sign => VN_sign_out(597),
        VN2CN4_sign => VN_sign_out(598),
        VN2CN5_sign => VN_sign_out(599),
        codeword => codeword(99),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN100 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(605 downto 600),
        Din0 => VN100_in0,
        Din1 => VN100_in1,
        Din2 => VN100_in2,
        Din3 => VN100_in3,
        Din4 => VN100_in4,
        Din5 => VN100_in5,
        VN2CN0_bit => VN_data_out(600),
        VN2CN1_bit => VN_data_out(601),
        VN2CN2_bit => VN_data_out(602),
        VN2CN3_bit => VN_data_out(603),
        VN2CN4_bit => VN_data_out(604),
        VN2CN5_bit => VN_data_out(605),
        VN2CN0_sign => VN_sign_out(600),
        VN2CN1_sign => VN_sign_out(601),
        VN2CN2_sign => VN_sign_out(602),
        VN2CN3_sign => VN_sign_out(603),
        VN2CN4_sign => VN_sign_out(604),
        VN2CN5_sign => VN_sign_out(605),
        codeword => codeword(100),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN101 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(611 downto 606),
        Din0 => VN101_in0,
        Din1 => VN101_in1,
        Din2 => VN101_in2,
        Din3 => VN101_in3,
        Din4 => VN101_in4,
        Din5 => VN101_in5,
        VN2CN0_bit => VN_data_out(606),
        VN2CN1_bit => VN_data_out(607),
        VN2CN2_bit => VN_data_out(608),
        VN2CN3_bit => VN_data_out(609),
        VN2CN4_bit => VN_data_out(610),
        VN2CN5_bit => VN_data_out(611),
        VN2CN0_sign => VN_sign_out(606),
        VN2CN1_sign => VN_sign_out(607),
        VN2CN2_sign => VN_sign_out(608),
        VN2CN3_sign => VN_sign_out(609),
        VN2CN4_sign => VN_sign_out(610),
        VN2CN5_sign => VN_sign_out(611),
        codeword => codeword(101),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN102 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(617 downto 612),
        Din0 => VN102_in0,
        Din1 => VN102_in1,
        Din2 => VN102_in2,
        Din3 => VN102_in3,
        Din4 => VN102_in4,
        Din5 => VN102_in5,
        VN2CN0_bit => VN_data_out(612),
        VN2CN1_bit => VN_data_out(613),
        VN2CN2_bit => VN_data_out(614),
        VN2CN3_bit => VN_data_out(615),
        VN2CN4_bit => VN_data_out(616),
        VN2CN5_bit => VN_data_out(617),
        VN2CN0_sign => VN_sign_out(612),
        VN2CN1_sign => VN_sign_out(613),
        VN2CN2_sign => VN_sign_out(614),
        VN2CN3_sign => VN_sign_out(615),
        VN2CN4_sign => VN_sign_out(616),
        VN2CN5_sign => VN_sign_out(617),
        codeword => codeword(102),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN103 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(623 downto 618),
        Din0 => VN103_in0,
        Din1 => VN103_in1,
        Din2 => VN103_in2,
        Din3 => VN103_in3,
        Din4 => VN103_in4,
        Din5 => VN103_in5,
        VN2CN0_bit => VN_data_out(618),
        VN2CN1_bit => VN_data_out(619),
        VN2CN2_bit => VN_data_out(620),
        VN2CN3_bit => VN_data_out(621),
        VN2CN4_bit => VN_data_out(622),
        VN2CN5_bit => VN_data_out(623),
        VN2CN0_sign => VN_sign_out(618),
        VN2CN1_sign => VN_sign_out(619),
        VN2CN2_sign => VN_sign_out(620),
        VN2CN3_sign => VN_sign_out(621),
        VN2CN4_sign => VN_sign_out(622),
        VN2CN5_sign => VN_sign_out(623),
        codeword => codeword(103),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN104 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(629 downto 624),
        Din0 => VN104_in0,
        Din1 => VN104_in1,
        Din2 => VN104_in2,
        Din3 => VN104_in3,
        Din4 => VN104_in4,
        Din5 => VN104_in5,
        VN2CN0_bit => VN_data_out(624),
        VN2CN1_bit => VN_data_out(625),
        VN2CN2_bit => VN_data_out(626),
        VN2CN3_bit => VN_data_out(627),
        VN2CN4_bit => VN_data_out(628),
        VN2CN5_bit => VN_data_out(629),
        VN2CN0_sign => VN_sign_out(624),
        VN2CN1_sign => VN_sign_out(625),
        VN2CN2_sign => VN_sign_out(626),
        VN2CN3_sign => VN_sign_out(627),
        VN2CN4_sign => VN_sign_out(628),
        VN2CN5_sign => VN_sign_out(629),
        codeword => codeword(104),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN105 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(635 downto 630),
        Din0 => VN105_in0,
        Din1 => VN105_in1,
        Din2 => VN105_in2,
        Din3 => VN105_in3,
        Din4 => VN105_in4,
        Din5 => VN105_in5,
        VN2CN0_bit => VN_data_out(630),
        VN2CN1_bit => VN_data_out(631),
        VN2CN2_bit => VN_data_out(632),
        VN2CN3_bit => VN_data_out(633),
        VN2CN4_bit => VN_data_out(634),
        VN2CN5_bit => VN_data_out(635),
        VN2CN0_sign => VN_sign_out(630),
        VN2CN1_sign => VN_sign_out(631),
        VN2CN2_sign => VN_sign_out(632),
        VN2CN3_sign => VN_sign_out(633),
        VN2CN4_sign => VN_sign_out(634),
        VN2CN5_sign => VN_sign_out(635),
        codeword => codeword(105),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN106 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(641 downto 636),
        Din0 => VN106_in0,
        Din1 => VN106_in1,
        Din2 => VN106_in2,
        Din3 => VN106_in3,
        Din4 => VN106_in4,
        Din5 => VN106_in5,
        VN2CN0_bit => VN_data_out(636),
        VN2CN1_bit => VN_data_out(637),
        VN2CN2_bit => VN_data_out(638),
        VN2CN3_bit => VN_data_out(639),
        VN2CN4_bit => VN_data_out(640),
        VN2CN5_bit => VN_data_out(641),
        VN2CN0_sign => VN_sign_out(636),
        VN2CN1_sign => VN_sign_out(637),
        VN2CN2_sign => VN_sign_out(638),
        VN2CN3_sign => VN_sign_out(639),
        VN2CN4_sign => VN_sign_out(640),
        VN2CN5_sign => VN_sign_out(641),
        codeword => codeword(106),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN107 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(647 downto 642),
        Din0 => VN107_in0,
        Din1 => VN107_in1,
        Din2 => VN107_in2,
        Din3 => VN107_in3,
        Din4 => VN107_in4,
        Din5 => VN107_in5,
        VN2CN0_bit => VN_data_out(642),
        VN2CN1_bit => VN_data_out(643),
        VN2CN2_bit => VN_data_out(644),
        VN2CN3_bit => VN_data_out(645),
        VN2CN4_bit => VN_data_out(646),
        VN2CN5_bit => VN_data_out(647),
        VN2CN0_sign => VN_sign_out(642),
        VN2CN1_sign => VN_sign_out(643),
        VN2CN2_sign => VN_sign_out(644),
        VN2CN3_sign => VN_sign_out(645),
        VN2CN4_sign => VN_sign_out(646),
        VN2CN5_sign => VN_sign_out(647),
        codeword => codeword(107),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN108 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(653 downto 648),
        Din0 => VN108_in0,
        Din1 => VN108_in1,
        Din2 => VN108_in2,
        Din3 => VN108_in3,
        Din4 => VN108_in4,
        Din5 => VN108_in5,
        VN2CN0_bit => VN_data_out(648),
        VN2CN1_bit => VN_data_out(649),
        VN2CN2_bit => VN_data_out(650),
        VN2CN3_bit => VN_data_out(651),
        VN2CN4_bit => VN_data_out(652),
        VN2CN5_bit => VN_data_out(653),
        VN2CN0_sign => VN_sign_out(648),
        VN2CN1_sign => VN_sign_out(649),
        VN2CN2_sign => VN_sign_out(650),
        VN2CN3_sign => VN_sign_out(651),
        VN2CN4_sign => VN_sign_out(652),
        VN2CN5_sign => VN_sign_out(653),
        codeword => codeword(108),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN109 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(659 downto 654),
        Din0 => VN109_in0,
        Din1 => VN109_in1,
        Din2 => VN109_in2,
        Din3 => VN109_in3,
        Din4 => VN109_in4,
        Din5 => VN109_in5,
        VN2CN0_bit => VN_data_out(654),
        VN2CN1_bit => VN_data_out(655),
        VN2CN2_bit => VN_data_out(656),
        VN2CN3_bit => VN_data_out(657),
        VN2CN4_bit => VN_data_out(658),
        VN2CN5_bit => VN_data_out(659),
        VN2CN0_sign => VN_sign_out(654),
        VN2CN1_sign => VN_sign_out(655),
        VN2CN2_sign => VN_sign_out(656),
        VN2CN3_sign => VN_sign_out(657),
        VN2CN4_sign => VN_sign_out(658),
        VN2CN5_sign => VN_sign_out(659),
        codeword => codeword(109),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN110 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(665 downto 660),
        Din0 => VN110_in0,
        Din1 => VN110_in1,
        Din2 => VN110_in2,
        Din3 => VN110_in3,
        Din4 => VN110_in4,
        Din5 => VN110_in5,
        VN2CN0_bit => VN_data_out(660),
        VN2CN1_bit => VN_data_out(661),
        VN2CN2_bit => VN_data_out(662),
        VN2CN3_bit => VN_data_out(663),
        VN2CN4_bit => VN_data_out(664),
        VN2CN5_bit => VN_data_out(665),
        VN2CN0_sign => VN_sign_out(660),
        VN2CN1_sign => VN_sign_out(661),
        VN2CN2_sign => VN_sign_out(662),
        VN2CN3_sign => VN_sign_out(663),
        VN2CN4_sign => VN_sign_out(664),
        VN2CN5_sign => VN_sign_out(665),
        codeword => codeword(110),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN111 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(671 downto 666),
        Din0 => VN111_in0,
        Din1 => VN111_in1,
        Din2 => VN111_in2,
        Din3 => VN111_in3,
        Din4 => VN111_in4,
        Din5 => VN111_in5,
        VN2CN0_bit => VN_data_out(666),
        VN2CN1_bit => VN_data_out(667),
        VN2CN2_bit => VN_data_out(668),
        VN2CN3_bit => VN_data_out(669),
        VN2CN4_bit => VN_data_out(670),
        VN2CN5_bit => VN_data_out(671),
        VN2CN0_sign => VN_sign_out(666),
        VN2CN1_sign => VN_sign_out(667),
        VN2CN2_sign => VN_sign_out(668),
        VN2CN3_sign => VN_sign_out(669),
        VN2CN4_sign => VN_sign_out(670),
        VN2CN5_sign => VN_sign_out(671),
        codeword => codeword(111),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN112 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(677 downto 672),
        Din0 => VN112_in0,
        Din1 => VN112_in1,
        Din2 => VN112_in2,
        Din3 => VN112_in3,
        Din4 => VN112_in4,
        Din5 => VN112_in5,
        VN2CN0_bit => VN_data_out(672),
        VN2CN1_bit => VN_data_out(673),
        VN2CN2_bit => VN_data_out(674),
        VN2CN3_bit => VN_data_out(675),
        VN2CN4_bit => VN_data_out(676),
        VN2CN5_bit => VN_data_out(677),
        VN2CN0_sign => VN_sign_out(672),
        VN2CN1_sign => VN_sign_out(673),
        VN2CN2_sign => VN_sign_out(674),
        VN2CN3_sign => VN_sign_out(675),
        VN2CN4_sign => VN_sign_out(676),
        VN2CN5_sign => VN_sign_out(677),
        codeword => codeword(112),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN113 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(683 downto 678),
        Din0 => VN113_in0,
        Din1 => VN113_in1,
        Din2 => VN113_in2,
        Din3 => VN113_in3,
        Din4 => VN113_in4,
        Din5 => VN113_in5,
        VN2CN0_bit => VN_data_out(678),
        VN2CN1_bit => VN_data_out(679),
        VN2CN2_bit => VN_data_out(680),
        VN2CN3_bit => VN_data_out(681),
        VN2CN4_bit => VN_data_out(682),
        VN2CN5_bit => VN_data_out(683),
        VN2CN0_sign => VN_sign_out(678),
        VN2CN1_sign => VN_sign_out(679),
        VN2CN2_sign => VN_sign_out(680),
        VN2CN3_sign => VN_sign_out(681),
        VN2CN4_sign => VN_sign_out(682),
        VN2CN5_sign => VN_sign_out(683),
        codeword => codeword(113),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN114 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(689 downto 684),
        Din0 => VN114_in0,
        Din1 => VN114_in1,
        Din2 => VN114_in2,
        Din3 => VN114_in3,
        Din4 => VN114_in4,
        Din5 => VN114_in5,
        VN2CN0_bit => VN_data_out(684),
        VN2CN1_bit => VN_data_out(685),
        VN2CN2_bit => VN_data_out(686),
        VN2CN3_bit => VN_data_out(687),
        VN2CN4_bit => VN_data_out(688),
        VN2CN5_bit => VN_data_out(689),
        VN2CN0_sign => VN_sign_out(684),
        VN2CN1_sign => VN_sign_out(685),
        VN2CN2_sign => VN_sign_out(686),
        VN2CN3_sign => VN_sign_out(687),
        VN2CN4_sign => VN_sign_out(688),
        VN2CN5_sign => VN_sign_out(689),
        codeword => codeword(114),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN115 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(695 downto 690),
        Din0 => VN115_in0,
        Din1 => VN115_in1,
        Din2 => VN115_in2,
        Din3 => VN115_in3,
        Din4 => VN115_in4,
        Din5 => VN115_in5,
        VN2CN0_bit => VN_data_out(690),
        VN2CN1_bit => VN_data_out(691),
        VN2CN2_bit => VN_data_out(692),
        VN2CN3_bit => VN_data_out(693),
        VN2CN4_bit => VN_data_out(694),
        VN2CN5_bit => VN_data_out(695),
        VN2CN0_sign => VN_sign_out(690),
        VN2CN1_sign => VN_sign_out(691),
        VN2CN2_sign => VN_sign_out(692),
        VN2CN3_sign => VN_sign_out(693),
        VN2CN4_sign => VN_sign_out(694),
        VN2CN5_sign => VN_sign_out(695),
        codeword => codeword(115),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN116 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(701 downto 696),
        Din0 => VN116_in0,
        Din1 => VN116_in1,
        Din2 => VN116_in2,
        Din3 => VN116_in3,
        Din4 => VN116_in4,
        Din5 => VN116_in5,
        VN2CN0_bit => VN_data_out(696),
        VN2CN1_bit => VN_data_out(697),
        VN2CN2_bit => VN_data_out(698),
        VN2CN3_bit => VN_data_out(699),
        VN2CN4_bit => VN_data_out(700),
        VN2CN5_bit => VN_data_out(701),
        VN2CN0_sign => VN_sign_out(696),
        VN2CN1_sign => VN_sign_out(697),
        VN2CN2_sign => VN_sign_out(698),
        VN2CN3_sign => VN_sign_out(699),
        VN2CN4_sign => VN_sign_out(700),
        VN2CN5_sign => VN_sign_out(701),
        codeword => codeword(116),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN117 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(707 downto 702),
        Din0 => VN117_in0,
        Din1 => VN117_in1,
        Din2 => VN117_in2,
        Din3 => VN117_in3,
        Din4 => VN117_in4,
        Din5 => VN117_in5,
        VN2CN0_bit => VN_data_out(702),
        VN2CN1_bit => VN_data_out(703),
        VN2CN2_bit => VN_data_out(704),
        VN2CN3_bit => VN_data_out(705),
        VN2CN4_bit => VN_data_out(706),
        VN2CN5_bit => VN_data_out(707),
        VN2CN0_sign => VN_sign_out(702),
        VN2CN1_sign => VN_sign_out(703),
        VN2CN2_sign => VN_sign_out(704),
        VN2CN3_sign => VN_sign_out(705),
        VN2CN4_sign => VN_sign_out(706),
        VN2CN5_sign => VN_sign_out(707),
        codeword => codeword(117),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN118 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(713 downto 708),
        Din0 => VN118_in0,
        Din1 => VN118_in1,
        Din2 => VN118_in2,
        Din3 => VN118_in3,
        Din4 => VN118_in4,
        Din5 => VN118_in5,
        VN2CN0_bit => VN_data_out(708),
        VN2CN1_bit => VN_data_out(709),
        VN2CN2_bit => VN_data_out(710),
        VN2CN3_bit => VN_data_out(711),
        VN2CN4_bit => VN_data_out(712),
        VN2CN5_bit => VN_data_out(713),
        VN2CN0_sign => VN_sign_out(708),
        VN2CN1_sign => VN_sign_out(709),
        VN2CN2_sign => VN_sign_out(710),
        VN2CN3_sign => VN_sign_out(711),
        VN2CN4_sign => VN_sign_out(712),
        VN2CN5_sign => VN_sign_out(713),
        codeword => codeword(118),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN119 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(719 downto 714),
        Din0 => VN119_in0,
        Din1 => VN119_in1,
        Din2 => VN119_in2,
        Din3 => VN119_in3,
        Din4 => VN119_in4,
        Din5 => VN119_in5,
        VN2CN0_bit => VN_data_out(714),
        VN2CN1_bit => VN_data_out(715),
        VN2CN2_bit => VN_data_out(716),
        VN2CN3_bit => VN_data_out(717),
        VN2CN4_bit => VN_data_out(718),
        VN2CN5_bit => VN_data_out(719),
        VN2CN0_sign => VN_sign_out(714),
        VN2CN1_sign => VN_sign_out(715),
        VN2CN2_sign => VN_sign_out(716),
        VN2CN3_sign => VN_sign_out(717),
        VN2CN4_sign => VN_sign_out(718),
        VN2CN5_sign => VN_sign_out(719),
        codeword => codeword(119),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN120 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(725 downto 720),
        Din0 => VN120_in0,
        Din1 => VN120_in1,
        Din2 => VN120_in2,
        Din3 => VN120_in3,
        Din4 => VN120_in4,
        Din5 => VN120_in5,
        VN2CN0_bit => VN_data_out(720),
        VN2CN1_bit => VN_data_out(721),
        VN2CN2_bit => VN_data_out(722),
        VN2CN3_bit => VN_data_out(723),
        VN2CN4_bit => VN_data_out(724),
        VN2CN5_bit => VN_data_out(725),
        VN2CN0_sign => VN_sign_out(720),
        VN2CN1_sign => VN_sign_out(721),
        VN2CN2_sign => VN_sign_out(722),
        VN2CN3_sign => VN_sign_out(723),
        VN2CN4_sign => VN_sign_out(724),
        VN2CN5_sign => VN_sign_out(725),
        codeword => codeword(120),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN121 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(731 downto 726),
        Din0 => VN121_in0,
        Din1 => VN121_in1,
        Din2 => VN121_in2,
        Din3 => VN121_in3,
        Din4 => VN121_in4,
        Din5 => VN121_in5,
        VN2CN0_bit => VN_data_out(726),
        VN2CN1_bit => VN_data_out(727),
        VN2CN2_bit => VN_data_out(728),
        VN2CN3_bit => VN_data_out(729),
        VN2CN4_bit => VN_data_out(730),
        VN2CN5_bit => VN_data_out(731),
        VN2CN0_sign => VN_sign_out(726),
        VN2CN1_sign => VN_sign_out(727),
        VN2CN2_sign => VN_sign_out(728),
        VN2CN3_sign => VN_sign_out(729),
        VN2CN4_sign => VN_sign_out(730),
        VN2CN5_sign => VN_sign_out(731),
        codeword => codeword(121),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN122 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(737 downto 732),
        Din0 => VN122_in0,
        Din1 => VN122_in1,
        Din2 => VN122_in2,
        Din3 => VN122_in3,
        Din4 => VN122_in4,
        Din5 => VN122_in5,
        VN2CN0_bit => VN_data_out(732),
        VN2CN1_bit => VN_data_out(733),
        VN2CN2_bit => VN_data_out(734),
        VN2CN3_bit => VN_data_out(735),
        VN2CN4_bit => VN_data_out(736),
        VN2CN5_bit => VN_data_out(737),
        VN2CN0_sign => VN_sign_out(732),
        VN2CN1_sign => VN_sign_out(733),
        VN2CN2_sign => VN_sign_out(734),
        VN2CN3_sign => VN_sign_out(735),
        VN2CN4_sign => VN_sign_out(736),
        VN2CN5_sign => VN_sign_out(737),
        codeword => codeword(122),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN123 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(743 downto 738),
        Din0 => VN123_in0,
        Din1 => VN123_in1,
        Din2 => VN123_in2,
        Din3 => VN123_in3,
        Din4 => VN123_in4,
        Din5 => VN123_in5,
        VN2CN0_bit => VN_data_out(738),
        VN2CN1_bit => VN_data_out(739),
        VN2CN2_bit => VN_data_out(740),
        VN2CN3_bit => VN_data_out(741),
        VN2CN4_bit => VN_data_out(742),
        VN2CN5_bit => VN_data_out(743),
        VN2CN0_sign => VN_sign_out(738),
        VN2CN1_sign => VN_sign_out(739),
        VN2CN2_sign => VN_sign_out(740),
        VN2CN3_sign => VN_sign_out(741),
        VN2CN4_sign => VN_sign_out(742),
        VN2CN5_sign => VN_sign_out(743),
        codeword => codeword(123),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN124 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(749 downto 744),
        Din0 => VN124_in0,
        Din1 => VN124_in1,
        Din2 => VN124_in2,
        Din3 => VN124_in3,
        Din4 => VN124_in4,
        Din5 => VN124_in5,
        VN2CN0_bit => VN_data_out(744),
        VN2CN1_bit => VN_data_out(745),
        VN2CN2_bit => VN_data_out(746),
        VN2CN3_bit => VN_data_out(747),
        VN2CN4_bit => VN_data_out(748),
        VN2CN5_bit => VN_data_out(749),
        VN2CN0_sign => VN_sign_out(744),
        VN2CN1_sign => VN_sign_out(745),
        VN2CN2_sign => VN_sign_out(746),
        VN2CN3_sign => VN_sign_out(747),
        VN2CN4_sign => VN_sign_out(748),
        VN2CN5_sign => VN_sign_out(749),
        codeword => codeword(124),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN125 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(755 downto 750),
        Din0 => VN125_in0,
        Din1 => VN125_in1,
        Din2 => VN125_in2,
        Din3 => VN125_in3,
        Din4 => VN125_in4,
        Din5 => VN125_in5,
        VN2CN0_bit => VN_data_out(750),
        VN2CN1_bit => VN_data_out(751),
        VN2CN2_bit => VN_data_out(752),
        VN2CN3_bit => VN_data_out(753),
        VN2CN4_bit => VN_data_out(754),
        VN2CN5_bit => VN_data_out(755),
        VN2CN0_sign => VN_sign_out(750),
        VN2CN1_sign => VN_sign_out(751),
        VN2CN2_sign => VN_sign_out(752),
        VN2CN3_sign => VN_sign_out(753),
        VN2CN4_sign => VN_sign_out(754),
        VN2CN5_sign => VN_sign_out(755),
        codeword => codeword(125),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN126 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(761 downto 756),
        Din0 => VN126_in0,
        Din1 => VN126_in1,
        Din2 => VN126_in2,
        Din3 => VN126_in3,
        Din4 => VN126_in4,
        Din5 => VN126_in5,
        VN2CN0_bit => VN_data_out(756),
        VN2CN1_bit => VN_data_out(757),
        VN2CN2_bit => VN_data_out(758),
        VN2CN3_bit => VN_data_out(759),
        VN2CN4_bit => VN_data_out(760),
        VN2CN5_bit => VN_data_out(761),
        VN2CN0_sign => VN_sign_out(756),
        VN2CN1_sign => VN_sign_out(757),
        VN2CN2_sign => VN_sign_out(758),
        VN2CN3_sign => VN_sign_out(759),
        VN2CN4_sign => VN_sign_out(760),
        VN2CN5_sign => VN_sign_out(761),
        codeword => codeword(126),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN127 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(767 downto 762),
        Din0 => VN127_in0,
        Din1 => VN127_in1,
        Din2 => VN127_in2,
        Din3 => VN127_in3,
        Din4 => VN127_in4,
        Din5 => VN127_in5,
        VN2CN0_bit => VN_data_out(762),
        VN2CN1_bit => VN_data_out(763),
        VN2CN2_bit => VN_data_out(764),
        VN2CN3_bit => VN_data_out(765),
        VN2CN4_bit => VN_data_out(766),
        VN2CN5_bit => VN_data_out(767),
        VN2CN0_sign => VN_sign_out(762),
        VN2CN1_sign => VN_sign_out(763),
        VN2CN2_sign => VN_sign_out(764),
        VN2CN3_sign => VN_sign_out(765),
        VN2CN4_sign => VN_sign_out(766),
        VN2CN5_sign => VN_sign_out(767),
        codeword => codeword(127),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN128 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(773 downto 768),
        Din0 => VN128_in0,
        Din1 => VN128_in1,
        Din2 => VN128_in2,
        Din3 => VN128_in3,
        Din4 => VN128_in4,
        Din5 => VN128_in5,
        VN2CN0_bit => VN_data_out(768),
        VN2CN1_bit => VN_data_out(769),
        VN2CN2_bit => VN_data_out(770),
        VN2CN3_bit => VN_data_out(771),
        VN2CN4_bit => VN_data_out(772),
        VN2CN5_bit => VN_data_out(773),
        VN2CN0_sign => VN_sign_out(768),
        VN2CN1_sign => VN_sign_out(769),
        VN2CN2_sign => VN_sign_out(770),
        VN2CN3_sign => VN_sign_out(771),
        VN2CN4_sign => VN_sign_out(772),
        VN2CN5_sign => VN_sign_out(773),
        codeword => codeword(128),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN129 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(779 downto 774),
        Din0 => VN129_in0,
        Din1 => VN129_in1,
        Din2 => VN129_in2,
        Din3 => VN129_in3,
        Din4 => VN129_in4,
        Din5 => VN129_in5,
        VN2CN0_bit => VN_data_out(774),
        VN2CN1_bit => VN_data_out(775),
        VN2CN2_bit => VN_data_out(776),
        VN2CN3_bit => VN_data_out(777),
        VN2CN4_bit => VN_data_out(778),
        VN2CN5_bit => VN_data_out(779),
        VN2CN0_sign => VN_sign_out(774),
        VN2CN1_sign => VN_sign_out(775),
        VN2CN2_sign => VN_sign_out(776),
        VN2CN3_sign => VN_sign_out(777),
        VN2CN4_sign => VN_sign_out(778),
        VN2CN5_sign => VN_sign_out(779),
        codeword => codeword(129),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN130 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(785 downto 780),
        Din0 => VN130_in0,
        Din1 => VN130_in1,
        Din2 => VN130_in2,
        Din3 => VN130_in3,
        Din4 => VN130_in4,
        Din5 => VN130_in5,
        VN2CN0_bit => VN_data_out(780),
        VN2CN1_bit => VN_data_out(781),
        VN2CN2_bit => VN_data_out(782),
        VN2CN3_bit => VN_data_out(783),
        VN2CN4_bit => VN_data_out(784),
        VN2CN5_bit => VN_data_out(785),
        VN2CN0_sign => VN_sign_out(780),
        VN2CN1_sign => VN_sign_out(781),
        VN2CN2_sign => VN_sign_out(782),
        VN2CN3_sign => VN_sign_out(783),
        VN2CN4_sign => VN_sign_out(784),
        VN2CN5_sign => VN_sign_out(785),
        codeword => codeword(130),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN131 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(791 downto 786),
        Din0 => VN131_in0,
        Din1 => VN131_in1,
        Din2 => VN131_in2,
        Din3 => VN131_in3,
        Din4 => VN131_in4,
        Din5 => VN131_in5,
        VN2CN0_bit => VN_data_out(786),
        VN2CN1_bit => VN_data_out(787),
        VN2CN2_bit => VN_data_out(788),
        VN2CN3_bit => VN_data_out(789),
        VN2CN4_bit => VN_data_out(790),
        VN2CN5_bit => VN_data_out(791),
        VN2CN0_sign => VN_sign_out(786),
        VN2CN1_sign => VN_sign_out(787),
        VN2CN2_sign => VN_sign_out(788),
        VN2CN3_sign => VN_sign_out(789),
        VN2CN4_sign => VN_sign_out(790),
        VN2CN5_sign => VN_sign_out(791),
        codeword => codeword(131),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN132 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(797 downto 792),
        Din0 => VN132_in0,
        Din1 => VN132_in1,
        Din2 => VN132_in2,
        Din3 => VN132_in3,
        Din4 => VN132_in4,
        Din5 => VN132_in5,
        VN2CN0_bit => VN_data_out(792),
        VN2CN1_bit => VN_data_out(793),
        VN2CN2_bit => VN_data_out(794),
        VN2CN3_bit => VN_data_out(795),
        VN2CN4_bit => VN_data_out(796),
        VN2CN5_bit => VN_data_out(797),
        VN2CN0_sign => VN_sign_out(792),
        VN2CN1_sign => VN_sign_out(793),
        VN2CN2_sign => VN_sign_out(794),
        VN2CN3_sign => VN_sign_out(795),
        VN2CN4_sign => VN_sign_out(796),
        VN2CN5_sign => VN_sign_out(797),
        codeword => codeword(132),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN133 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(803 downto 798),
        Din0 => VN133_in0,
        Din1 => VN133_in1,
        Din2 => VN133_in2,
        Din3 => VN133_in3,
        Din4 => VN133_in4,
        Din5 => VN133_in5,
        VN2CN0_bit => VN_data_out(798),
        VN2CN1_bit => VN_data_out(799),
        VN2CN2_bit => VN_data_out(800),
        VN2CN3_bit => VN_data_out(801),
        VN2CN4_bit => VN_data_out(802),
        VN2CN5_bit => VN_data_out(803),
        VN2CN0_sign => VN_sign_out(798),
        VN2CN1_sign => VN_sign_out(799),
        VN2CN2_sign => VN_sign_out(800),
        VN2CN3_sign => VN_sign_out(801),
        VN2CN4_sign => VN_sign_out(802),
        VN2CN5_sign => VN_sign_out(803),
        codeword => codeword(133),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN134 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(809 downto 804),
        Din0 => VN134_in0,
        Din1 => VN134_in1,
        Din2 => VN134_in2,
        Din3 => VN134_in3,
        Din4 => VN134_in4,
        Din5 => VN134_in5,
        VN2CN0_bit => VN_data_out(804),
        VN2CN1_bit => VN_data_out(805),
        VN2CN2_bit => VN_data_out(806),
        VN2CN3_bit => VN_data_out(807),
        VN2CN4_bit => VN_data_out(808),
        VN2CN5_bit => VN_data_out(809),
        VN2CN0_sign => VN_sign_out(804),
        VN2CN1_sign => VN_sign_out(805),
        VN2CN2_sign => VN_sign_out(806),
        VN2CN3_sign => VN_sign_out(807),
        VN2CN4_sign => VN_sign_out(808),
        VN2CN5_sign => VN_sign_out(809),
        codeword => codeword(134),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN135 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(815 downto 810),
        Din0 => VN135_in0,
        Din1 => VN135_in1,
        Din2 => VN135_in2,
        Din3 => VN135_in3,
        Din4 => VN135_in4,
        Din5 => VN135_in5,
        VN2CN0_bit => VN_data_out(810),
        VN2CN1_bit => VN_data_out(811),
        VN2CN2_bit => VN_data_out(812),
        VN2CN3_bit => VN_data_out(813),
        VN2CN4_bit => VN_data_out(814),
        VN2CN5_bit => VN_data_out(815),
        VN2CN0_sign => VN_sign_out(810),
        VN2CN1_sign => VN_sign_out(811),
        VN2CN2_sign => VN_sign_out(812),
        VN2CN3_sign => VN_sign_out(813),
        VN2CN4_sign => VN_sign_out(814),
        VN2CN5_sign => VN_sign_out(815),
        codeword => codeword(135),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN136 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(821 downto 816),
        Din0 => VN136_in0,
        Din1 => VN136_in1,
        Din2 => VN136_in2,
        Din3 => VN136_in3,
        Din4 => VN136_in4,
        Din5 => VN136_in5,
        VN2CN0_bit => VN_data_out(816),
        VN2CN1_bit => VN_data_out(817),
        VN2CN2_bit => VN_data_out(818),
        VN2CN3_bit => VN_data_out(819),
        VN2CN4_bit => VN_data_out(820),
        VN2CN5_bit => VN_data_out(821),
        VN2CN0_sign => VN_sign_out(816),
        VN2CN1_sign => VN_sign_out(817),
        VN2CN2_sign => VN_sign_out(818),
        VN2CN3_sign => VN_sign_out(819),
        VN2CN4_sign => VN_sign_out(820),
        VN2CN5_sign => VN_sign_out(821),
        codeword => codeword(136),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN137 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(827 downto 822),
        Din0 => VN137_in0,
        Din1 => VN137_in1,
        Din2 => VN137_in2,
        Din3 => VN137_in3,
        Din4 => VN137_in4,
        Din5 => VN137_in5,
        VN2CN0_bit => VN_data_out(822),
        VN2CN1_bit => VN_data_out(823),
        VN2CN2_bit => VN_data_out(824),
        VN2CN3_bit => VN_data_out(825),
        VN2CN4_bit => VN_data_out(826),
        VN2CN5_bit => VN_data_out(827),
        VN2CN0_sign => VN_sign_out(822),
        VN2CN1_sign => VN_sign_out(823),
        VN2CN2_sign => VN_sign_out(824),
        VN2CN3_sign => VN_sign_out(825),
        VN2CN4_sign => VN_sign_out(826),
        VN2CN5_sign => VN_sign_out(827),
        codeword => codeword(137),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN138 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(833 downto 828),
        Din0 => VN138_in0,
        Din1 => VN138_in1,
        Din2 => VN138_in2,
        Din3 => VN138_in3,
        Din4 => VN138_in4,
        Din5 => VN138_in5,
        VN2CN0_bit => VN_data_out(828),
        VN2CN1_bit => VN_data_out(829),
        VN2CN2_bit => VN_data_out(830),
        VN2CN3_bit => VN_data_out(831),
        VN2CN4_bit => VN_data_out(832),
        VN2CN5_bit => VN_data_out(833),
        VN2CN0_sign => VN_sign_out(828),
        VN2CN1_sign => VN_sign_out(829),
        VN2CN2_sign => VN_sign_out(830),
        VN2CN3_sign => VN_sign_out(831),
        VN2CN4_sign => VN_sign_out(832),
        VN2CN5_sign => VN_sign_out(833),
        codeword => codeword(138),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN139 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(839 downto 834),
        Din0 => VN139_in0,
        Din1 => VN139_in1,
        Din2 => VN139_in2,
        Din3 => VN139_in3,
        Din4 => VN139_in4,
        Din5 => VN139_in5,
        VN2CN0_bit => VN_data_out(834),
        VN2CN1_bit => VN_data_out(835),
        VN2CN2_bit => VN_data_out(836),
        VN2CN3_bit => VN_data_out(837),
        VN2CN4_bit => VN_data_out(838),
        VN2CN5_bit => VN_data_out(839),
        VN2CN0_sign => VN_sign_out(834),
        VN2CN1_sign => VN_sign_out(835),
        VN2CN2_sign => VN_sign_out(836),
        VN2CN3_sign => VN_sign_out(837),
        VN2CN4_sign => VN_sign_out(838),
        VN2CN5_sign => VN_sign_out(839),
        codeword => codeword(139),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN140 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(845 downto 840),
        Din0 => VN140_in0,
        Din1 => VN140_in1,
        Din2 => VN140_in2,
        Din3 => VN140_in3,
        Din4 => VN140_in4,
        Din5 => VN140_in5,
        VN2CN0_bit => VN_data_out(840),
        VN2CN1_bit => VN_data_out(841),
        VN2CN2_bit => VN_data_out(842),
        VN2CN3_bit => VN_data_out(843),
        VN2CN4_bit => VN_data_out(844),
        VN2CN5_bit => VN_data_out(845),
        VN2CN0_sign => VN_sign_out(840),
        VN2CN1_sign => VN_sign_out(841),
        VN2CN2_sign => VN_sign_out(842),
        VN2CN3_sign => VN_sign_out(843),
        VN2CN4_sign => VN_sign_out(844),
        VN2CN5_sign => VN_sign_out(845),
        codeword => codeword(140),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN141 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(851 downto 846),
        Din0 => VN141_in0,
        Din1 => VN141_in1,
        Din2 => VN141_in2,
        Din3 => VN141_in3,
        Din4 => VN141_in4,
        Din5 => VN141_in5,
        VN2CN0_bit => VN_data_out(846),
        VN2CN1_bit => VN_data_out(847),
        VN2CN2_bit => VN_data_out(848),
        VN2CN3_bit => VN_data_out(849),
        VN2CN4_bit => VN_data_out(850),
        VN2CN5_bit => VN_data_out(851),
        VN2CN0_sign => VN_sign_out(846),
        VN2CN1_sign => VN_sign_out(847),
        VN2CN2_sign => VN_sign_out(848),
        VN2CN3_sign => VN_sign_out(849),
        VN2CN4_sign => VN_sign_out(850),
        VN2CN5_sign => VN_sign_out(851),
        codeword => codeword(141),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN142 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(857 downto 852),
        Din0 => VN142_in0,
        Din1 => VN142_in1,
        Din2 => VN142_in2,
        Din3 => VN142_in3,
        Din4 => VN142_in4,
        Din5 => VN142_in5,
        VN2CN0_bit => VN_data_out(852),
        VN2CN1_bit => VN_data_out(853),
        VN2CN2_bit => VN_data_out(854),
        VN2CN3_bit => VN_data_out(855),
        VN2CN4_bit => VN_data_out(856),
        VN2CN5_bit => VN_data_out(857),
        VN2CN0_sign => VN_sign_out(852),
        VN2CN1_sign => VN_sign_out(853),
        VN2CN2_sign => VN_sign_out(854),
        VN2CN3_sign => VN_sign_out(855),
        VN2CN4_sign => VN_sign_out(856),
        VN2CN5_sign => VN_sign_out(857),
        codeword => codeword(142),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN143 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(863 downto 858),
        Din0 => VN143_in0,
        Din1 => VN143_in1,
        Din2 => VN143_in2,
        Din3 => VN143_in3,
        Din4 => VN143_in4,
        Din5 => VN143_in5,
        VN2CN0_bit => VN_data_out(858),
        VN2CN1_bit => VN_data_out(859),
        VN2CN2_bit => VN_data_out(860),
        VN2CN3_bit => VN_data_out(861),
        VN2CN4_bit => VN_data_out(862),
        VN2CN5_bit => VN_data_out(863),
        VN2CN0_sign => VN_sign_out(858),
        VN2CN1_sign => VN_sign_out(859),
        VN2CN2_sign => VN_sign_out(860),
        VN2CN3_sign => VN_sign_out(861),
        VN2CN4_sign => VN_sign_out(862),
        VN2CN5_sign => VN_sign_out(863),
        codeword => codeword(143),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN144 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(869 downto 864),
        Din0 => VN144_in0,
        Din1 => VN144_in1,
        Din2 => VN144_in2,
        Din3 => VN144_in3,
        Din4 => VN144_in4,
        Din5 => VN144_in5,
        VN2CN0_bit => VN_data_out(864),
        VN2CN1_bit => VN_data_out(865),
        VN2CN2_bit => VN_data_out(866),
        VN2CN3_bit => VN_data_out(867),
        VN2CN4_bit => VN_data_out(868),
        VN2CN5_bit => VN_data_out(869),
        VN2CN0_sign => VN_sign_out(864),
        VN2CN1_sign => VN_sign_out(865),
        VN2CN2_sign => VN_sign_out(866),
        VN2CN3_sign => VN_sign_out(867),
        VN2CN4_sign => VN_sign_out(868),
        VN2CN5_sign => VN_sign_out(869),
        codeword => codeword(144),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN145 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(875 downto 870),
        Din0 => VN145_in0,
        Din1 => VN145_in1,
        Din2 => VN145_in2,
        Din3 => VN145_in3,
        Din4 => VN145_in4,
        Din5 => VN145_in5,
        VN2CN0_bit => VN_data_out(870),
        VN2CN1_bit => VN_data_out(871),
        VN2CN2_bit => VN_data_out(872),
        VN2CN3_bit => VN_data_out(873),
        VN2CN4_bit => VN_data_out(874),
        VN2CN5_bit => VN_data_out(875),
        VN2CN0_sign => VN_sign_out(870),
        VN2CN1_sign => VN_sign_out(871),
        VN2CN2_sign => VN_sign_out(872),
        VN2CN3_sign => VN_sign_out(873),
        VN2CN4_sign => VN_sign_out(874),
        VN2CN5_sign => VN_sign_out(875),
        codeword => codeword(145),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN146 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(881 downto 876),
        Din0 => VN146_in0,
        Din1 => VN146_in1,
        Din2 => VN146_in2,
        Din3 => VN146_in3,
        Din4 => VN146_in4,
        Din5 => VN146_in5,
        VN2CN0_bit => VN_data_out(876),
        VN2CN1_bit => VN_data_out(877),
        VN2CN2_bit => VN_data_out(878),
        VN2CN3_bit => VN_data_out(879),
        VN2CN4_bit => VN_data_out(880),
        VN2CN5_bit => VN_data_out(881),
        VN2CN0_sign => VN_sign_out(876),
        VN2CN1_sign => VN_sign_out(877),
        VN2CN2_sign => VN_sign_out(878),
        VN2CN3_sign => VN_sign_out(879),
        VN2CN4_sign => VN_sign_out(880),
        VN2CN5_sign => VN_sign_out(881),
        codeword => codeword(146),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN147 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(887 downto 882),
        Din0 => VN147_in0,
        Din1 => VN147_in1,
        Din2 => VN147_in2,
        Din3 => VN147_in3,
        Din4 => VN147_in4,
        Din5 => VN147_in5,
        VN2CN0_bit => VN_data_out(882),
        VN2CN1_bit => VN_data_out(883),
        VN2CN2_bit => VN_data_out(884),
        VN2CN3_bit => VN_data_out(885),
        VN2CN4_bit => VN_data_out(886),
        VN2CN5_bit => VN_data_out(887),
        VN2CN0_sign => VN_sign_out(882),
        VN2CN1_sign => VN_sign_out(883),
        VN2CN2_sign => VN_sign_out(884),
        VN2CN3_sign => VN_sign_out(885),
        VN2CN4_sign => VN_sign_out(886),
        VN2CN5_sign => VN_sign_out(887),
        codeword => codeword(147),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN148 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(893 downto 888),
        Din0 => VN148_in0,
        Din1 => VN148_in1,
        Din2 => VN148_in2,
        Din3 => VN148_in3,
        Din4 => VN148_in4,
        Din5 => VN148_in5,
        VN2CN0_bit => VN_data_out(888),
        VN2CN1_bit => VN_data_out(889),
        VN2CN2_bit => VN_data_out(890),
        VN2CN3_bit => VN_data_out(891),
        VN2CN4_bit => VN_data_out(892),
        VN2CN5_bit => VN_data_out(893),
        VN2CN0_sign => VN_sign_out(888),
        VN2CN1_sign => VN_sign_out(889),
        VN2CN2_sign => VN_sign_out(890),
        VN2CN3_sign => VN_sign_out(891),
        VN2CN4_sign => VN_sign_out(892),
        VN2CN5_sign => VN_sign_out(893),
        codeword => codeword(148),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN149 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(899 downto 894),
        Din0 => VN149_in0,
        Din1 => VN149_in1,
        Din2 => VN149_in2,
        Din3 => VN149_in3,
        Din4 => VN149_in4,
        Din5 => VN149_in5,
        VN2CN0_bit => VN_data_out(894),
        VN2CN1_bit => VN_data_out(895),
        VN2CN2_bit => VN_data_out(896),
        VN2CN3_bit => VN_data_out(897),
        VN2CN4_bit => VN_data_out(898),
        VN2CN5_bit => VN_data_out(899),
        VN2CN0_sign => VN_sign_out(894),
        VN2CN1_sign => VN_sign_out(895),
        VN2CN2_sign => VN_sign_out(896),
        VN2CN3_sign => VN_sign_out(897),
        VN2CN4_sign => VN_sign_out(898),
        VN2CN5_sign => VN_sign_out(899),
        codeword => codeword(149),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN150 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(905 downto 900),
        Din0 => VN150_in0,
        Din1 => VN150_in1,
        Din2 => VN150_in2,
        Din3 => VN150_in3,
        Din4 => VN150_in4,
        Din5 => VN150_in5,
        VN2CN0_bit => VN_data_out(900),
        VN2CN1_bit => VN_data_out(901),
        VN2CN2_bit => VN_data_out(902),
        VN2CN3_bit => VN_data_out(903),
        VN2CN4_bit => VN_data_out(904),
        VN2CN5_bit => VN_data_out(905),
        VN2CN0_sign => VN_sign_out(900),
        VN2CN1_sign => VN_sign_out(901),
        VN2CN2_sign => VN_sign_out(902),
        VN2CN3_sign => VN_sign_out(903),
        VN2CN4_sign => VN_sign_out(904),
        VN2CN5_sign => VN_sign_out(905),
        codeword => codeword(150),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN151 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(911 downto 906),
        Din0 => VN151_in0,
        Din1 => VN151_in1,
        Din2 => VN151_in2,
        Din3 => VN151_in3,
        Din4 => VN151_in4,
        Din5 => VN151_in5,
        VN2CN0_bit => VN_data_out(906),
        VN2CN1_bit => VN_data_out(907),
        VN2CN2_bit => VN_data_out(908),
        VN2CN3_bit => VN_data_out(909),
        VN2CN4_bit => VN_data_out(910),
        VN2CN5_bit => VN_data_out(911),
        VN2CN0_sign => VN_sign_out(906),
        VN2CN1_sign => VN_sign_out(907),
        VN2CN2_sign => VN_sign_out(908),
        VN2CN3_sign => VN_sign_out(909),
        VN2CN4_sign => VN_sign_out(910),
        VN2CN5_sign => VN_sign_out(911),
        codeword => codeword(151),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN152 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(917 downto 912),
        Din0 => VN152_in0,
        Din1 => VN152_in1,
        Din2 => VN152_in2,
        Din3 => VN152_in3,
        Din4 => VN152_in4,
        Din5 => VN152_in5,
        VN2CN0_bit => VN_data_out(912),
        VN2CN1_bit => VN_data_out(913),
        VN2CN2_bit => VN_data_out(914),
        VN2CN3_bit => VN_data_out(915),
        VN2CN4_bit => VN_data_out(916),
        VN2CN5_bit => VN_data_out(917),
        VN2CN0_sign => VN_sign_out(912),
        VN2CN1_sign => VN_sign_out(913),
        VN2CN2_sign => VN_sign_out(914),
        VN2CN3_sign => VN_sign_out(915),
        VN2CN4_sign => VN_sign_out(916),
        VN2CN5_sign => VN_sign_out(917),
        codeword => codeword(152),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN153 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(923 downto 918),
        Din0 => VN153_in0,
        Din1 => VN153_in1,
        Din2 => VN153_in2,
        Din3 => VN153_in3,
        Din4 => VN153_in4,
        Din5 => VN153_in5,
        VN2CN0_bit => VN_data_out(918),
        VN2CN1_bit => VN_data_out(919),
        VN2CN2_bit => VN_data_out(920),
        VN2CN3_bit => VN_data_out(921),
        VN2CN4_bit => VN_data_out(922),
        VN2CN5_bit => VN_data_out(923),
        VN2CN0_sign => VN_sign_out(918),
        VN2CN1_sign => VN_sign_out(919),
        VN2CN2_sign => VN_sign_out(920),
        VN2CN3_sign => VN_sign_out(921),
        VN2CN4_sign => VN_sign_out(922),
        VN2CN5_sign => VN_sign_out(923),
        codeword => codeword(153),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN154 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(929 downto 924),
        Din0 => VN154_in0,
        Din1 => VN154_in1,
        Din2 => VN154_in2,
        Din3 => VN154_in3,
        Din4 => VN154_in4,
        Din5 => VN154_in5,
        VN2CN0_bit => VN_data_out(924),
        VN2CN1_bit => VN_data_out(925),
        VN2CN2_bit => VN_data_out(926),
        VN2CN3_bit => VN_data_out(927),
        VN2CN4_bit => VN_data_out(928),
        VN2CN5_bit => VN_data_out(929),
        VN2CN0_sign => VN_sign_out(924),
        VN2CN1_sign => VN_sign_out(925),
        VN2CN2_sign => VN_sign_out(926),
        VN2CN3_sign => VN_sign_out(927),
        VN2CN4_sign => VN_sign_out(928),
        VN2CN5_sign => VN_sign_out(929),
        codeword => codeword(154),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN155 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(935 downto 930),
        Din0 => VN155_in0,
        Din1 => VN155_in1,
        Din2 => VN155_in2,
        Din3 => VN155_in3,
        Din4 => VN155_in4,
        Din5 => VN155_in5,
        VN2CN0_bit => VN_data_out(930),
        VN2CN1_bit => VN_data_out(931),
        VN2CN2_bit => VN_data_out(932),
        VN2CN3_bit => VN_data_out(933),
        VN2CN4_bit => VN_data_out(934),
        VN2CN5_bit => VN_data_out(935),
        VN2CN0_sign => VN_sign_out(930),
        VN2CN1_sign => VN_sign_out(931),
        VN2CN2_sign => VN_sign_out(932),
        VN2CN3_sign => VN_sign_out(933),
        VN2CN4_sign => VN_sign_out(934),
        VN2CN5_sign => VN_sign_out(935),
        codeword => codeword(155),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN156 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(941 downto 936),
        Din0 => VN156_in0,
        Din1 => VN156_in1,
        Din2 => VN156_in2,
        Din3 => VN156_in3,
        Din4 => VN156_in4,
        Din5 => VN156_in5,
        VN2CN0_bit => VN_data_out(936),
        VN2CN1_bit => VN_data_out(937),
        VN2CN2_bit => VN_data_out(938),
        VN2CN3_bit => VN_data_out(939),
        VN2CN4_bit => VN_data_out(940),
        VN2CN5_bit => VN_data_out(941),
        VN2CN0_sign => VN_sign_out(936),
        VN2CN1_sign => VN_sign_out(937),
        VN2CN2_sign => VN_sign_out(938),
        VN2CN3_sign => VN_sign_out(939),
        VN2CN4_sign => VN_sign_out(940),
        VN2CN5_sign => VN_sign_out(941),
        codeword => codeword(156),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN157 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(947 downto 942),
        Din0 => VN157_in0,
        Din1 => VN157_in1,
        Din2 => VN157_in2,
        Din3 => VN157_in3,
        Din4 => VN157_in4,
        Din5 => VN157_in5,
        VN2CN0_bit => VN_data_out(942),
        VN2CN1_bit => VN_data_out(943),
        VN2CN2_bit => VN_data_out(944),
        VN2CN3_bit => VN_data_out(945),
        VN2CN4_bit => VN_data_out(946),
        VN2CN5_bit => VN_data_out(947),
        VN2CN0_sign => VN_sign_out(942),
        VN2CN1_sign => VN_sign_out(943),
        VN2CN2_sign => VN_sign_out(944),
        VN2CN3_sign => VN_sign_out(945),
        VN2CN4_sign => VN_sign_out(946),
        VN2CN5_sign => VN_sign_out(947),
        codeword => codeword(157),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN158 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(953 downto 948),
        Din0 => VN158_in0,
        Din1 => VN158_in1,
        Din2 => VN158_in2,
        Din3 => VN158_in3,
        Din4 => VN158_in4,
        Din5 => VN158_in5,
        VN2CN0_bit => VN_data_out(948),
        VN2CN1_bit => VN_data_out(949),
        VN2CN2_bit => VN_data_out(950),
        VN2CN3_bit => VN_data_out(951),
        VN2CN4_bit => VN_data_out(952),
        VN2CN5_bit => VN_data_out(953),
        VN2CN0_sign => VN_sign_out(948),
        VN2CN1_sign => VN_sign_out(949),
        VN2CN2_sign => VN_sign_out(950),
        VN2CN3_sign => VN_sign_out(951),
        VN2CN4_sign => VN_sign_out(952),
        VN2CN5_sign => VN_sign_out(953),
        codeword => codeword(158),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN159 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(959 downto 954),
        Din0 => VN159_in0,
        Din1 => VN159_in1,
        Din2 => VN159_in2,
        Din3 => VN159_in3,
        Din4 => VN159_in4,
        Din5 => VN159_in5,
        VN2CN0_bit => VN_data_out(954),
        VN2CN1_bit => VN_data_out(955),
        VN2CN2_bit => VN_data_out(956),
        VN2CN3_bit => VN_data_out(957),
        VN2CN4_bit => VN_data_out(958),
        VN2CN5_bit => VN_data_out(959),
        VN2CN0_sign => VN_sign_out(954),
        VN2CN1_sign => VN_sign_out(955),
        VN2CN2_sign => VN_sign_out(956),
        VN2CN3_sign => VN_sign_out(957),
        VN2CN4_sign => VN_sign_out(958),
        VN2CN5_sign => VN_sign_out(959),
        codeword => codeword(159),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN160 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(965 downto 960),
        Din0 => VN160_in0,
        Din1 => VN160_in1,
        Din2 => VN160_in2,
        Din3 => VN160_in3,
        Din4 => VN160_in4,
        Din5 => VN160_in5,
        VN2CN0_bit => VN_data_out(960),
        VN2CN1_bit => VN_data_out(961),
        VN2CN2_bit => VN_data_out(962),
        VN2CN3_bit => VN_data_out(963),
        VN2CN4_bit => VN_data_out(964),
        VN2CN5_bit => VN_data_out(965),
        VN2CN0_sign => VN_sign_out(960),
        VN2CN1_sign => VN_sign_out(961),
        VN2CN2_sign => VN_sign_out(962),
        VN2CN3_sign => VN_sign_out(963),
        VN2CN4_sign => VN_sign_out(964),
        VN2CN5_sign => VN_sign_out(965),
        codeword => codeword(160),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN161 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(971 downto 966),
        Din0 => VN161_in0,
        Din1 => VN161_in1,
        Din2 => VN161_in2,
        Din3 => VN161_in3,
        Din4 => VN161_in4,
        Din5 => VN161_in5,
        VN2CN0_bit => VN_data_out(966),
        VN2CN1_bit => VN_data_out(967),
        VN2CN2_bit => VN_data_out(968),
        VN2CN3_bit => VN_data_out(969),
        VN2CN4_bit => VN_data_out(970),
        VN2CN5_bit => VN_data_out(971),
        VN2CN0_sign => VN_sign_out(966),
        VN2CN1_sign => VN_sign_out(967),
        VN2CN2_sign => VN_sign_out(968),
        VN2CN3_sign => VN_sign_out(969),
        VN2CN4_sign => VN_sign_out(970),
        VN2CN5_sign => VN_sign_out(971),
        codeword => codeword(161),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN162 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(977 downto 972),
        Din0 => VN162_in0,
        Din1 => VN162_in1,
        Din2 => VN162_in2,
        Din3 => VN162_in3,
        Din4 => VN162_in4,
        Din5 => VN162_in5,
        VN2CN0_bit => VN_data_out(972),
        VN2CN1_bit => VN_data_out(973),
        VN2CN2_bit => VN_data_out(974),
        VN2CN3_bit => VN_data_out(975),
        VN2CN4_bit => VN_data_out(976),
        VN2CN5_bit => VN_data_out(977),
        VN2CN0_sign => VN_sign_out(972),
        VN2CN1_sign => VN_sign_out(973),
        VN2CN2_sign => VN_sign_out(974),
        VN2CN3_sign => VN_sign_out(975),
        VN2CN4_sign => VN_sign_out(976),
        VN2CN5_sign => VN_sign_out(977),
        codeword => codeword(162),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN163 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(983 downto 978),
        Din0 => VN163_in0,
        Din1 => VN163_in1,
        Din2 => VN163_in2,
        Din3 => VN163_in3,
        Din4 => VN163_in4,
        Din5 => VN163_in5,
        VN2CN0_bit => VN_data_out(978),
        VN2CN1_bit => VN_data_out(979),
        VN2CN2_bit => VN_data_out(980),
        VN2CN3_bit => VN_data_out(981),
        VN2CN4_bit => VN_data_out(982),
        VN2CN5_bit => VN_data_out(983),
        VN2CN0_sign => VN_sign_out(978),
        VN2CN1_sign => VN_sign_out(979),
        VN2CN2_sign => VN_sign_out(980),
        VN2CN3_sign => VN_sign_out(981),
        VN2CN4_sign => VN_sign_out(982),
        VN2CN5_sign => VN_sign_out(983),
        codeword => codeword(163),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN164 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(989 downto 984),
        Din0 => VN164_in0,
        Din1 => VN164_in1,
        Din2 => VN164_in2,
        Din3 => VN164_in3,
        Din4 => VN164_in4,
        Din5 => VN164_in5,
        VN2CN0_bit => VN_data_out(984),
        VN2CN1_bit => VN_data_out(985),
        VN2CN2_bit => VN_data_out(986),
        VN2CN3_bit => VN_data_out(987),
        VN2CN4_bit => VN_data_out(988),
        VN2CN5_bit => VN_data_out(989),
        VN2CN0_sign => VN_sign_out(984),
        VN2CN1_sign => VN_sign_out(985),
        VN2CN2_sign => VN_sign_out(986),
        VN2CN3_sign => VN_sign_out(987),
        VN2CN4_sign => VN_sign_out(988),
        VN2CN5_sign => VN_sign_out(989),
        codeword => codeword(164),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN165 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(995 downto 990),
        Din0 => VN165_in0,
        Din1 => VN165_in1,
        Din2 => VN165_in2,
        Din3 => VN165_in3,
        Din4 => VN165_in4,
        Din5 => VN165_in5,
        VN2CN0_bit => VN_data_out(990),
        VN2CN1_bit => VN_data_out(991),
        VN2CN2_bit => VN_data_out(992),
        VN2CN3_bit => VN_data_out(993),
        VN2CN4_bit => VN_data_out(994),
        VN2CN5_bit => VN_data_out(995),
        VN2CN0_sign => VN_sign_out(990),
        VN2CN1_sign => VN_sign_out(991),
        VN2CN2_sign => VN_sign_out(992),
        VN2CN3_sign => VN_sign_out(993),
        VN2CN4_sign => VN_sign_out(994),
        VN2CN5_sign => VN_sign_out(995),
        codeword => codeword(165),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN166 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1001 downto 996),
        Din0 => VN166_in0,
        Din1 => VN166_in1,
        Din2 => VN166_in2,
        Din3 => VN166_in3,
        Din4 => VN166_in4,
        Din5 => VN166_in5,
        VN2CN0_bit => VN_data_out(996),
        VN2CN1_bit => VN_data_out(997),
        VN2CN2_bit => VN_data_out(998),
        VN2CN3_bit => VN_data_out(999),
        VN2CN4_bit => VN_data_out(1000),
        VN2CN5_bit => VN_data_out(1001),
        VN2CN0_sign => VN_sign_out(996),
        VN2CN1_sign => VN_sign_out(997),
        VN2CN2_sign => VN_sign_out(998),
        VN2CN3_sign => VN_sign_out(999),
        VN2CN4_sign => VN_sign_out(1000),
        VN2CN5_sign => VN_sign_out(1001),
        codeword => codeword(166),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN167 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1007 downto 1002),
        Din0 => VN167_in0,
        Din1 => VN167_in1,
        Din2 => VN167_in2,
        Din3 => VN167_in3,
        Din4 => VN167_in4,
        Din5 => VN167_in5,
        VN2CN0_bit => VN_data_out(1002),
        VN2CN1_bit => VN_data_out(1003),
        VN2CN2_bit => VN_data_out(1004),
        VN2CN3_bit => VN_data_out(1005),
        VN2CN4_bit => VN_data_out(1006),
        VN2CN5_bit => VN_data_out(1007),
        VN2CN0_sign => VN_sign_out(1002),
        VN2CN1_sign => VN_sign_out(1003),
        VN2CN2_sign => VN_sign_out(1004),
        VN2CN3_sign => VN_sign_out(1005),
        VN2CN4_sign => VN_sign_out(1006),
        VN2CN5_sign => VN_sign_out(1007),
        codeword => codeword(167),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN168 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1013 downto 1008),
        Din0 => VN168_in0,
        Din1 => VN168_in1,
        Din2 => VN168_in2,
        Din3 => VN168_in3,
        Din4 => VN168_in4,
        Din5 => VN168_in5,
        VN2CN0_bit => VN_data_out(1008),
        VN2CN1_bit => VN_data_out(1009),
        VN2CN2_bit => VN_data_out(1010),
        VN2CN3_bit => VN_data_out(1011),
        VN2CN4_bit => VN_data_out(1012),
        VN2CN5_bit => VN_data_out(1013),
        VN2CN0_sign => VN_sign_out(1008),
        VN2CN1_sign => VN_sign_out(1009),
        VN2CN2_sign => VN_sign_out(1010),
        VN2CN3_sign => VN_sign_out(1011),
        VN2CN4_sign => VN_sign_out(1012),
        VN2CN5_sign => VN_sign_out(1013),
        codeword => codeword(168),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN169 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1019 downto 1014),
        Din0 => VN169_in0,
        Din1 => VN169_in1,
        Din2 => VN169_in2,
        Din3 => VN169_in3,
        Din4 => VN169_in4,
        Din5 => VN169_in5,
        VN2CN0_bit => VN_data_out(1014),
        VN2CN1_bit => VN_data_out(1015),
        VN2CN2_bit => VN_data_out(1016),
        VN2CN3_bit => VN_data_out(1017),
        VN2CN4_bit => VN_data_out(1018),
        VN2CN5_bit => VN_data_out(1019),
        VN2CN0_sign => VN_sign_out(1014),
        VN2CN1_sign => VN_sign_out(1015),
        VN2CN2_sign => VN_sign_out(1016),
        VN2CN3_sign => VN_sign_out(1017),
        VN2CN4_sign => VN_sign_out(1018),
        VN2CN5_sign => VN_sign_out(1019),
        codeword => codeword(169),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN170 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1025 downto 1020),
        Din0 => VN170_in0,
        Din1 => VN170_in1,
        Din2 => VN170_in2,
        Din3 => VN170_in3,
        Din4 => VN170_in4,
        Din5 => VN170_in5,
        VN2CN0_bit => VN_data_out(1020),
        VN2CN1_bit => VN_data_out(1021),
        VN2CN2_bit => VN_data_out(1022),
        VN2CN3_bit => VN_data_out(1023),
        VN2CN4_bit => VN_data_out(1024),
        VN2CN5_bit => VN_data_out(1025),
        VN2CN0_sign => VN_sign_out(1020),
        VN2CN1_sign => VN_sign_out(1021),
        VN2CN2_sign => VN_sign_out(1022),
        VN2CN3_sign => VN_sign_out(1023),
        VN2CN4_sign => VN_sign_out(1024),
        VN2CN5_sign => VN_sign_out(1025),
        codeword => codeword(170),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN171 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1031 downto 1026),
        Din0 => VN171_in0,
        Din1 => VN171_in1,
        Din2 => VN171_in2,
        Din3 => VN171_in3,
        Din4 => VN171_in4,
        Din5 => VN171_in5,
        VN2CN0_bit => VN_data_out(1026),
        VN2CN1_bit => VN_data_out(1027),
        VN2CN2_bit => VN_data_out(1028),
        VN2CN3_bit => VN_data_out(1029),
        VN2CN4_bit => VN_data_out(1030),
        VN2CN5_bit => VN_data_out(1031),
        VN2CN0_sign => VN_sign_out(1026),
        VN2CN1_sign => VN_sign_out(1027),
        VN2CN2_sign => VN_sign_out(1028),
        VN2CN3_sign => VN_sign_out(1029),
        VN2CN4_sign => VN_sign_out(1030),
        VN2CN5_sign => VN_sign_out(1031),
        codeword => codeword(171),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN172 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1037 downto 1032),
        Din0 => VN172_in0,
        Din1 => VN172_in1,
        Din2 => VN172_in2,
        Din3 => VN172_in3,
        Din4 => VN172_in4,
        Din5 => VN172_in5,
        VN2CN0_bit => VN_data_out(1032),
        VN2CN1_bit => VN_data_out(1033),
        VN2CN2_bit => VN_data_out(1034),
        VN2CN3_bit => VN_data_out(1035),
        VN2CN4_bit => VN_data_out(1036),
        VN2CN5_bit => VN_data_out(1037),
        VN2CN0_sign => VN_sign_out(1032),
        VN2CN1_sign => VN_sign_out(1033),
        VN2CN2_sign => VN_sign_out(1034),
        VN2CN3_sign => VN_sign_out(1035),
        VN2CN4_sign => VN_sign_out(1036),
        VN2CN5_sign => VN_sign_out(1037),
        codeword => codeword(172),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN173 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1043 downto 1038),
        Din0 => VN173_in0,
        Din1 => VN173_in1,
        Din2 => VN173_in2,
        Din3 => VN173_in3,
        Din4 => VN173_in4,
        Din5 => VN173_in5,
        VN2CN0_bit => VN_data_out(1038),
        VN2CN1_bit => VN_data_out(1039),
        VN2CN2_bit => VN_data_out(1040),
        VN2CN3_bit => VN_data_out(1041),
        VN2CN4_bit => VN_data_out(1042),
        VN2CN5_bit => VN_data_out(1043),
        VN2CN0_sign => VN_sign_out(1038),
        VN2CN1_sign => VN_sign_out(1039),
        VN2CN2_sign => VN_sign_out(1040),
        VN2CN3_sign => VN_sign_out(1041),
        VN2CN4_sign => VN_sign_out(1042),
        VN2CN5_sign => VN_sign_out(1043),
        codeword => codeword(173),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN174 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1049 downto 1044),
        Din0 => VN174_in0,
        Din1 => VN174_in1,
        Din2 => VN174_in2,
        Din3 => VN174_in3,
        Din4 => VN174_in4,
        Din5 => VN174_in5,
        VN2CN0_bit => VN_data_out(1044),
        VN2CN1_bit => VN_data_out(1045),
        VN2CN2_bit => VN_data_out(1046),
        VN2CN3_bit => VN_data_out(1047),
        VN2CN4_bit => VN_data_out(1048),
        VN2CN5_bit => VN_data_out(1049),
        VN2CN0_sign => VN_sign_out(1044),
        VN2CN1_sign => VN_sign_out(1045),
        VN2CN2_sign => VN_sign_out(1046),
        VN2CN3_sign => VN_sign_out(1047),
        VN2CN4_sign => VN_sign_out(1048),
        VN2CN5_sign => VN_sign_out(1049),
        codeword => codeword(174),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN175 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1055 downto 1050),
        Din0 => VN175_in0,
        Din1 => VN175_in1,
        Din2 => VN175_in2,
        Din3 => VN175_in3,
        Din4 => VN175_in4,
        Din5 => VN175_in5,
        VN2CN0_bit => VN_data_out(1050),
        VN2CN1_bit => VN_data_out(1051),
        VN2CN2_bit => VN_data_out(1052),
        VN2CN3_bit => VN_data_out(1053),
        VN2CN4_bit => VN_data_out(1054),
        VN2CN5_bit => VN_data_out(1055),
        VN2CN0_sign => VN_sign_out(1050),
        VN2CN1_sign => VN_sign_out(1051),
        VN2CN2_sign => VN_sign_out(1052),
        VN2CN3_sign => VN_sign_out(1053),
        VN2CN4_sign => VN_sign_out(1054),
        VN2CN5_sign => VN_sign_out(1055),
        codeword => codeword(175),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN176 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1061 downto 1056),
        Din0 => VN176_in0,
        Din1 => VN176_in1,
        Din2 => VN176_in2,
        Din3 => VN176_in3,
        Din4 => VN176_in4,
        Din5 => VN176_in5,
        VN2CN0_bit => VN_data_out(1056),
        VN2CN1_bit => VN_data_out(1057),
        VN2CN2_bit => VN_data_out(1058),
        VN2CN3_bit => VN_data_out(1059),
        VN2CN4_bit => VN_data_out(1060),
        VN2CN5_bit => VN_data_out(1061),
        VN2CN0_sign => VN_sign_out(1056),
        VN2CN1_sign => VN_sign_out(1057),
        VN2CN2_sign => VN_sign_out(1058),
        VN2CN3_sign => VN_sign_out(1059),
        VN2CN4_sign => VN_sign_out(1060),
        VN2CN5_sign => VN_sign_out(1061),
        codeword => codeword(176),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN177 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1067 downto 1062),
        Din0 => VN177_in0,
        Din1 => VN177_in1,
        Din2 => VN177_in2,
        Din3 => VN177_in3,
        Din4 => VN177_in4,
        Din5 => VN177_in5,
        VN2CN0_bit => VN_data_out(1062),
        VN2CN1_bit => VN_data_out(1063),
        VN2CN2_bit => VN_data_out(1064),
        VN2CN3_bit => VN_data_out(1065),
        VN2CN4_bit => VN_data_out(1066),
        VN2CN5_bit => VN_data_out(1067),
        VN2CN0_sign => VN_sign_out(1062),
        VN2CN1_sign => VN_sign_out(1063),
        VN2CN2_sign => VN_sign_out(1064),
        VN2CN3_sign => VN_sign_out(1065),
        VN2CN4_sign => VN_sign_out(1066),
        VN2CN5_sign => VN_sign_out(1067),
        codeword => codeword(177),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN178 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1073 downto 1068),
        Din0 => VN178_in0,
        Din1 => VN178_in1,
        Din2 => VN178_in2,
        Din3 => VN178_in3,
        Din4 => VN178_in4,
        Din5 => VN178_in5,
        VN2CN0_bit => VN_data_out(1068),
        VN2CN1_bit => VN_data_out(1069),
        VN2CN2_bit => VN_data_out(1070),
        VN2CN3_bit => VN_data_out(1071),
        VN2CN4_bit => VN_data_out(1072),
        VN2CN5_bit => VN_data_out(1073),
        VN2CN0_sign => VN_sign_out(1068),
        VN2CN1_sign => VN_sign_out(1069),
        VN2CN2_sign => VN_sign_out(1070),
        VN2CN3_sign => VN_sign_out(1071),
        VN2CN4_sign => VN_sign_out(1072),
        VN2CN5_sign => VN_sign_out(1073),
        codeword => codeword(178),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN179 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1079 downto 1074),
        Din0 => VN179_in0,
        Din1 => VN179_in1,
        Din2 => VN179_in2,
        Din3 => VN179_in3,
        Din4 => VN179_in4,
        Din5 => VN179_in5,
        VN2CN0_bit => VN_data_out(1074),
        VN2CN1_bit => VN_data_out(1075),
        VN2CN2_bit => VN_data_out(1076),
        VN2CN3_bit => VN_data_out(1077),
        VN2CN4_bit => VN_data_out(1078),
        VN2CN5_bit => VN_data_out(1079),
        VN2CN0_sign => VN_sign_out(1074),
        VN2CN1_sign => VN_sign_out(1075),
        VN2CN2_sign => VN_sign_out(1076),
        VN2CN3_sign => VN_sign_out(1077),
        VN2CN4_sign => VN_sign_out(1078),
        VN2CN5_sign => VN_sign_out(1079),
        codeword => codeword(179),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN180 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1085 downto 1080),
        Din0 => VN180_in0,
        Din1 => VN180_in1,
        Din2 => VN180_in2,
        Din3 => VN180_in3,
        Din4 => VN180_in4,
        Din5 => VN180_in5,
        VN2CN0_bit => VN_data_out(1080),
        VN2CN1_bit => VN_data_out(1081),
        VN2CN2_bit => VN_data_out(1082),
        VN2CN3_bit => VN_data_out(1083),
        VN2CN4_bit => VN_data_out(1084),
        VN2CN5_bit => VN_data_out(1085),
        VN2CN0_sign => VN_sign_out(1080),
        VN2CN1_sign => VN_sign_out(1081),
        VN2CN2_sign => VN_sign_out(1082),
        VN2CN3_sign => VN_sign_out(1083),
        VN2CN4_sign => VN_sign_out(1084),
        VN2CN5_sign => VN_sign_out(1085),
        codeword => codeword(180),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN181 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1091 downto 1086),
        Din0 => VN181_in0,
        Din1 => VN181_in1,
        Din2 => VN181_in2,
        Din3 => VN181_in3,
        Din4 => VN181_in4,
        Din5 => VN181_in5,
        VN2CN0_bit => VN_data_out(1086),
        VN2CN1_bit => VN_data_out(1087),
        VN2CN2_bit => VN_data_out(1088),
        VN2CN3_bit => VN_data_out(1089),
        VN2CN4_bit => VN_data_out(1090),
        VN2CN5_bit => VN_data_out(1091),
        VN2CN0_sign => VN_sign_out(1086),
        VN2CN1_sign => VN_sign_out(1087),
        VN2CN2_sign => VN_sign_out(1088),
        VN2CN3_sign => VN_sign_out(1089),
        VN2CN4_sign => VN_sign_out(1090),
        VN2CN5_sign => VN_sign_out(1091),
        codeword => codeword(181),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN182 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1097 downto 1092),
        Din0 => VN182_in0,
        Din1 => VN182_in1,
        Din2 => VN182_in2,
        Din3 => VN182_in3,
        Din4 => VN182_in4,
        Din5 => VN182_in5,
        VN2CN0_bit => VN_data_out(1092),
        VN2CN1_bit => VN_data_out(1093),
        VN2CN2_bit => VN_data_out(1094),
        VN2CN3_bit => VN_data_out(1095),
        VN2CN4_bit => VN_data_out(1096),
        VN2CN5_bit => VN_data_out(1097),
        VN2CN0_sign => VN_sign_out(1092),
        VN2CN1_sign => VN_sign_out(1093),
        VN2CN2_sign => VN_sign_out(1094),
        VN2CN3_sign => VN_sign_out(1095),
        VN2CN4_sign => VN_sign_out(1096),
        VN2CN5_sign => VN_sign_out(1097),
        codeword => codeword(182),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN183 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1103 downto 1098),
        Din0 => VN183_in0,
        Din1 => VN183_in1,
        Din2 => VN183_in2,
        Din3 => VN183_in3,
        Din4 => VN183_in4,
        Din5 => VN183_in5,
        VN2CN0_bit => VN_data_out(1098),
        VN2CN1_bit => VN_data_out(1099),
        VN2CN2_bit => VN_data_out(1100),
        VN2CN3_bit => VN_data_out(1101),
        VN2CN4_bit => VN_data_out(1102),
        VN2CN5_bit => VN_data_out(1103),
        VN2CN0_sign => VN_sign_out(1098),
        VN2CN1_sign => VN_sign_out(1099),
        VN2CN2_sign => VN_sign_out(1100),
        VN2CN3_sign => VN_sign_out(1101),
        VN2CN4_sign => VN_sign_out(1102),
        VN2CN5_sign => VN_sign_out(1103),
        codeword => codeword(183),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN184 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1109 downto 1104),
        Din0 => VN184_in0,
        Din1 => VN184_in1,
        Din2 => VN184_in2,
        Din3 => VN184_in3,
        Din4 => VN184_in4,
        Din5 => VN184_in5,
        VN2CN0_bit => VN_data_out(1104),
        VN2CN1_bit => VN_data_out(1105),
        VN2CN2_bit => VN_data_out(1106),
        VN2CN3_bit => VN_data_out(1107),
        VN2CN4_bit => VN_data_out(1108),
        VN2CN5_bit => VN_data_out(1109),
        VN2CN0_sign => VN_sign_out(1104),
        VN2CN1_sign => VN_sign_out(1105),
        VN2CN2_sign => VN_sign_out(1106),
        VN2CN3_sign => VN_sign_out(1107),
        VN2CN4_sign => VN_sign_out(1108),
        VN2CN5_sign => VN_sign_out(1109),
        codeword => codeword(184),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN185 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1115 downto 1110),
        Din0 => VN185_in0,
        Din1 => VN185_in1,
        Din2 => VN185_in2,
        Din3 => VN185_in3,
        Din4 => VN185_in4,
        Din5 => VN185_in5,
        VN2CN0_bit => VN_data_out(1110),
        VN2CN1_bit => VN_data_out(1111),
        VN2CN2_bit => VN_data_out(1112),
        VN2CN3_bit => VN_data_out(1113),
        VN2CN4_bit => VN_data_out(1114),
        VN2CN5_bit => VN_data_out(1115),
        VN2CN0_sign => VN_sign_out(1110),
        VN2CN1_sign => VN_sign_out(1111),
        VN2CN2_sign => VN_sign_out(1112),
        VN2CN3_sign => VN_sign_out(1113),
        VN2CN4_sign => VN_sign_out(1114),
        VN2CN5_sign => VN_sign_out(1115),
        codeword => codeword(185),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN186 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1121 downto 1116),
        Din0 => VN186_in0,
        Din1 => VN186_in1,
        Din2 => VN186_in2,
        Din3 => VN186_in3,
        Din4 => VN186_in4,
        Din5 => VN186_in5,
        VN2CN0_bit => VN_data_out(1116),
        VN2CN1_bit => VN_data_out(1117),
        VN2CN2_bit => VN_data_out(1118),
        VN2CN3_bit => VN_data_out(1119),
        VN2CN4_bit => VN_data_out(1120),
        VN2CN5_bit => VN_data_out(1121),
        VN2CN0_sign => VN_sign_out(1116),
        VN2CN1_sign => VN_sign_out(1117),
        VN2CN2_sign => VN_sign_out(1118),
        VN2CN3_sign => VN_sign_out(1119),
        VN2CN4_sign => VN_sign_out(1120),
        VN2CN5_sign => VN_sign_out(1121),
        codeword => codeword(186),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN187 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1127 downto 1122),
        Din0 => VN187_in0,
        Din1 => VN187_in1,
        Din2 => VN187_in2,
        Din3 => VN187_in3,
        Din4 => VN187_in4,
        Din5 => VN187_in5,
        VN2CN0_bit => VN_data_out(1122),
        VN2CN1_bit => VN_data_out(1123),
        VN2CN2_bit => VN_data_out(1124),
        VN2CN3_bit => VN_data_out(1125),
        VN2CN4_bit => VN_data_out(1126),
        VN2CN5_bit => VN_data_out(1127),
        VN2CN0_sign => VN_sign_out(1122),
        VN2CN1_sign => VN_sign_out(1123),
        VN2CN2_sign => VN_sign_out(1124),
        VN2CN3_sign => VN_sign_out(1125),
        VN2CN4_sign => VN_sign_out(1126),
        VN2CN5_sign => VN_sign_out(1127),
        codeword => codeword(187),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN188 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1133 downto 1128),
        Din0 => VN188_in0,
        Din1 => VN188_in1,
        Din2 => VN188_in2,
        Din3 => VN188_in3,
        Din4 => VN188_in4,
        Din5 => VN188_in5,
        VN2CN0_bit => VN_data_out(1128),
        VN2CN1_bit => VN_data_out(1129),
        VN2CN2_bit => VN_data_out(1130),
        VN2CN3_bit => VN_data_out(1131),
        VN2CN4_bit => VN_data_out(1132),
        VN2CN5_bit => VN_data_out(1133),
        VN2CN0_sign => VN_sign_out(1128),
        VN2CN1_sign => VN_sign_out(1129),
        VN2CN2_sign => VN_sign_out(1130),
        VN2CN3_sign => VN_sign_out(1131),
        VN2CN4_sign => VN_sign_out(1132),
        VN2CN5_sign => VN_sign_out(1133),
        codeword => codeword(188),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN189 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1139 downto 1134),
        Din0 => VN189_in0,
        Din1 => VN189_in1,
        Din2 => VN189_in2,
        Din3 => VN189_in3,
        Din4 => VN189_in4,
        Din5 => VN189_in5,
        VN2CN0_bit => VN_data_out(1134),
        VN2CN1_bit => VN_data_out(1135),
        VN2CN2_bit => VN_data_out(1136),
        VN2CN3_bit => VN_data_out(1137),
        VN2CN4_bit => VN_data_out(1138),
        VN2CN5_bit => VN_data_out(1139),
        VN2CN0_sign => VN_sign_out(1134),
        VN2CN1_sign => VN_sign_out(1135),
        VN2CN2_sign => VN_sign_out(1136),
        VN2CN3_sign => VN_sign_out(1137),
        VN2CN4_sign => VN_sign_out(1138),
        VN2CN5_sign => VN_sign_out(1139),
        codeword => codeword(189),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN190 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1145 downto 1140),
        Din0 => VN190_in0,
        Din1 => VN190_in1,
        Din2 => VN190_in2,
        Din3 => VN190_in3,
        Din4 => VN190_in4,
        Din5 => VN190_in5,
        VN2CN0_bit => VN_data_out(1140),
        VN2CN1_bit => VN_data_out(1141),
        VN2CN2_bit => VN_data_out(1142),
        VN2CN3_bit => VN_data_out(1143),
        VN2CN4_bit => VN_data_out(1144),
        VN2CN5_bit => VN_data_out(1145),
        VN2CN0_sign => VN_sign_out(1140),
        VN2CN1_sign => VN_sign_out(1141),
        VN2CN2_sign => VN_sign_out(1142),
        VN2CN3_sign => VN_sign_out(1143),
        VN2CN4_sign => VN_sign_out(1144),
        VN2CN5_sign => VN_sign_out(1145),
        codeword => codeword(190),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN191 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1151 downto 1146),
        Din0 => VN191_in0,
        Din1 => VN191_in1,
        Din2 => VN191_in2,
        Din3 => VN191_in3,
        Din4 => VN191_in4,
        Din5 => VN191_in5,
        VN2CN0_bit => VN_data_out(1146),
        VN2CN1_bit => VN_data_out(1147),
        VN2CN2_bit => VN_data_out(1148),
        VN2CN3_bit => VN_data_out(1149),
        VN2CN4_bit => VN_data_out(1150),
        VN2CN5_bit => VN_data_out(1151),
        VN2CN0_sign => VN_sign_out(1146),
        VN2CN1_sign => VN_sign_out(1147),
        VN2CN2_sign => VN_sign_out(1148),
        VN2CN3_sign => VN_sign_out(1149),
        VN2CN4_sign => VN_sign_out(1150),
        VN2CN5_sign => VN_sign_out(1151),
        codeword => codeword(191),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN192 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1157 downto 1152),
        Din0 => VN192_in0,
        Din1 => VN192_in1,
        Din2 => VN192_in2,
        Din3 => VN192_in3,
        Din4 => VN192_in4,
        Din5 => VN192_in5,
        VN2CN0_bit => VN_data_out(1152),
        VN2CN1_bit => VN_data_out(1153),
        VN2CN2_bit => VN_data_out(1154),
        VN2CN3_bit => VN_data_out(1155),
        VN2CN4_bit => VN_data_out(1156),
        VN2CN5_bit => VN_data_out(1157),
        VN2CN0_sign => VN_sign_out(1152),
        VN2CN1_sign => VN_sign_out(1153),
        VN2CN2_sign => VN_sign_out(1154),
        VN2CN3_sign => VN_sign_out(1155),
        VN2CN4_sign => VN_sign_out(1156),
        VN2CN5_sign => VN_sign_out(1157),
        codeword => codeword(192),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN193 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1163 downto 1158),
        Din0 => VN193_in0,
        Din1 => VN193_in1,
        Din2 => VN193_in2,
        Din3 => VN193_in3,
        Din4 => VN193_in4,
        Din5 => VN193_in5,
        VN2CN0_bit => VN_data_out(1158),
        VN2CN1_bit => VN_data_out(1159),
        VN2CN2_bit => VN_data_out(1160),
        VN2CN3_bit => VN_data_out(1161),
        VN2CN4_bit => VN_data_out(1162),
        VN2CN5_bit => VN_data_out(1163),
        VN2CN0_sign => VN_sign_out(1158),
        VN2CN1_sign => VN_sign_out(1159),
        VN2CN2_sign => VN_sign_out(1160),
        VN2CN3_sign => VN_sign_out(1161),
        VN2CN4_sign => VN_sign_out(1162),
        VN2CN5_sign => VN_sign_out(1163),
        codeword => codeword(193),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN194 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1169 downto 1164),
        Din0 => VN194_in0,
        Din1 => VN194_in1,
        Din2 => VN194_in2,
        Din3 => VN194_in3,
        Din4 => VN194_in4,
        Din5 => VN194_in5,
        VN2CN0_bit => VN_data_out(1164),
        VN2CN1_bit => VN_data_out(1165),
        VN2CN2_bit => VN_data_out(1166),
        VN2CN3_bit => VN_data_out(1167),
        VN2CN4_bit => VN_data_out(1168),
        VN2CN5_bit => VN_data_out(1169),
        VN2CN0_sign => VN_sign_out(1164),
        VN2CN1_sign => VN_sign_out(1165),
        VN2CN2_sign => VN_sign_out(1166),
        VN2CN3_sign => VN_sign_out(1167),
        VN2CN4_sign => VN_sign_out(1168),
        VN2CN5_sign => VN_sign_out(1169),
        codeword => codeword(194),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN195 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1175 downto 1170),
        Din0 => VN195_in0,
        Din1 => VN195_in1,
        Din2 => VN195_in2,
        Din3 => VN195_in3,
        Din4 => VN195_in4,
        Din5 => VN195_in5,
        VN2CN0_bit => VN_data_out(1170),
        VN2CN1_bit => VN_data_out(1171),
        VN2CN2_bit => VN_data_out(1172),
        VN2CN3_bit => VN_data_out(1173),
        VN2CN4_bit => VN_data_out(1174),
        VN2CN5_bit => VN_data_out(1175),
        VN2CN0_sign => VN_sign_out(1170),
        VN2CN1_sign => VN_sign_out(1171),
        VN2CN2_sign => VN_sign_out(1172),
        VN2CN3_sign => VN_sign_out(1173),
        VN2CN4_sign => VN_sign_out(1174),
        VN2CN5_sign => VN_sign_out(1175),
        codeword => codeword(195),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN196 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1181 downto 1176),
        Din0 => VN196_in0,
        Din1 => VN196_in1,
        Din2 => VN196_in2,
        Din3 => VN196_in3,
        Din4 => VN196_in4,
        Din5 => VN196_in5,
        VN2CN0_bit => VN_data_out(1176),
        VN2CN1_bit => VN_data_out(1177),
        VN2CN2_bit => VN_data_out(1178),
        VN2CN3_bit => VN_data_out(1179),
        VN2CN4_bit => VN_data_out(1180),
        VN2CN5_bit => VN_data_out(1181),
        VN2CN0_sign => VN_sign_out(1176),
        VN2CN1_sign => VN_sign_out(1177),
        VN2CN2_sign => VN_sign_out(1178),
        VN2CN3_sign => VN_sign_out(1179),
        VN2CN4_sign => VN_sign_out(1180),
        VN2CN5_sign => VN_sign_out(1181),
        codeword => codeword(196),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN197 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1187 downto 1182),
        Din0 => VN197_in0,
        Din1 => VN197_in1,
        Din2 => VN197_in2,
        Din3 => VN197_in3,
        Din4 => VN197_in4,
        Din5 => VN197_in5,
        VN2CN0_bit => VN_data_out(1182),
        VN2CN1_bit => VN_data_out(1183),
        VN2CN2_bit => VN_data_out(1184),
        VN2CN3_bit => VN_data_out(1185),
        VN2CN4_bit => VN_data_out(1186),
        VN2CN5_bit => VN_data_out(1187),
        VN2CN0_sign => VN_sign_out(1182),
        VN2CN1_sign => VN_sign_out(1183),
        VN2CN2_sign => VN_sign_out(1184),
        VN2CN3_sign => VN_sign_out(1185),
        VN2CN4_sign => VN_sign_out(1186),
        VN2CN5_sign => VN_sign_out(1187),
        codeword => codeword(197),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN198 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1193 downto 1188),
        Din0 => VN198_in0,
        Din1 => VN198_in1,
        Din2 => VN198_in2,
        Din3 => VN198_in3,
        Din4 => VN198_in4,
        Din5 => VN198_in5,
        VN2CN0_bit => VN_data_out(1188),
        VN2CN1_bit => VN_data_out(1189),
        VN2CN2_bit => VN_data_out(1190),
        VN2CN3_bit => VN_data_out(1191),
        VN2CN4_bit => VN_data_out(1192),
        VN2CN5_bit => VN_data_out(1193),
        VN2CN0_sign => VN_sign_out(1188),
        VN2CN1_sign => VN_sign_out(1189),
        VN2CN2_sign => VN_sign_out(1190),
        VN2CN3_sign => VN_sign_out(1191),
        VN2CN4_sign => VN_sign_out(1192),
        VN2CN5_sign => VN_sign_out(1193),
        codeword => codeword(198),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN199 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1199 downto 1194),
        Din0 => VN199_in0,
        Din1 => VN199_in1,
        Din2 => VN199_in2,
        Din3 => VN199_in3,
        Din4 => VN199_in4,
        Din5 => VN199_in5,
        VN2CN0_bit => VN_data_out(1194),
        VN2CN1_bit => VN_data_out(1195),
        VN2CN2_bit => VN_data_out(1196),
        VN2CN3_bit => VN_data_out(1197),
        VN2CN4_bit => VN_data_out(1198),
        VN2CN5_bit => VN_data_out(1199),
        VN2CN0_sign => VN_sign_out(1194),
        VN2CN1_sign => VN_sign_out(1195),
        VN2CN2_sign => VN_sign_out(1196),
        VN2CN3_sign => VN_sign_out(1197),
        VN2CN4_sign => VN_sign_out(1198),
        VN2CN5_sign => VN_sign_out(1199),
        codeword => codeword(199),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN200 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1205 downto 1200),
        Din0 => VN200_in0,
        Din1 => VN200_in1,
        Din2 => VN200_in2,
        Din3 => VN200_in3,
        Din4 => VN200_in4,
        Din5 => VN200_in5,
        VN2CN0_bit => VN_data_out(1200),
        VN2CN1_bit => VN_data_out(1201),
        VN2CN2_bit => VN_data_out(1202),
        VN2CN3_bit => VN_data_out(1203),
        VN2CN4_bit => VN_data_out(1204),
        VN2CN5_bit => VN_data_out(1205),
        VN2CN0_sign => VN_sign_out(1200),
        VN2CN1_sign => VN_sign_out(1201),
        VN2CN2_sign => VN_sign_out(1202),
        VN2CN3_sign => VN_sign_out(1203),
        VN2CN4_sign => VN_sign_out(1204),
        VN2CN5_sign => VN_sign_out(1205),
        codeword => codeword(200),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN201 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1211 downto 1206),
        Din0 => VN201_in0,
        Din1 => VN201_in1,
        Din2 => VN201_in2,
        Din3 => VN201_in3,
        Din4 => VN201_in4,
        Din5 => VN201_in5,
        VN2CN0_bit => VN_data_out(1206),
        VN2CN1_bit => VN_data_out(1207),
        VN2CN2_bit => VN_data_out(1208),
        VN2CN3_bit => VN_data_out(1209),
        VN2CN4_bit => VN_data_out(1210),
        VN2CN5_bit => VN_data_out(1211),
        VN2CN0_sign => VN_sign_out(1206),
        VN2CN1_sign => VN_sign_out(1207),
        VN2CN2_sign => VN_sign_out(1208),
        VN2CN3_sign => VN_sign_out(1209),
        VN2CN4_sign => VN_sign_out(1210),
        VN2CN5_sign => VN_sign_out(1211),
        codeword => codeword(201),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN202 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1217 downto 1212),
        Din0 => VN202_in0,
        Din1 => VN202_in1,
        Din2 => VN202_in2,
        Din3 => VN202_in3,
        Din4 => VN202_in4,
        Din5 => VN202_in5,
        VN2CN0_bit => VN_data_out(1212),
        VN2CN1_bit => VN_data_out(1213),
        VN2CN2_bit => VN_data_out(1214),
        VN2CN3_bit => VN_data_out(1215),
        VN2CN4_bit => VN_data_out(1216),
        VN2CN5_bit => VN_data_out(1217),
        VN2CN0_sign => VN_sign_out(1212),
        VN2CN1_sign => VN_sign_out(1213),
        VN2CN2_sign => VN_sign_out(1214),
        VN2CN3_sign => VN_sign_out(1215),
        VN2CN4_sign => VN_sign_out(1216),
        VN2CN5_sign => VN_sign_out(1217),
        codeword => codeword(202),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN203 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1223 downto 1218),
        Din0 => VN203_in0,
        Din1 => VN203_in1,
        Din2 => VN203_in2,
        Din3 => VN203_in3,
        Din4 => VN203_in4,
        Din5 => VN203_in5,
        VN2CN0_bit => VN_data_out(1218),
        VN2CN1_bit => VN_data_out(1219),
        VN2CN2_bit => VN_data_out(1220),
        VN2CN3_bit => VN_data_out(1221),
        VN2CN4_bit => VN_data_out(1222),
        VN2CN5_bit => VN_data_out(1223),
        VN2CN0_sign => VN_sign_out(1218),
        VN2CN1_sign => VN_sign_out(1219),
        VN2CN2_sign => VN_sign_out(1220),
        VN2CN3_sign => VN_sign_out(1221),
        VN2CN4_sign => VN_sign_out(1222),
        VN2CN5_sign => VN_sign_out(1223),
        codeword => codeword(203),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN204 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1229 downto 1224),
        Din0 => VN204_in0,
        Din1 => VN204_in1,
        Din2 => VN204_in2,
        Din3 => VN204_in3,
        Din4 => VN204_in4,
        Din5 => VN204_in5,
        VN2CN0_bit => VN_data_out(1224),
        VN2CN1_bit => VN_data_out(1225),
        VN2CN2_bit => VN_data_out(1226),
        VN2CN3_bit => VN_data_out(1227),
        VN2CN4_bit => VN_data_out(1228),
        VN2CN5_bit => VN_data_out(1229),
        VN2CN0_sign => VN_sign_out(1224),
        VN2CN1_sign => VN_sign_out(1225),
        VN2CN2_sign => VN_sign_out(1226),
        VN2CN3_sign => VN_sign_out(1227),
        VN2CN4_sign => VN_sign_out(1228),
        VN2CN5_sign => VN_sign_out(1229),
        codeword => codeword(204),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN205 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1235 downto 1230),
        Din0 => VN205_in0,
        Din1 => VN205_in1,
        Din2 => VN205_in2,
        Din3 => VN205_in3,
        Din4 => VN205_in4,
        Din5 => VN205_in5,
        VN2CN0_bit => VN_data_out(1230),
        VN2CN1_bit => VN_data_out(1231),
        VN2CN2_bit => VN_data_out(1232),
        VN2CN3_bit => VN_data_out(1233),
        VN2CN4_bit => VN_data_out(1234),
        VN2CN5_bit => VN_data_out(1235),
        VN2CN0_sign => VN_sign_out(1230),
        VN2CN1_sign => VN_sign_out(1231),
        VN2CN2_sign => VN_sign_out(1232),
        VN2CN3_sign => VN_sign_out(1233),
        VN2CN4_sign => VN_sign_out(1234),
        VN2CN5_sign => VN_sign_out(1235),
        codeword => codeword(205),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN206 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1241 downto 1236),
        Din0 => VN206_in0,
        Din1 => VN206_in1,
        Din2 => VN206_in2,
        Din3 => VN206_in3,
        Din4 => VN206_in4,
        Din5 => VN206_in5,
        VN2CN0_bit => VN_data_out(1236),
        VN2CN1_bit => VN_data_out(1237),
        VN2CN2_bit => VN_data_out(1238),
        VN2CN3_bit => VN_data_out(1239),
        VN2CN4_bit => VN_data_out(1240),
        VN2CN5_bit => VN_data_out(1241),
        VN2CN0_sign => VN_sign_out(1236),
        VN2CN1_sign => VN_sign_out(1237),
        VN2CN2_sign => VN_sign_out(1238),
        VN2CN3_sign => VN_sign_out(1239),
        VN2CN4_sign => VN_sign_out(1240),
        VN2CN5_sign => VN_sign_out(1241),
        codeword => codeword(206),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN207 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1247 downto 1242),
        Din0 => VN207_in0,
        Din1 => VN207_in1,
        Din2 => VN207_in2,
        Din3 => VN207_in3,
        Din4 => VN207_in4,
        Din5 => VN207_in5,
        VN2CN0_bit => VN_data_out(1242),
        VN2CN1_bit => VN_data_out(1243),
        VN2CN2_bit => VN_data_out(1244),
        VN2CN3_bit => VN_data_out(1245),
        VN2CN4_bit => VN_data_out(1246),
        VN2CN5_bit => VN_data_out(1247),
        VN2CN0_sign => VN_sign_out(1242),
        VN2CN1_sign => VN_sign_out(1243),
        VN2CN2_sign => VN_sign_out(1244),
        VN2CN3_sign => VN_sign_out(1245),
        VN2CN4_sign => VN_sign_out(1246),
        VN2CN5_sign => VN_sign_out(1247),
        codeword => codeword(207),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN208 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1253 downto 1248),
        Din0 => VN208_in0,
        Din1 => VN208_in1,
        Din2 => VN208_in2,
        Din3 => VN208_in3,
        Din4 => VN208_in4,
        Din5 => VN208_in5,
        VN2CN0_bit => VN_data_out(1248),
        VN2CN1_bit => VN_data_out(1249),
        VN2CN2_bit => VN_data_out(1250),
        VN2CN3_bit => VN_data_out(1251),
        VN2CN4_bit => VN_data_out(1252),
        VN2CN5_bit => VN_data_out(1253),
        VN2CN0_sign => VN_sign_out(1248),
        VN2CN1_sign => VN_sign_out(1249),
        VN2CN2_sign => VN_sign_out(1250),
        VN2CN3_sign => VN_sign_out(1251),
        VN2CN4_sign => VN_sign_out(1252),
        VN2CN5_sign => VN_sign_out(1253),
        codeword => codeword(208),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN209 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1259 downto 1254),
        Din0 => VN209_in0,
        Din1 => VN209_in1,
        Din2 => VN209_in2,
        Din3 => VN209_in3,
        Din4 => VN209_in4,
        Din5 => VN209_in5,
        VN2CN0_bit => VN_data_out(1254),
        VN2CN1_bit => VN_data_out(1255),
        VN2CN2_bit => VN_data_out(1256),
        VN2CN3_bit => VN_data_out(1257),
        VN2CN4_bit => VN_data_out(1258),
        VN2CN5_bit => VN_data_out(1259),
        VN2CN0_sign => VN_sign_out(1254),
        VN2CN1_sign => VN_sign_out(1255),
        VN2CN2_sign => VN_sign_out(1256),
        VN2CN3_sign => VN_sign_out(1257),
        VN2CN4_sign => VN_sign_out(1258),
        VN2CN5_sign => VN_sign_out(1259),
        codeword => codeword(209),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN210 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1265 downto 1260),
        Din0 => VN210_in0,
        Din1 => VN210_in1,
        Din2 => VN210_in2,
        Din3 => VN210_in3,
        Din4 => VN210_in4,
        Din5 => VN210_in5,
        VN2CN0_bit => VN_data_out(1260),
        VN2CN1_bit => VN_data_out(1261),
        VN2CN2_bit => VN_data_out(1262),
        VN2CN3_bit => VN_data_out(1263),
        VN2CN4_bit => VN_data_out(1264),
        VN2CN5_bit => VN_data_out(1265),
        VN2CN0_sign => VN_sign_out(1260),
        VN2CN1_sign => VN_sign_out(1261),
        VN2CN2_sign => VN_sign_out(1262),
        VN2CN3_sign => VN_sign_out(1263),
        VN2CN4_sign => VN_sign_out(1264),
        VN2CN5_sign => VN_sign_out(1265),
        codeword => codeword(210),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN211 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1271 downto 1266),
        Din0 => VN211_in0,
        Din1 => VN211_in1,
        Din2 => VN211_in2,
        Din3 => VN211_in3,
        Din4 => VN211_in4,
        Din5 => VN211_in5,
        VN2CN0_bit => VN_data_out(1266),
        VN2CN1_bit => VN_data_out(1267),
        VN2CN2_bit => VN_data_out(1268),
        VN2CN3_bit => VN_data_out(1269),
        VN2CN4_bit => VN_data_out(1270),
        VN2CN5_bit => VN_data_out(1271),
        VN2CN0_sign => VN_sign_out(1266),
        VN2CN1_sign => VN_sign_out(1267),
        VN2CN2_sign => VN_sign_out(1268),
        VN2CN3_sign => VN_sign_out(1269),
        VN2CN4_sign => VN_sign_out(1270),
        VN2CN5_sign => VN_sign_out(1271),
        codeword => codeword(211),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN212 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1277 downto 1272),
        Din0 => VN212_in0,
        Din1 => VN212_in1,
        Din2 => VN212_in2,
        Din3 => VN212_in3,
        Din4 => VN212_in4,
        Din5 => VN212_in5,
        VN2CN0_bit => VN_data_out(1272),
        VN2CN1_bit => VN_data_out(1273),
        VN2CN2_bit => VN_data_out(1274),
        VN2CN3_bit => VN_data_out(1275),
        VN2CN4_bit => VN_data_out(1276),
        VN2CN5_bit => VN_data_out(1277),
        VN2CN0_sign => VN_sign_out(1272),
        VN2CN1_sign => VN_sign_out(1273),
        VN2CN2_sign => VN_sign_out(1274),
        VN2CN3_sign => VN_sign_out(1275),
        VN2CN4_sign => VN_sign_out(1276),
        VN2CN5_sign => VN_sign_out(1277),
        codeword => codeword(212),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN213 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1283 downto 1278),
        Din0 => VN213_in0,
        Din1 => VN213_in1,
        Din2 => VN213_in2,
        Din3 => VN213_in3,
        Din4 => VN213_in4,
        Din5 => VN213_in5,
        VN2CN0_bit => VN_data_out(1278),
        VN2CN1_bit => VN_data_out(1279),
        VN2CN2_bit => VN_data_out(1280),
        VN2CN3_bit => VN_data_out(1281),
        VN2CN4_bit => VN_data_out(1282),
        VN2CN5_bit => VN_data_out(1283),
        VN2CN0_sign => VN_sign_out(1278),
        VN2CN1_sign => VN_sign_out(1279),
        VN2CN2_sign => VN_sign_out(1280),
        VN2CN3_sign => VN_sign_out(1281),
        VN2CN4_sign => VN_sign_out(1282),
        VN2CN5_sign => VN_sign_out(1283),
        codeword => codeword(213),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN214 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1289 downto 1284),
        Din0 => VN214_in0,
        Din1 => VN214_in1,
        Din2 => VN214_in2,
        Din3 => VN214_in3,
        Din4 => VN214_in4,
        Din5 => VN214_in5,
        VN2CN0_bit => VN_data_out(1284),
        VN2CN1_bit => VN_data_out(1285),
        VN2CN2_bit => VN_data_out(1286),
        VN2CN3_bit => VN_data_out(1287),
        VN2CN4_bit => VN_data_out(1288),
        VN2CN5_bit => VN_data_out(1289),
        VN2CN0_sign => VN_sign_out(1284),
        VN2CN1_sign => VN_sign_out(1285),
        VN2CN2_sign => VN_sign_out(1286),
        VN2CN3_sign => VN_sign_out(1287),
        VN2CN4_sign => VN_sign_out(1288),
        VN2CN5_sign => VN_sign_out(1289),
        codeword => codeword(214),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN215 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1295 downto 1290),
        Din0 => VN215_in0,
        Din1 => VN215_in1,
        Din2 => VN215_in2,
        Din3 => VN215_in3,
        Din4 => VN215_in4,
        Din5 => VN215_in5,
        VN2CN0_bit => VN_data_out(1290),
        VN2CN1_bit => VN_data_out(1291),
        VN2CN2_bit => VN_data_out(1292),
        VN2CN3_bit => VN_data_out(1293),
        VN2CN4_bit => VN_data_out(1294),
        VN2CN5_bit => VN_data_out(1295),
        VN2CN0_sign => VN_sign_out(1290),
        VN2CN1_sign => VN_sign_out(1291),
        VN2CN2_sign => VN_sign_out(1292),
        VN2CN3_sign => VN_sign_out(1293),
        VN2CN4_sign => VN_sign_out(1294),
        VN2CN5_sign => VN_sign_out(1295),
        codeword => codeword(215),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN216 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1301 downto 1296),
        Din0 => VN216_in0,
        Din1 => VN216_in1,
        Din2 => VN216_in2,
        Din3 => VN216_in3,
        Din4 => VN216_in4,
        Din5 => VN216_in5,
        VN2CN0_bit => VN_data_out(1296),
        VN2CN1_bit => VN_data_out(1297),
        VN2CN2_bit => VN_data_out(1298),
        VN2CN3_bit => VN_data_out(1299),
        VN2CN4_bit => VN_data_out(1300),
        VN2CN5_bit => VN_data_out(1301),
        VN2CN0_sign => VN_sign_out(1296),
        VN2CN1_sign => VN_sign_out(1297),
        VN2CN2_sign => VN_sign_out(1298),
        VN2CN3_sign => VN_sign_out(1299),
        VN2CN4_sign => VN_sign_out(1300),
        VN2CN5_sign => VN_sign_out(1301),
        codeword => codeword(216),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN217 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1307 downto 1302),
        Din0 => VN217_in0,
        Din1 => VN217_in1,
        Din2 => VN217_in2,
        Din3 => VN217_in3,
        Din4 => VN217_in4,
        Din5 => VN217_in5,
        VN2CN0_bit => VN_data_out(1302),
        VN2CN1_bit => VN_data_out(1303),
        VN2CN2_bit => VN_data_out(1304),
        VN2CN3_bit => VN_data_out(1305),
        VN2CN4_bit => VN_data_out(1306),
        VN2CN5_bit => VN_data_out(1307),
        VN2CN0_sign => VN_sign_out(1302),
        VN2CN1_sign => VN_sign_out(1303),
        VN2CN2_sign => VN_sign_out(1304),
        VN2CN3_sign => VN_sign_out(1305),
        VN2CN4_sign => VN_sign_out(1306),
        VN2CN5_sign => VN_sign_out(1307),
        codeword => codeword(217),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN218 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1313 downto 1308),
        Din0 => VN218_in0,
        Din1 => VN218_in1,
        Din2 => VN218_in2,
        Din3 => VN218_in3,
        Din4 => VN218_in4,
        Din5 => VN218_in5,
        VN2CN0_bit => VN_data_out(1308),
        VN2CN1_bit => VN_data_out(1309),
        VN2CN2_bit => VN_data_out(1310),
        VN2CN3_bit => VN_data_out(1311),
        VN2CN4_bit => VN_data_out(1312),
        VN2CN5_bit => VN_data_out(1313),
        VN2CN0_sign => VN_sign_out(1308),
        VN2CN1_sign => VN_sign_out(1309),
        VN2CN2_sign => VN_sign_out(1310),
        VN2CN3_sign => VN_sign_out(1311),
        VN2CN4_sign => VN_sign_out(1312),
        VN2CN5_sign => VN_sign_out(1313),
        codeword => codeword(218),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN219 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1319 downto 1314),
        Din0 => VN219_in0,
        Din1 => VN219_in1,
        Din2 => VN219_in2,
        Din3 => VN219_in3,
        Din4 => VN219_in4,
        Din5 => VN219_in5,
        VN2CN0_bit => VN_data_out(1314),
        VN2CN1_bit => VN_data_out(1315),
        VN2CN2_bit => VN_data_out(1316),
        VN2CN3_bit => VN_data_out(1317),
        VN2CN4_bit => VN_data_out(1318),
        VN2CN5_bit => VN_data_out(1319),
        VN2CN0_sign => VN_sign_out(1314),
        VN2CN1_sign => VN_sign_out(1315),
        VN2CN2_sign => VN_sign_out(1316),
        VN2CN3_sign => VN_sign_out(1317),
        VN2CN4_sign => VN_sign_out(1318),
        VN2CN5_sign => VN_sign_out(1319),
        codeword => codeword(219),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN220 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1325 downto 1320),
        Din0 => VN220_in0,
        Din1 => VN220_in1,
        Din2 => VN220_in2,
        Din3 => VN220_in3,
        Din4 => VN220_in4,
        Din5 => VN220_in5,
        VN2CN0_bit => VN_data_out(1320),
        VN2CN1_bit => VN_data_out(1321),
        VN2CN2_bit => VN_data_out(1322),
        VN2CN3_bit => VN_data_out(1323),
        VN2CN4_bit => VN_data_out(1324),
        VN2CN5_bit => VN_data_out(1325),
        VN2CN0_sign => VN_sign_out(1320),
        VN2CN1_sign => VN_sign_out(1321),
        VN2CN2_sign => VN_sign_out(1322),
        VN2CN3_sign => VN_sign_out(1323),
        VN2CN4_sign => VN_sign_out(1324),
        VN2CN5_sign => VN_sign_out(1325),
        codeword => codeword(220),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN221 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1331 downto 1326),
        Din0 => VN221_in0,
        Din1 => VN221_in1,
        Din2 => VN221_in2,
        Din3 => VN221_in3,
        Din4 => VN221_in4,
        Din5 => VN221_in5,
        VN2CN0_bit => VN_data_out(1326),
        VN2CN1_bit => VN_data_out(1327),
        VN2CN2_bit => VN_data_out(1328),
        VN2CN3_bit => VN_data_out(1329),
        VN2CN4_bit => VN_data_out(1330),
        VN2CN5_bit => VN_data_out(1331),
        VN2CN0_sign => VN_sign_out(1326),
        VN2CN1_sign => VN_sign_out(1327),
        VN2CN2_sign => VN_sign_out(1328),
        VN2CN3_sign => VN_sign_out(1329),
        VN2CN4_sign => VN_sign_out(1330),
        VN2CN5_sign => VN_sign_out(1331),
        codeword => codeword(221),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN222 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1337 downto 1332),
        Din0 => VN222_in0,
        Din1 => VN222_in1,
        Din2 => VN222_in2,
        Din3 => VN222_in3,
        Din4 => VN222_in4,
        Din5 => VN222_in5,
        VN2CN0_bit => VN_data_out(1332),
        VN2CN1_bit => VN_data_out(1333),
        VN2CN2_bit => VN_data_out(1334),
        VN2CN3_bit => VN_data_out(1335),
        VN2CN4_bit => VN_data_out(1336),
        VN2CN5_bit => VN_data_out(1337),
        VN2CN0_sign => VN_sign_out(1332),
        VN2CN1_sign => VN_sign_out(1333),
        VN2CN2_sign => VN_sign_out(1334),
        VN2CN3_sign => VN_sign_out(1335),
        VN2CN4_sign => VN_sign_out(1336),
        VN2CN5_sign => VN_sign_out(1337),
        codeword => codeword(222),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN223 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1343 downto 1338),
        Din0 => VN223_in0,
        Din1 => VN223_in1,
        Din2 => VN223_in2,
        Din3 => VN223_in3,
        Din4 => VN223_in4,
        Din5 => VN223_in5,
        VN2CN0_bit => VN_data_out(1338),
        VN2CN1_bit => VN_data_out(1339),
        VN2CN2_bit => VN_data_out(1340),
        VN2CN3_bit => VN_data_out(1341),
        VN2CN4_bit => VN_data_out(1342),
        VN2CN5_bit => VN_data_out(1343),
        VN2CN0_sign => VN_sign_out(1338),
        VN2CN1_sign => VN_sign_out(1339),
        VN2CN2_sign => VN_sign_out(1340),
        VN2CN3_sign => VN_sign_out(1341),
        VN2CN4_sign => VN_sign_out(1342),
        VN2CN5_sign => VN_sign_out(1343),
        codeword => codeword(223),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN224 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1349 downto 1344),
        Din0 => VN224_in0,
        Din1 => VN224_in1,
        Din2 => VN224_in2,
        Din3 => VN224_in3,
        Din4 => VN224_in4,
        Din5 => VN224_in5,
        VN2CN0_bit => VN_data_out(1344),
        VN2CN1_bit => VN_data_out(1345),
        VN2CN2_bit => VN_data_out(1346),
        VN2CN3_bit => VN_data_out(1347),
        VN2CN4_bit => VN_data_out(1348),
        VN2CN5_bit => VN_data_out(1349),
        VN2CN0_sign => VN_sign_out(1344),
        VN2CN1_sign => VN_sign_out(1345),
        VN2CN2_sign => VN_sign_out(1346),
        VN2CN3_sign => VN_sign_out(1347),
        VN2CN4_sign => VN_sign_out(1348),
        VN2CN5_sign => VN_sign_out(1349),
        codeword => codeword(224),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN225 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1355 downto 1350),
        Din0 => VN225_in0,
        Din1 => VN225_in1,
        Din2 => VN225_in2,
        Din3 => VN225_in3,
        Din4 => VN225_in4,
        Din5 => VN225_in5,
        VN2CN0_bit => VN_data_out(1350),
        VN2CN1_bit => VN_data_out(1351),
        VN2CN2_bit => VN_data_out(1352),
        VN2CN3_bit => VN_data_out(1353),
        VN2CN4_bit => VN_data_out(1354),
        VN2CN5_bit => VN_data_out(1355),
        VN2CN0_sign => VN_sign_out(1350),
        VN2CN1_sign => VN_sign_out(1351),
        VN2CN2_sign => VN_sign_out(1352),
        VN2CN3_sign => VN_sign_out(1353),
        VN2CN4_sign => VN_sign_out(1354),
        VN2CN5_sign => VN_sign_out(1355),
        codeword => codeword(225),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN226 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1361 downto 1356),
        Din0 => VN226_in0,
        Din1 => VN226_in1,
        Din2 => VN226_in2,
        Din3 => VN226_in3,
        Din4 => VN226_in4,
        Din5 => VN226_in5,
        VN2CN0_bit => VN_data_out(1356),
        VN2CN1_bit => VN_data_out(1357),
        VN2CN2_bit => VN_data_out(1358),
        VN2CN3_bit => VN_data_out(1359),
        VN2CN4_bit => VN_data_out(1360),
        VN2CN5_bit => VN_data_out(1361),
        VN2CN0_sign => VN_sign_out(1356),
        VN2CN1_sign => VN_sign_out(1357),
        VN2CN2_sign => VN_sign_out(1358),
        VN2CN3_sign => VN_sign_out(1359),
        VN2CN4_sign => VN_sign_out(1360),
        VN2CN5_sign => VN_sign_out(1361),
        codeword => codeword(226),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN227 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1367 downto 1362),
        Din0 => VN227_in0,
        Din1 => VN227_in1,
        Din2 => VN227_in2,
        Din3 => VN227_in3,
        Din4 => VN227_in4,
        Din5 => VN227_in5,
        VN2CN0_bit => VN_data_out(1362),
        VN2CN1_bit => VN_data_out(1363),
        VN2CN2_bit => VN_data_out(1364),
        VN2CN3_bit => VN_data_out(1365),
        VN2CN4_bit => VN_data_out(1366),
        VN2CN5_bit => VN_data_out(1367),
        VN2CN0_sign => VN_sign_out(1362),
        VN2CN1_sign => VN_sign_out(1363),
        VN2CN2_sign => VN_sign_out(1364),
        VN2CN3_sign => VN_sign_out(1365),
        VN2CN4_sign => VN_sign_out(1366),
        VN2CN5_sign => VN_sign_out(1367),
        codeword => codeword(227),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN228 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1373 downto 1368),
        Din0 => VN228_in0,
        Din1 => VN228_in1,
        Din2 => VN228_in2,
        Din3 => VN228_in3,
        Din4 => VN228_in4,
        Din5 => VN228_in5,
        VN2CN0_bit => VN_data_out(1368),
        VN2CN1_bit => VN_data_out(1369),
        VN2CN2_bit => VN_data_out(1370),
        VN2CN3_bit => VN_data_out(1371),
        VN2CN4_bit => VN_data_out(1372),
        VN2CN5_bit => VN_data_out(1373),
        VN2CN0_sign => VN_sign_out(1368),
        VN2CN1_sign => VN_sign_out(1369),
        VN2CN2_sign => VN_sign_out(1370),
        VN2CN3_sign => VN_sign_out(1371),
        VN2CN4_sign => VN_sign_out(1372),
        VN2CN5_sign => VN_sign_out(1373),
        codeword => codeword(228),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN229 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1379 downto 1374),
        Din0 => VN229_in0,
        Din1 => VN229_in1,
        Din2 => VN229_in2,
        Din3 => VN229_in3,
        Din4 => VN229_in4,
        Din5 => VN229_in5,
        VN2CN0_bit => VN_data_out(1374),
        VN2CN1_bit => VN_data_out(1375),
        VN2CN2_bit => VN_data_out(1376),
        VN2CN3_bit => VN_data_out(1377),
        VN2CN4_bit => VN_data_out(1378),
        VN2CN5_bit => VN_data_out(1379),
        VN2CN0_sign => VN_sign_out(1374),
        VN2CN1_sign => VN_sign_out(1375),
        VN2CN2_sign => VN_sign_out(1376),
        VN2CN3_sign => VN_sign_out(1377),
        VN2CN4_sign => VN_sign_out(1378),
        VN2CN5_sign => VN_sign_out(1379),
        codeword => codeword(229),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN230 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1385 downto 1380),
        Din0 => VN230_in0,
        Din1 => VN230_in1,
        Din2 => VN230_in2,
        Din3 => VN230_in3,
        Din4 => VN230_in4,
        Din5 => VN230_in5,
        VN2CN0_bit => VN_data_out(1380),
        VN2CN1_bit => VN_data_out(1381),
        VN2CN2_bit => VN_data_out(1382),
        VN2CN3_bit => VN_data_out(1383),
        VN2CN4_bit => VN_data_out(1384),
        VN2CN5_bit => VN_data_out(1385),
        VN2CN0_sign => VN_sign_out(1380),
        VN2CN1_sign => VN_sign_out(1381),
        VN2CN2_sign => VN_sign_out(1382),
        VN2CN3_sign => VN_sign_out(1383),
        VN2CN4_sign => VN_sign_out(1384),
        VN2CN5_sign => VN_sign_out(1385),
        codeword => codeword(230),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN231 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1391 downto 1386),
        Din0 => VN231_in0,
        Din1 => VN231_in1,
        Din2 => VN231_in2,
        Din3 => VN231_in3,
        Din4 => VN231_in4,
        Din5 => VN231_in5,
        VN2CN0_bit => VN_data_out(1386),
        VN2CN1_bit => VN_data_out(1387),
        VN2CN2_bit => VN_data_out(1388),
        VN2CN3_bit => VN_data_out(1389),
        VN2CN4_bit => VN_data_out(1390),
        VN2CN5_bit => VN_data_out(1391),
        VN2CN0_sign => VN_sign_out(1386),
        VN2CN1_sign => VN_sign_out(1387),
        VN2CN2_sign => VN_sign_out(1388),
        VN2CN3_sign => VN_sign_out(1389),
        VN2CN4_sign => VN_sign_out(1390),
        VN2CN5_sign => VN_sign_out(1391),
        codeword => codeword(231),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN232 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1397 downto 1392),
        Din0 => VN232_in0,
        Din1 => VN232_in1,
        Din2 => VN232_in2,
        Din3 => VN232_in3,
        Din4 => VN232_in4,
        Din5 => VN232_in5,
        VN2CN0_bit => VN_data_out(1392),
        VN2CN1_bit => VN_data_out(1393),
        VN2CN2_bit => VN_data_out(1394),
        VN2CN3_bit => VN_data_out(1395),
        VN2CN4_bit => VN_data_out(1396),
        VN2CN5_bit => VN_data_out(1397),
        VN2CN0_sign => VN_sign_out(1392),
        VN2CN1_sign => VN_sign_out(1393),
        VN2CN2_sign => VN_sign_out(1394),
        VN2CN3_sign => VN_sign_out(1395),
        VN2CN4_sign => VN_sign_out(1396),
        VN2CN5_sign => VN_sign_out(1397),
        codeword => codeword(232),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN233 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1403 downto 1398),
        Din0 => VN233_in0,
        Din1 => VN233_in1,
        Din2 => VN233_in2,
        Din3 => VN233_in3,
        Din4 => VN233_in4,
        Din5 => VN233_in5,
        VN2CN0_bit => VN_data_out(1398),
        VN2CN1_bit => VN_data_out(1399),
        VN2CN2_bit => VN_data_out(1400),
        VN2CN3_bit => VN_data_out(1401),
        VN2CN4_bit => VN_data_out(1402),
        VN2CN5_bit => VN_data_out(1403),
        VN2CN0_sign => VN_sign_out(1398),
        VN2CN1_sign => VN_sign_out(1399),
        VN2CN2_sign => VN_sign_out(1400),
        VN2CN3_sign => VN_sign_out(1401),
        VN2CN4_sign => VN_sign_out(1402),
        VN2CN5_sign => VN_sign_out(1403),
        codeword => codeword(233),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN234 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1409 downto 1404),
        Din0 => VN234_in0,
        Din1 => VN234_in1,
        Din2 => VN234_in2,
        Din3 => VN234_in3,
        Din4 => VN234_in4,
        Din5 => VN234_in5,
        VN2CN0_bit => VN_data_out(1404),
        VN2CN1_bit => VN_data_out(1405),
        VN2CN2_bit => VN_data_out(1406),
        VN2CN3_bit => VN_data_out(1407),
        VN2CN4_bit => VN_data_out(1408),
        VN2CN5_bit => VN_data_out(1409),
        VN2CN0_sign => VN_sign_out(1404),
        VN2CN1_sign => VN_sign_out(1405),
        VN2CN2_sign => VN_sign_out(1406),
        VN2CN3_sign => VN_sign_out(1407),
        VN2CN4_sign => VN_sign_out(1408),
        VN2CN5_sign => VN_sign_out(1409),
        codeword => codeword(234),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN235 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1415 downto 1410),
        Din0 => VN235_in0,
        Din1 => VN235_in1,
        Din2 => VN235_in2,
        Din3 => VN235_in3,
        Din4 => VN235_in4,
        Din5 => VN235_in5,
        VN2CN0_bit => VN_data_out(1410),
        VN2CN1_bit => VN_data_out(1411),
        VN2CN2_bit => VN_data_out(1412),
        VN2CN3_bit => VN_data_out(1413),
        VN2CN4_bit => VN_data_out(1414),
        VN2CN5_bit => VN_data_out(1415),
        VN2CN0_sign => VN_sign_out(1410),
        VN2CN1_sign => VN_sign_out(1411),
        VN2CN2_sign => VN_sign_out(1412),
        VN2CN3_sign => VN_sign_out(1413),
        VN2CN4_sign => VN_sign_out(1414),
        VN2CN5_sign => VN_sign_out(1415),
        codeword => codeword(235),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN236 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1421 downto 1416),
        Din0 => VN236_in0,
        Din1 => VN236_in1,
        Din2 => VN236_in2,
        Din3 => VN236_in3,
        Din4 => VN236_in4,
        Din5 => VN236_in5,
        VN2CN0_bit => VN_data_out(1416),
        VN2CN1_bit => VN_data_out(1417),
        VN2CN2_bit => VN_data_out(1418),
        VN2CN3_bit => VN_data_out(1419),
        VN2CN4_bit => VN_data_out(1420),
        VN2CN5_bit => VN_data_out(1421),
        VN2CN0_sign => VN_sign_out(1416),
        VN2CN1_sign => VN_sign_out(1417),
        VN2CN2_sign => VN_sign_out(1418),
        VN2CN3_sign => VN_sign_out(1419),
        VN2CN4_sign => VN_sign_out(1420),
        VN2CN5_sign => VN_sign_out(1421),
        codeword => codeword(236),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN237 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1427 downto 1422),
        Din0 => VN237_in0,
        Din1 => VN237_in1,
        Din2 => VN237_in2,
        Din3 => VN237_in3,
        Din4 => VN237_in4,
        Din5 => VN237_in5,
        VN2CN0_bit => VN_data_out(1422),
        VN2CN1_bit => VN_data_out(1423),
        VN2CN2_bit => VN_data_out(1424),
        VN2CN3_bit => VN_data_out(1425),
        VN2CN4_bit => VN_data_out(1426),
        VN2CN5_bit => VN_data_out(1427),
        VN2CN0_sign => VN_sign_out(1422),
        VN2CN1_sign => VN_sign_out(1423),
        VN2CN2_sign => VN_sign_out(1424),
        VN2CN3_sign => VN_sign_out(1425),
        VN2CN4_sign => VN_sign_out(1426),
        VN2CN5_sign => VN_sign_out(1427),
        codeword => codeword(237),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN238 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1433 downto 1428),
        Din0 => VN238_in0,
        Din1 => VN238_in1,
        Din2 => VN238_in2,
        Din3 => VN238_in3,
        Din4 => VN238_in4,
        Din5 => VN238_in5,
        VN2CN0_bit => VN_data_out(1428),
        VN2CN1_bit => VN_data_out(1429),
        VN2CN2_bit => VN_data_out(1430),
        VN2CN3_bit => VN_data_out(1431),
        VN2CN4_bit => VN_data_out(1432),
        VN2CN5_bit => VN_data_out(1433),
        VN2CN0_sign => VN_sign_out(1428),
        VN2CN1_sign => VN_sign_out(1429),
        VN2CN2_sign => VN_sign_out(1430),
        VN2CN3_sign => VN_sign_out(1431),
        VN2CN4_sign => VN_sign_out(1432),
        VN2CN5_sign => VN_sign_out(1433),
        codeword => codeword(238),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN239 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1439 downto 1434),
        Din0 => VN239_in0,
        Din1 => VN239_in1,
        Din2 => VN239_in2,
        Din3 => VN239_in3,
        Din4 => VN239_in4,
        Din5 => VN239_in5,
        VN2CN0_bit => VN_data_out(1434),
        VN2CN1_bit => VN_data_out(1435),
        VN2CN2_bit => VN_data_out(1436),
        VN2CN3_bit => VN_data_out(1437),
        VN2CN4_bit => VN_data_out(1438),
        VN2CN5_bit => VN_data_out(1439),
        VN2CN0_sign => VN_sign_out(1434),
        VN2CN1_sign => VN_sign_out(1435),
        VN2CN2_sign => VN_sign_out(1436),
        VN2CN3_sign => VN_sign_out(1437),
        VN2CN4_sign => VN_sign_out(1438),
        VN2CN5_sign => VN_sign_out(1439),
        codeword => codeword(239),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN240 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1445 downto 1440),
        Din0 => VN240_in0,
        Din1 => VN240_in1,
        Din2 => VN240_in2,
        Din3 => VN240_in3,
        Din4 => VN240_in4,
        Din5 => VN240_in5,
        VN2CN0_bit => VN_data_out(1440),
        VN2CN1_bit => VN_data_out(1441),
        VN2CN2_bit => VN_data_out(1442),
        VN2CN3_bit => VN_data_out(1443),
        VN2CN4_bit => VN_data_out(1444),
        VN2CN5_bit => VN_data_out(1445),
        VN2CN0_sign => VN_sign_out(1440),
        VN2CN1_sign => VN_sign_out(1441),
        VN2CN2_sign => VN_sign_out(1442),
        VN2CN3_sign => VN_sign_out(1443),
        VN2CN4_sign => VN_sign_out(1444),
        VN2CN5_sign => VN_sign_out(1445),
        codeword => codeword(240),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN241 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1451 downto 1446),
        Din0 => VN241_in0,
        Din1 => VN241_in1,
        Din2 => VN241_in2,
        Din3 => VN241_in3,
        Din4 => VN241_in4,
        Din5 => VN241_in5,
        VN2CN0_bit => VN_data_out(1446),
        VN2CN1_bit => VN_data_out(1447),
        VN2CN2_bit => VN_data_out(1448),
        VN2CN3_bit => VN_data_out(1449),
        VN2CN4_bit => VN_data_out(1450),
        VN2CN5_bit => VN_data_out(1451),
        VN2CN0_sign => VN_sign_out(1446),
        VN2CN1_sign => VN_sign_out(1447),
        VN2CN2_sign => VN_sign_out(1448),
        VN2CN3_sign => VN_sign_out(1449),
        VN2CN4_sign => VN_sign_out(1450),
        VN2CN5_sign => VN_sign_out(1451),
        codeword => codeword(241),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN242 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1457 downto 1452),
        Din0 => VN242_in0,
        Din1 => VN242_in1,
        Din2 => VN242_in2,
        Din3 => VN242_in3,
        Din4 => VN242_in4,
        Din5 => VN242_in5,
        VN2CN0_bit => VN_data_out(1452),
        VN2CN1_bit => VN_data_out(1453),
        VN2CN2_bit => VN_data_out(1454),
        VN2CN3_bit => VN_data_out(1455),
        VN2CN4_bit => VN_data_out(1456),
        VN2CN5_bit => VN_data_out(1457),
        VN2CN0_sign => VN_sign_out(1452),
        VN2CN1_sign => VN_sign_out(1453),
        VN2CN2_sign => VN_sign_out(1454),
        VN2CN3_sign => VN_sign_out(1455),
        VN2CN4_sign => VN_sign_out(1456),
        VN2CN5_sign => VN_sign_out(1457),
        codeword => codeword(242),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN243 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1463 downto 1458),
        Din0 => VN243_in0,
        Din1 => VN243_in1,
        Din2 => VN243_in2,
        Din3 => VN243_in3,
        Din4 => VN243_in4,
        Din5 => VN243_in5,
        VN2CN0_bit => VN_data_out(1458),
        VN2CN1_bit => VN_data_out(1459),
        VN2CN2_bit => VN_data_out(1460),
        VN2CN3_bit => VN_data_out(1461),
        VN2CN4_bit => VN_data_out(1462),
        VN2CN5_bit => VN_data_out(1463),
        VN2CN0_sign => VN_sign_out(1458),
        VN2CN1_sign => VN_sign_out(1459),
        VN2CN2_sign => VN_sign_out(1460),
        VN2CN3_sign => VN_sign_out(1461),
        VN2CN4_sign => VN_sign_out(1462),
        VN2CN5_sign => VN_sign_out(1463),
        codeword => codeword(243),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN244 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1469 downto 1464),
        Din0 => VN244_in0,
        Din1 => VN244_in1,
        Din2 => VN244_in2,
        Din3 => VN244_in3,
        Din4 => VN244_in4,
        Din5 => VN244_in5,
        VN2CN0_bit => VN_data_out(1464),
        VN2CN1_bit => VN_data_out(1465),
        VN2CN2_bit => VN_data_out(1466),
        VN2CN3_bit => VN_data_out(1467),
        VN2CN4_bit => VN_data_out(1468),
        VN2CN5_bit => VN_data_out(1469),
        VN2CN0_sign => VN_sign_out(1464),
        VN2CN1_sign => VN_sign_out(1465),
        VN2CN2_sign => VN_sign_out(1466),
        VN2CN3_sign => VN_sign_out(1467),
        VN2CN4_sign => VN_sign_out(1468),
        VN2CN5_sign => VN_sign_out(1469),
        codeword => codeword(244),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN245 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1475 downto 1470),
        Din0 => VN245_in0,
        Din1 => VN245_in1,
        Din2 => VN245_in2,
        Din3 => VN245_in3,
        Din4 => VN245_in4,
        Din5 => VN245_in5,
        VN2CN0_bit => VN_data_out(1470),
        VN2CN1_bit => VN_data_out(1471),
        VN2CN2_bit => VN_data_out(1472),
        VN2CN3_bit => VN_data_out(1473),
        VN2CN4_bit => VN_data_out(1474),
        VN2CN5_bit => VN_data_out(1475),
        VN2CN0_sign => VN_sign_out(1470),
        VN2CN1_sign => VN_sign_out(1471),
        VN2CN2_sign => VN_sign_out(1472),
        VN2CN3_sign => VN_sign_out(1473),
        VN2CN4_sign => VN_sign_out(1474),
        VN2CN5_sign => VN_sign_out(1475),
        codeword => codeword(245),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN246 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1481 downto 1476),
        Din0 => VN246_in0,
        Din1 => VN246_in1,
        Din2 => VN246_in2,
        Din3 => VN246_in3,
        Din4 => VN246_in4,
        Din5 => VN246_in5,
        VN2CN0_bit => VN_data_out(1476),
        VN2CN1_bit => VN_data_out(1477),
        VN2CN2_bit => VN_data_out(1478),
        VN2CN3_bit => VN_data_out(1479),
        VN2CN4_bit => VN_data_out(1480),
        VN2CN5_bit => VN_data_out(1481),
        VN2CN0_sign => VN_sign_out(1476),
        VN2CN1_sign => VN_sign_out(1477),
        VN2CN2_sign => VN_sign_out(1478),
        VN2CN3_sign => VN_sign_out(1479),
        VN2CN4_sign => VN_sign_out(1480),
        VN2CN5_sign => VN_sign_out(1481),
        codeword => codeword(246),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN247 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1487 downto 1482),
        Din0 => VN247_in0,
        Din1 => VN247_in1,
        Din2 => VN247_in2,
        Din3 => VN247_in3,
        Din4 => VN247_in4,
        Din5 => VN247_in5,
        VN2CN0_bit => VN_data_out(1482),
        VN2CN1_bit => VN_data_out(1483),
        VN2CN2_bit => VN_data_out(1484),
        VN2CN3_bit => VN_data_out(1485),
        VN2CN4_bit => VN_data_out(1486),
        VN2CN5_bit => VN_data_out(1487),
        VN2CN0_sign => VN_sign_out(1482),
        VN2CN1_sign => VN_sign_out(1483),
        VN2CN2_sign => VN_sign_out(1484),
        VN2CN3_sign => VN_sign_out(1485),
        VN2CN4_sign => VN_sign_out(1486),
        VN2CN5_sign => VN_sign_out(1487),
        codeword => codeword(247),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN248 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1493 downto 1488),
        Din0 => VN248_in0,
        Din1 => VN248_in1,
        Din2 => VN248_in2,
        Din3 => VN248_in3,
        Din4 => VN248_in4,
        Din5 => VN248_in5,
        VN2CN0_bit => VN_data_out(1488),
        VN2CN1_bit => VN_data_out(1489),
        VN2CN2_bit => VN_data_out(1490),
        VN2CN3_bit => VN_data_out(1491),
        VN2CN4_bit => VN_data_out(1492),
        VN2CN5_bit => VN_data_out(1493),
        VN2CN0_sign => VN_sign_out(1488),
        VN2CN1_sign => VN_sign_out(1489),
        VN2CN2_sign => VN_sign_out(1490),
        VN2CN3_sign => VN_sign_out(1491),
        VN2CN4_sign => VN_sign_out(1492),
        VN2CN5_sign => VN_sign_out(1493),
        codeword => codeword(248),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN249 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1499 downto 1494),
        Din0 => VN249_in0,
        Din1 => VN249_in1,
        Din2 => VN249_in2,
        Din3 => VN249_in3,
        Din4 => VN249_in4,
        Din5 => VN249_in5,
        VN2CN0_bit => VN_data_out(1494),
        VN2CN1_bit => VN_data_out(1495),
        VN2CN2_bit => VN_data_out(1496),
        VN2CN3_bit => VN_data_out(1497),
        VN2CN4_bit => VN_data_out(1498),
        VN2CN5_bit => VN_data_out(1499),
        VN2CN0_sign => VN_sign_out(1494),
        VN2CN1_sign => VN_sign_out(1495),
        VN2CN2_sign => VN_sign_out(1496),
        VN2CN3_sign => VN_sign_out(1497),
        VN2CN4_sign => VN_sign_out(1498),
        VN2CN5_sign => VN_sign_out(1499),
        codeword => codeword(249),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN250 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1505 downto 1500),
        Din0 => VN250_in0,
        Din1 => VN250_in1,
        Din2 => VN250_in2,
        Din3 => VN250_in3,
        Din4 => VN250_in4,
        Din5 => VN250_in5,
        VN2CN0_bit => VN_data_out(1500),
        VN2CN1_bit => VN_data_out(1501),
        VN2CN2_bit => VN_data_out(1502),
        VN2CN3_bit => VN_data_out(1503),
        VN2CN4_bit => VN_data_out(1504),
        VN2CN5_bit => VN_data_out(1505),
        VN2CN0_sign => VN_sign_out(1500),
        VN2CN1_sign => VN_sign_out(1501),
        VN2CN2_sign => VN_sign_out(1502),
        VN2CN3_sign => VN_sign_out(1503),
        VN2CN4_sign => VN_sign_out(1504),
        VN2CN5_sign => VN_sign_out(1505),
        codeword => codeword(250),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN251 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1511 downto 1506),
        Din0 => VN251_in0,
        Din1 => VN251_in1,
        Din2 => VN251_in2,
        Din3 => VN251_in3,
        Din4 => VN251_in4,
        Din5 => VN251_in5,
        VN2CN0_bit => VN_data_out(1506),
        VN2CN1_bit => VN_data_out(1507),
        VN2CN2_bit => VN_data_out(1508),
        VN2CN3_bit => VN_data_out(1509),
        VN2CN4_bit => VN_data_out(1510),
        VN2CN5_bit => VN_data_out(1511),
        VN2CN0_sign => VN_sign_out(1506),
        VN2CN1_sign => VN_sign_out(1507),
        VN2CN2_sign => VN_sign_out(1508),
        VN2CN3_sign => VN_sign_out(1509),
        VN2CN4_sign => VN_sign_out(1510),
        VN2CN5_sign => VN_sign_out(1511),
        codeword => codeword(251),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN252 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1517 downto 1512),
        Din0 => VN252_in0,
        Din1 => VN252_in1,
        Din2 => VN252_in2,
        Din3 => VN252_in3,
        Din4 => VN252_in4,
        Din5 => VN252_in5,
        VN2CN0_bit => VN_data_out(1512),
        VN2CN1_bit => VN_data_out(1513),
        VN2CN2_bit => VN_data_out(1514),
        VN2CN3_bit => VN_data_out(1515),
        VN2CN4_bit => VN_data_out(1516),
        VN2CN5_bit => VN_data_out(1517),
        VN2CN0_sign => VN_sign_out(1512),
        VN2CN1_sign => VN_sign_out(1513),
        VN2CN2_sign => VN_sign_out(1514),
        VN2CN3_sign => VN_sign_out(1515),
        VN2CN4_sign => VN_sign_out(1516),
        VN2CN5_sign => VN_sign_out(1517),
        codeword => codeword(252),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN253 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1523 downto 1518),
        Din0 => VN253_in0,
        Din1 => VN253_in1,
        Din2 => VN253_in2,
        Din3 => VN253_in3,
        Din4 => VN253_in4,
        Din5 => VN253_in5,
        VN2CN0_bit => VN_data_out(1518),
        VN2CN1_bit => VN_data_out(1519),
        VN2CN2_bit => VN_data_out(1520),
        VN2CN3_bit => VN_data_out(1521),
        VN2CN4_bit => VN_data_out(1522),
        VN2CN5_bit => VN_data_out(1523),
        VN2CN0_sign => VN_sign_out(1518),
        VN2CN1_sign => VN_sign_out(1519),
        VN2CN2_sign => VN_sign_out(1520),
        VN2CN3_sign => VN_sign_out(1521),
        VN2CN4_sign => VN_sign_out(1522),
        VN2CN5_sign => VN_sign_out(1523),
        codeword => codeword(253),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN254 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1529 downto 1524),
        Din0 => VN254_in0,
        Din1 => VN254_in1,
        Din2 => VN254_in2,
        Din3 => VN254_in3,
        Din4 => VN254_in4,
        Din5 => VN254_in5,
        VN2CN0_bit => VN_data_out(1524),
        VN2CN1_bit => VN_data_out(1525),
        VN2CN2_bit => VN_data_out(1526),
        VN2CN3_bit => VN_data_out(1527),
        VN2CN4_bit => VN_data_out(1528),
        VN2CN5_bit => VN_data_out(1529),
        VN2CN0_sign => VN_sign_out(1524),
        VN2CN1_sign => VN_sign_out(1525),
        VN2CN2_sign => VN_sign_out(1526),
        VN2CN3_sign => VN_sign_out(1527),
        VN2CN4_sign => VN_sign_out(1528),
        VN2CN5_sign => VN_sign_out(1529),
        codeword => codeword(254),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN255 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1535 downto 1530),
        Din0 => VN255_in0,
        Din1 => VN255_in1,
        Din2 => VN255_in2,
        Din3 => VN255_in3,
        Din4 => VN255_in4,
        Din5 => VN255_in5,
        VN2CN0_bit => VN_data_out(1530),
        VN2CN1_bit => VN_data_out(1531),
        VN2CN2_bit => VN_data_out(1532),
        VN2CN3_bit => VN_data_out(1533),
        VN2CN4_bit => VN_data_out(1534),
        VN2CN5_bit => VN_data_out(1535),
        VN2CN0_sign => VN_sign_out(1530),
        VN2CN1_sign => VN_sign_out(1531),
        VN2CN2_sign => VN_sign_out(1532),
        VN2CN3_sign => VN_sign_out(1533),
        VN2CN4_sign => VN_sign_out(1534),
        VN2CN5_sign => VN_sign_out(1535),
        codeword => codeword(255),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN256 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1541 downto 1536),
        Din0 => VN256_in0,
        Din1 => VN256_in1,
        Din2 => VN256_in2,
        Din3 => VN256_in3,
        Din4 => VN256_in4,
        Din5 => VN256_in5,
        VN2CN0_bit => VN_data_out(1536),
        VN2CN1_bit => VN_data_out(1537),
        VN2CN2_bit => VN_data_out(1538),
        VN2CN3_bit => VN_data_out(1539),
        VN2CN4_bit => VN_data_out(1540),
        VN2CN5_bit => VN_data_out(1541),
        VN2CN0_sign => VN_sign_out(1536),
        VN2CN1_sign => VN_sign_out(1537),
        VN2CN2_sign => VN_sign_out(1538),
        VN2CN3_sign => VN_sign_out(1539),
        VN2CN4_sign => VN_sign_out(1540),
        VN2CN5_sign => VN_sign_out(1541),
        codeword => codeword(256),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN257 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1547 downto 1542),
        Din0 => VN257_in0,
        Din1 => VN257_in1,
        Din2 => VN257_in2,
        Din3 => VN257_in3,
        Din4 => VN257_in4,
        Din5 => VN257_in5,
        VN2CN0_bit => VN_data_out(1542),
        VN2CN1_bit => VN_data_out(1543),
        VN2CN2_bit => VN_data_out(1544),
        VN2CN3_bit => VN_data_out(1545),
        VN2CN4_bit => VN_data_out(1546),
        VN2CN5_bit => VN_data_out(1547),
        VN2CN0_sign => VN_sign_out(1542),
        VN2CN1_sign => VN_sign_out(1543),
        VN2CN2_sign => VN_sign_out(1544),
        VN2CN3_sign => VN_sign_out(1545),
        VN2CN4_sign => VN_sign_out(1546),
        VN2CN5_sign => VN_sign_out(1547),
        codeword => codeword(257),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN258 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1553 downto 1548),
        Din0 => VN258_in0,
        Din1 => VN258_in1,
        Din2 => VN258_in2,
        Din3 => VN258_in3,
        Din4 => VN258_in4,
        Din5 => VN258_in5,
        VN2CN0_bit => VN_data_out(1548),
        VN2CN1_bit => VN_data_out(1549),
        VN2CN2_bit => VN_data_out(1550),
        VN2CN3_bit => VN_data_out(1551),
        VN2CN4_bit => VN_data_out(1552),
        VN2CN5_bit => VN_data_out(1553),
        VN2CN0_sign => VN_sign_out(1548),
        VN2CN1_sign => VN_sign_out(1549),
        VN2CN2_sign => VN_sign_out(1550),
        VN2CN3_sign => VN_sign_out(1551),
        VN2CN4_sign => VN_sign_out(1552),
        VN2CN5_sign => VN_sign_out(1553),
        codeword => codeword(258),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN259 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1559 downto 1554),
        Din0 => VN259_in0,
        Din1 => VN259_in1,
        Din2 => VN259_in2,
        Din3 => VN259_in3,
        Din4 => VN259_in4,
        Din5 => VN259_in5,
        VN2CN0_bit => VN_data_out(1554),
        VN2CN1_bit => VN_data_out(1555),
        VN2CN2_bit => VN_data_out(1556),
        VN2CN3_bit => VN_data_out(1557),
        VN2CN4_bit => VN_data_out(1558),
        VN2CN5_bit => VN_data_out(1559),
        VN2CN0_sign => VN_sign_out(1554),
        VN2CN1_sign => VN_sign_out(1555),
        VN2CN2_sign => VN_sign_out(1556),
        VN2CN3_sign => VN_sign_out(1557),
        VN2CN4_sign => VN_sign_out(1558),
        VN2CN5_sign => VN_sign_out(1559),
        codeword => codeword(259),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN260 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1565 downto 1560),
        Din0 => VN260_in0,
        Din1 => VN260_in1,
        Din2 => VN260_in2,
        Din3 => VN260_in3,
        Din4 => VN260_in4,
        Din5 => VN260_in5,
        VN2CN0_bit => VN_data_out(1560),
        VN2CN1_bit => VN_data_out(1561),
        VN2CN2_bit => VN_data_out(1562),
        VN2CN3_bit => VN_data_out(1563),
        VN2CN4_bit => VN_data_out(1564),
        VN2CN5_bit => VN_data_out(1565),
        VN2CN0_sign => VN_sign_out(1560),
        VN2CN1_sign => VN_sign_out(1561),
        VN2CN2_sign => VN_sign_out(1562),
        VN2CN3_sign => VN_sign_out(1563),
        VN2CN4_sign => VN_sign_out(1564),
        VN2CN5_sign => VN_sign_out(1565),
        codeword => codeword(260),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN261 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1571 downto 1566),
        Din0 => VN261_in0,
        Din1 => VN261_in1,
        Din2 => VN261_in2,
        Din3 => VN261_in3,
        Din4 => VN261_in4,
        Din5 => VN261_in5,
        VN2CN0_bit => VN_data_out(1566),
        VN2CN1_bit => VN_data_out(1567),
        VN2CN2_bit => VN_data_out(1568),
        VN2CN3_bit => VN_data_out(1569),
        VN2CN4_bit => VN_data_out(1570),
        VN2CN5_bit => VN_data_out(1571),
        VN2CN0_sign => VN_sign_out(1566),
        VN2CN1_sign => VN_sign_out(1567),
        VN2CN2_sign => VN_sign_out(1568),
        VN2CN3_sign => VN_sign_out(1569),
        VN2CN4_sign => VN_sign_out(1570),
        VN2CN5_sign => VN_sign_out(1571),
        codeword => codeword(261),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN262 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1577 downto 1572),
        Din0 => VN262_in0,
        Din1 => VN262_in1,
        Din2 => VN262_in2,
        Din3 => VN262_in3,
        Din4 => VN262_in4,
        Din5 => VN262_in5,
        VN2CN0_bit => VN_data_out(1572),
        VN2CN1_bit => VN_data_out(1573),
        VN2CN2_bit => VN_data_out(1574),
        VN2CN3_bit => VN_data_out(1575),
        VN2CN4_bit => VN_data_out(1576),
        VN2CN5_bit => VN_data_out(1577),
        VN2CN0_sign => VN_sign_out(1572),
        VN2CN1_sign => VN_sign_out(1573),
        VN2CN2_sign => VN_sign_out(1574),
        VN2CN3_sign => VN_sign_out(1575),
        VN2CN4_sign => VN_sign_out(1576),
        VN2CN5_sign => VN_sign_out(1577),
        codeword => codeword(262),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN263 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1583 downto 1578),
        Din0 => VN263_in0,
        Din1 => VN263_in1,
        Din2 => VN263_in2,
        Din3 => VN263_in3,
        Din4 => VN263_in4,
        Din5 => VN263_in5,
        VN2CN0_bit => VN_data_out(1578),
        VN2CN1_bit => VN_data_out(1579),
        VN2CN2_bit => VN_data_out(1580),
        VN2CN3_bit => VN_data_out(1581),
        VN2CN4_bit => VN_data_out(1582),
        VN2CN5_bit => VN_data_out(1583),
        VN2CN0_sign => VN_sign_out(1578),
        VN2CN1_sign => VN_sign_out(1579),
        VN2CN2_sign => VN_sign_out(1580),
        VN2CN3_sign => VN_sign_out(1581),
        VN2CN4_sign => VN_sign_out(1582),
        VN2CN5_sign => VN_sign_out(1583),
        codeword => codeword(263),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN264 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1589 downto 1584),
        Din0 => VN264_in0,
        Din1 => VN264_in1,
        Din2 => VN264_in2,
        Din3 => VN264_in3,
        Din4 => VN264_in4,
        Din5 => VN264_in5,
        VN2CN0_bit => VN_data_out(1584),
        VN2CN1_bit => VN_data_out(1585),
        VN2CN2_bit => VN_data_out(1586),
        VN2CN3_bit => VN_data_out(1587),
        VN2CN4_bit => VN_data_out(1588),
        VN2CN5_bit => VN_data_out(1589),
        VN2CN0_sign => VN_sign_out(1584),
        VN2CN1_sign => VN_sign_out(1585),
        VN2CN2_sign => VN_sign_out(1586),
        VN2CN3_sign => VN_sign_out(1587),
        VN2CN4_sign => VN_sign_out(1588),
        VN2CN5_sign => VN_sign_out(1589),
        codeword => codeword(264),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN265 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1595 downto 1590),
        Din0 => VN265_in0,
        Din1 => VN265_in1,
        Din2 => VN265_in2,
        Din3 => VN265_in3,
        Din4 => VN265_in4,
        Din5 => VN265_in5,
        VN2CN0_bit => VN_data_out(1590),
        VN2CN1_bit => VN_data_out(1591),
        VN2CN2_bit => VN_data_out(1592),
        VN2CN3_bit => VN_data_out(1593),
        VN2CN4_bit => VN_data_out(1594),
        VN2CN5_bit => VN_data_out(1595),
        VN2CN0_sign => VN_sign_out(1590),
        VN2CN1_sign => VN_sign_out(1591),
        VN2CN2_sign => VN_sign_out(1592),
        VN2CN3_sign => VN_sign_out(1593),
        VN2CN4_sign => VN_sign_out(1594),
        VN2CN5_sign => VN_sign_out(1595),
        codeword => codeword(265),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN266 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1601 downto 1596),
        Din0 => VN266_in0,
        Din1 => VN266_in1,
        Din2 => VN266_in2,
        Din3 => VN266_in3,
        Din4 => VN266_in4,
        Din5 => VN266_in5,
        VN2CN0_bit => VN_data_out(1596),
        VN2CN1_bit => VN_data_out(1597),
        VN2CN2_bit => VN_data_out(1598),
        VN2CN3_bit => VN_data_out(1599),
        VN2CN4_bit => VN_data_out(1600),
        VN2CN5_bit => VN_data_out(1601),
        VN2CN0_sign => VN_sign_out(1596),
        VN2CN1_sign => VN_sign_out(1597),
        VN2CN2_sign => VN_sign_out(1598),
        VN2CN3_sign => VN_sign_out(1599),
        VN2CN4_sign => VN_sign_out(1600),
        VN2CN5_sign => VN_sign_out(1601),
        codeword => codeword(266),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN267 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1607 downto 1602),
        Din0 => VN267_in0,
        Din1 => VN267_in1,
        Din2 => VN267_in2,
        Din3 => VN267_in3,
        Din4 => VN267_in4,
        Din5 => VN267_in5,
        VN2CN0_bit => VN_data_out(1602),
        VN2CN1_bit => VN_data_out(1603),
        VN2CN2_bit => VN_data_out(1604),
        VN2CN3_bit => VN_data_out(1605),
        VN2CN4_bit => VN_data_out(1606),
        VN2CN5_bit => VN_data_out(1607),
        VN2CN0_sign => VN_sign_out(1602),
        VN2CN1_sign => VN_sign_out(1603),
        VN2CN2_sign => VN_sign_out(1604),
        VN2CN3_sign => VN_sign_out(1605),
        VN2CN4_sign => VN_sign_out(1606),
        VN2CN5_sign => VN_sign_out(1607),
        codeword => codeword(267),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN268 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1613 downto 1608),
        Din0 => VN268_in0,
        Din1 => VN268_in1,
        Din2 => VN268_in2,
        Din3 => VN268_in3,
        Din4 => VN268_in4,
        Din5 => VN268_in5,
        VN2CN0_bit => VN_data_out(1608),
        VN2CN1_bit => VN_data_out(1609),
        VN2CN2_bit => VN_data_out(1610),
        VN2CN3_bit => VN_data_out(1611),
        VN2CN4_bit => VN_data_out(1612),
        VN2CN5_bit => VN_data_out(1613),
        VN2CN0_sign => VN_sign_out(1608),
        VN2CN1_sign => VN_sign_out(1609),
        VN2CN2_sign => VN_sign_out(1610),
        VN2CN3_sign => VN_sign_out(1611),
        VN2CN4_sign => VN_sign_out(1612),
        VN2CN5_sign => VN_sign_out(1613),
        codeword => codeword(268),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN269 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1619 downto 1614),
        Din0 => VN269_in0,
        Din1 => VN269_in1,
        Din2 => VN269_in2,
        Din3 => VN269_in3,
        Din4 => VN269_in4,
        Din5 => VN269_in5,
        VN2CN0_bit => VN_data_out(1614),
        VN2CN1_bit => VN_data_out(1615),
        VN2CN2_bit => VN_data_out(1616),
        VN2CN3_bit => VN_data_out(1617),
        VN2CN4_bit => VN_data_out(1618),
        VN2CN5_bit => VN_data_out(1619),
        VN2CN0_sign => VN_sign_out(1614),
        VN2CN1_sign => VN_sign_out(1615),
        VN2CN2_sign => VN_sign_out(1616),
        VN2CN3_sign => VN_sign_out(1617),
        VN2CN4_sign => VN_sign_out(1618),
        VN2CN5_sign => VN_sign_out(1619),
        codeword => codeword(269),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN270 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1625 downto 1620),
        Din0 => VN270_in0,
        Din1 => VN270_in1,
        Din2 => VN270_in2,
        Din3 => VN270_in3,
        Din4 => VN270_in4,
        Din5 => VN270_in5,
        VN2CN0_bit => VN_data_out(1620),
        VN2CN1_bit => VN_data_out(1621),
        VN2CN2_bit => VN_data_out(1622),
        VN2CN3_bit => VN_data_out(1623),
        VN2CN4_bit => VN_data_out(1624),
        VN2CN5_bit => VN_data_out(1625),
        VN2CN0_sign => VN_sign_out(1620),
        VN2CN1_sign => VN_sign_out(1621),
        VN2CN2_sign => VN_sign_out(1622),
        VN2CN3_sign => VN_sign_out(1623),
        VN2CN4_sign => VN_sign_out(1624),
        VN2CN5_sign => VN_sign_out(1625),
        codeword => codeword(270),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN271 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1631 downto 1626),
        Din0 => VN271_in0,
        Din1 => VN271_in1,
        Din2 => VN271_in2,
        Din3 => VN271_in3,
        Din4 => VN271_in4,
        Din5 => VN271_in5,
        VN2CN0_bit => VN_data_out(1626),
        VN2CN1_bit => VN_data_out(1627),
        VN2CN2_bit => VN_data_out(1628),
        VN2CN3_bit => VN_data_out(1629),
        VN2CN4_bit => VN_data_out(1630),
        VN2CN5_bit => VN_data_out(1631),
        VN2CN0_sign => VN_sign_out(1626),
        VN2CN1_sign => VN_sign_out(1627),
        VN2CN2_sign => VN_sign_out(1628),
        VN2CN3_sign => VN_sign_out(1629),
        VN2CN4_sign => VN_sign_out(1630),
        VN2CN5_sign => VN_sign_out(1631),
        codeword => codeword(271),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN272 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1637 downto 1632),
        Din0 => VN272_in0,
        Din1 => VN272_in1,
        Din2 => VN272_in2,
        Din3 => VN272_in3,
        Din4 => VN272_in4,
        Din5 => VN272_in5,
        VN2CN0_bit => VN_data_out(1632),
        VN2CN1_bit => VN_data_out(1633),
        VN2CN2_bit => VN_data_out(1634),
        VN2CN3_bit => VN_data_out(1635),
        VN2CN4_bit => VN_data_out(1636),
        VN2CN5_bit => VN_data_out(1637),
        VN2CN0_sign => VN_sign_out(1632),
        VN2CN1_sign => VN_sign_out(1633),
        VN2CN2_sign => VN_sign_out(1634),
        VN2CN3_sign => VN_sign_out(1635),
        VN2CN4_sign => VN_sign_out(1636),
        VN2CN5_sign => VN_sign_out(1637),
        codeword => codeword(272),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN273 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1643 downto 1638),
        Din0 => VN273_in0,
        Din1 => VN273_in1,
        Din2 => VN273_in2,
        Din3 => VN273_in3,
        Din4 => VN273_in4,
        Din5 => VN273_in5,
        VN2CN0_bit => VN_data_out(1638),
        VN2CN1_bit => VN_data_out(1639),
        VN2CN2_bit => VN_data_out(1640),
        VN2CN3_bit => VN_data_out(1641),
        VN2CN4_bit => VN_data_out(1642),
        VN2CN5_bit => VN_data_out(1643),
        VN2CN0_sign => VN_sign_out(1638),
        VN2CN1_sign => VN_sign_out(1639),
        VN2CN2_sign => VN_sign_out(1640),
        VN2CN3_sign => VN_sign_out(1641),
        VN2CN4_sign => VN_sign_out(1642),
        VN2CN5_sign => VN_sign_out(1643),
        codeword => codeword(273),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN274 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1649 downto 1644),
        Din0 => VN274_in0,
        Din1 => VN274_in1,
        Din2 => VN274_in2,
        Din3 => VN274_in3,
        Din4 => VN274_in4,
        Din5 => VN274_in5,
        VN2CN0_bit => VN_data_out(1644),
        VN2CN1_bit => VN_data_out(1645),
        VN2CN2_bit => VN_data_out(1646),
        VN2CN3_bit => VN_data_out(1647),
        VN2CN4_bit => VN_data_out(1648),
        VN2CN5_bit => VN_data_out(1649),
        VN2CN0_sign => VN_sign_out(1644),
        VN2CN1_sign => VN_sign_out(1645),
        VN2CN2_sign => VN_sign_out(1646),
        VN2CN3_sign => VN_sign_out(1647),
        VN2CN4_sign => VN_sign_out(1648),
        VN2CN5_sign => VN_sign_out(1649),
        codeword => codeword(274),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN275 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1655 downto 1650),
        Din0 => VN275_in0,
        Din1 => VN275_in1,
        Din2 => VN275_in2,
        Din3 => VN275_in3,
        Din4 => VN275_in4,
        Din5 => VN275_in5,
        VN2CN0_bit => VN_data_out(1650),
        VN2CN1_bit => VN_data_out(1651),
        VN2CN2_bit => VN_data_out(1652),
        VN2CN3_bit => VN_data_out(1653),
        VN2CN4_bit => VN_data_out(1654),
        VN2CN5_bit => VN_data_out(1655),
        VN2CN0_sign => VN_sign_out(1650),
        VN2CN1_sign => VN_sign_out(1651),
        VN2CN2_sign => VN_sign_out(1652),
        VN2CN3_sign => VN_sign_out(1653),
        VN2CN4_sign => VN_sign_out(1654),
        VN2CN5_sign => VN_sign_out(1655),
        codeword => codeword(275),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN276 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1661 downto 1656),
        Din0 => VN276_in0,
        Din1 => VN276_in1,
        Din2 => VN276_in2,
        Din3 => VN276_in3,
        Din4 => VN276_in4,
        Din5 => VN276_in5,
        VN2CN0_bit => VN_data_out(1656),
        VN2CN1_bit => VN_data_out(1657),
        VN2CN2_bit => VN_data_out(1658),
        VN2CN3_bit => VN_data_out(1659),
        VN2CN4_bit => VN_data_out(1660),
        VN2CN5_bit => VN_data_out(1661),
        VN2CN0_sign => VN_sign_out(1656),
        VN2CN1_sign => VN_sign_out(1657),
        VN2CN2_sign => VN_sign_out(1658),
        VN2CN3_sign => VN_sign_out(1659),
        VN2CN4_sign => VN_sign_out(1660),
        VN2CN5_sign => VN_sign_out(1661),
        codeword => codeword(276),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN277 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1667 downto 1662),
        Din0 => VN277_in0,
        Din1 => VN277_in1,
        Din2 => VN277_in2,
        Din3 => VN277_in3,
        Din4 => VN277_in4,
        Din5 => VN277_in5,
        VN2CN0_bit => VN_data_out(1662),
        VN2CN1_bit => VN_data_out(1663),
        VN2CN2_bit => VN_data_out(1664),
        VN2CN3_bit => VN_data_out(1665),
        VN2CN4_bit => VN_data_out(1666),
        VN2CN5_bit => VN_data_out(1667),
        VN2CN0_sign => VN_sign_out(1662),
        VN2CN1_sign => VN_sign_out(1663),
        VN2CN2_sign => VN_sign_out(1664),
        VN2CN3_sign => VN_sign_out(1665),
        VN2CN4_sign => VN_sign_out(1666),
        VN2CN5_sign => VN_sign_out(1667),
        codeword => codeword(277),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN278 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1673 downto 1668),
        Din0 => VN278_in0,
        Din1 => VN278_in1,
        Din2 => VN278_in2,
        Din3 => VN278_in3,
        Din4 => VN278_in4,
        Din5 => VN278_in5,
        VN2CN0_bit => VN_data_out(1668),
        VN2CN1_bit => VN_data_out(1669),
        VN2CN2_bit => VN_data_out(1670),
        VN2CN3_bit => VN_data_out(1671),
        VN2CN4_bit => VN_data_out(1672),
        VN2CN5_bit => VN_data_out(1673),
        VN2CN0_sign => VN_sign_out(1668),
        VN2CN1_sign => VN_sign_out(1669),
        VN2CN2_sign => VN_sign_out(1670),
        VN2CN3_sign => VN_sign_out(1671),
        VN2CN4_sign => VN_sign_out(1672),
        VN2CN5_sign => VN_sign_out(1673),
        codeword => codeword(278),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN279 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1679 downto 1674),
        Din0 => VN279_in0,
        Din1 => VN279_in1,
        Din2 => VN279_in2,
        Din3 => VN279_in3,
        Din4 => VN279_in4,
        Din5 => VN279_in5,
        VN2CN0_bit => VN_data_out(1674),
        VN2CN1_bit => VN_data_out(1675),
        VN2CN2_bit => VN_data_out(1676),
        VN2CN3_bit => VN_data_out(1677),
        VN2CN4_bit => VN_data_out(1678),
        VN2CN5_bit => VN_data_out(1679),
        VN2CN0_sign => VN_sign_out(1674),
        VN2CN1_sign => VN_sign_out(1675),
        VN2CN2_sign => VN_sign_out(1676),
        VN2CN3_sign => VN_sign_out(1677),
        VN2CN4_sign => VN_sign_out(1678),
        VN2CN5_sign => VN_sign_out(1679),
        codeword => codeword(279),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN280 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1685 downto 1680),
        Din0 => VN280_in0,
        Din1 => VN280_in1,
        Din2 => VN280_in2,
        Din3 => VN280_in3,
        Din4 => VN280_in4,
        Din5 => VN280_in5,
        VN2CN0_bit => VN_data_out(1680),
        VN2CN1_bit => VN_data_out(1681),
        VN2CN2_bit => VN_data_out(1682),
        VN2CN3_bit => VN_data_out(1683),
        VN2CN4_bit => VN_data_out(1684),
        VN2CN5_bit => VN_data_out(1685),
        VN2CN0_sign => VN_sign_out(1680),
        VN2CN1_sign => VN_sign_out(1681),
        VN2CN2_sign => VN_sign_out(1682),
        VN2CN3_sign => VN_sign_out(1683),
        VN2CN4_sign => VN_sign_out(1684),
        VN2CN5_sign => VN_sign_out(1685),
        codeword => codeword(280),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN281 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1691 downto 1686),
        Din0 => VN281_in0,
        Din1 => VN281_in1,
        Din2 => VN281_in2,
        Din3 => VN281_in3,
        Din4 => VN281_in4,
        Din5 => VN281_in5,
        VN2CN0_bit => VN_data_out(1686),
        VN2CN1_bit => VN_data_out(1687),
        VN2CN2_bit => VN_data_out(1688),
        VN2CN3_bit => VN_data_out(1689),
        VN2CN4_bit => VN_data_out(1690),
        VN2CN5_bit => VN_data_out(1691),
        VN2CN0_sign => VN_sign_out(1686),
        VN2CN1_sign => VN_sign_out(1687),
        VN2CN2_sign => VN_sign_out(1688),
        VN2CN3_sign => VN_sign_out(1689),
        VN2CN4_sign => VN_sign_out(1690),
        VN2CN5_sign => VN_sign_out(1691),
        codeword => codeword(281),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN282 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1697 downto 1692),
        Din0 => VN282_in0,
        Din1 => VN282_in1,
        Din2 => VN282_in2,
        Din3 => VN282_in3,
        Din4 => VN282_in4,
        Din5 => VN282_in5,
        VN2CN0_bit => VN_data_out(1692),
        VN2CN1_bit => VN_data_out(1693),
        VN2CN2_bit => VN_data_out(1694),
        VN2CN3_bit => VN_data_out(1695),
        VN2CN4_bit => VN_data_out(1696),
        VN2CN5_bit => VN_data_out(1697),
        VN2CN0_sign => VN_sign_out(1692),
        VN2CN1_sign => VN_sign_out(1693),
        VN2CN2_sign => VN_sign_out(1694),
        VN2CN3_sign => VN_sign_out(1695),
        VN2CN4_sign => VN_sign_out(1696),
        VN2CN5_sign => VN_sign_out(1697),
        codeword => codeword(282),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN283 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1703 downto 1698),
        Din0 => VN283_in0,
        Din1 => VN283_in1,
        Din2 => VN283_in2,
        Din3 => VN283_in3,
        Din4 => VN283_in4,
        Din5 => VN283_in5,
        VN2CN0_bit => VN_data_out(1698),
        VN2CN1_bit => VN_data_out(1699),
        VN2CN2_bit => VN_data_out(1700),
        VN2CN3_bit => VN_data_out(1701),
        VN2CN4_bit => VN_data_out(1702),
        VN2CN5_bit => VN_data_out(1703),
        VN2CN0_sign => VN_sign_out(1698),
        VN2CN1_sign => VN_sign_out(1699),
        VN2CN2_sign => VN_sign_out(1700),
        VN2CN3_sign => VN_sign_out(1701),
        VN2CN4_sign => VN_sign_out(1702),
        VN2CN5_sign => VN_sign_out(1703),
        codeword => codeword(283),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN284 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1709 downto 1704),
        Din0 => VN284_in0,
        Din1 => VN284_in1,
        Din2 => VN284_in2,
        Din3 => VN284_in3,
        Din4 => VN284_in4,
        Din5 => VN284_in5,
        VN2CN0_bit => VN_data_out(1704),
        VN2CN1_bit => VN_data_out(1705),
        VN2CN2_bit => VN_data_out(1706),
        VN2CN3_bit => VN_data_out(1707),
        VN2CN4_bit => VN_data_out(1708),
        VN2CN5_bit => VN_data_out(1709),
        VN2CN0_sign => VN_sign_out(1704),
        VN2CN1_sign => VN_sign_out(1705),
        VN2CN2_sign => VN_sign_out(1706),
        VN2CN3_sign => VN_sign_out(1707),
        VN2CN4_sign => VN_sign_out(1708),
        VN2CN5_sign => VN_sign_out(1709),
        codeword => codeword(284),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN285 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1715 downto 1710),
        Din0 => VN285_in0,
        Din1 => VN285_in1,
        Din2 => VN285_in2,
        Din3 => VN285_in3,
        Din4 => VN285_in4,
        Din5 => VN285_in5,
        VN2CN0_bit => VN_data_out(1710),
        VN2CN1_bit => VN_data_out(1711),
        VN2CN2_bit => VN_data_out(1712),
        VN2CN3_bit => VN_data_out(1713),
        VN2CN4_bit => VN_data_out(1714),
        VN2CN5_bit => VN_data_out(1715),
        VN2CN0_sign => VN_sign_out(1710),
        VN2CN1_sign => VN_sign_out(1711),
        VN2CN2_sign => VN_sign_out(1712),
        VN2CN3_sign => VN_sign_out(1713),
        VN2CN4_sign => VN_sign_out(1714),
        VN2CN5_sign => VN_sign_out(1715),
        codeword => codeword(285),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN286 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1721 downto 1716),
        Din0 => VN286_in0,
        Din1 => VN286_in1,
        Din2 => VN286_in2,
        Din3 => VN286_in3,
        Din4 => VN286_in4,
        Din5 => VN286_in5,
        VN2CN0_bit => VN_data_out(1716),
        VN2CN1_bit => VN_data_out(1717),
        VN2CN2_bit => VN_data_out(1718),
        VN2CN3_bit => VN_data_out(1719),
        VN2CN4_bit => VN_data_out(1720),
        VN2CN5_bit => VN_data_out(1721),
        VN2CN0_sign => VN_sign_out(1716),
        VN2CN1_sign => VN_sign_out(1717),
        VN2CN2_sign => VN_sign_out(1718),
        VN2CN3_sign => VN_sign_out(1719),
        VN2CN4_sign => VN_sign_out(1720),
        VN2CN5_sign => VN_sign_out(1721),
        codeword => codeword(286),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN287 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1727 downto 1722),
        Din0 => VN287_in0,
        Din1 => VN287_in1,
        Din2 => VN287_in2,
        Din3 => VN287_in3,
        Din4 => VN287_in4,
        Din5 => VN287_in5,
        VN2CN0_bit => VN_data_out(1722),
        VN2CN1_bit => VN_data_out(1723),
        VN2CN2_bit => VN_data_out(1724),
        VN2CN3_bit => VN_data_out(1725),
        VN2CN4_bit => VN_data_out(1726),
        VN2CN5_bit => VN_data_out(1727),
        VN2CN0_sign => VN_sign_out(1722),
        VN2CN1_sign => VN_sign_out(1723),
        VN2CN2_sign => VN_sign_out(1724),
        VN2CN3_sign => VN_sign_out(1725),
        VN2CN4_sign => VN_sign_out(1726),
        VN2CN5_sign => VN_sign_out(1727),
        codeword => codeword(287),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN288 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1733 downto 1728),
        Din0 => VN288_in0,
        Din1 => VN288_in1,
        Din2 => VN288_in2,
        Din3 => VN288_in3,
        Din4 => VN288_in4,
        Din5 => VN288_in5,
        VN2CN0_bit => VN_data_out(1728),
        VN2CN1_bit => VN_data_out(1729),
        VN2CN2_bit => VN_data_out(1730),
        VN2CN3_bit => VN_data_out(1731),
        VN2CN4_bit => VN_data_out(1732),
        VN2CN5_bit => VN_data_out(1733),
        VN2CN0_sign => VN_sign_out(1728),
        VN2CN1_sign => VN_sign_out(1729),
        VN2CN2_sign => VN_sign_out(1730),
        VN2CN3_sign => VN_sign_out(1731),
        VN2CN4_sign => VN_sign_out(1732),
        VN2CN5_sign => VN_sign_out(1733),
        codeword => codeword(288),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN289 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1739 downto 1734),
        Din0 => VN289_in0,
        Din1 => VN289_in1,
        Din2 => VN289_in2,
        Din3 => VN289_in3,
        Din4 => VN289_in4,
        Din5 => VN289_in5,
        VN2CN0_bit => VN_data_out(1734),
        VN2CN1_bit => VN_data_out(1735),
        VN2CN2_bit => VN_data_out(1736),
        VN2CN3_bit => VN_data_out(1737),
        VN2CN4_bit => VN_data_out(1738),
        VN2CN5_bit => VN_data_out(1739),
        VN2CN0_sign => VN_sign_out(1734),
        VN2CN1_sign => VN_sign_out(1735),
        VN2CN2_sign => VN_sign_out(1736),
        VN2CN3_sign => VN_sign_out(1737),
        VN2CN4_sign => VN_sign_out(1738),
        VN2CN5_sign => VN_sign_out(1739),
        codeword => codeword(289),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN290 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1745 downto 1740),
        Din0 => VN290_in0,
        Din1 => VN290_in1,
        Din2 => VN290_in2,
        Din3 => VN290_in3,
        Din4 => VN290_in4,
        Din5 => VN290_in5,
        VN2CN0_bit => VN_data_out(1740),
        VN2CN1_bit => VN_data_out(1741),
        VN2CN2_bit => VN_data_out(1742),
        VN2CN3_bit => VN_data_out(1743),
        VN2CN4_bit => VN_data_out(1744),
        VN2CN5_bit => VN_data_out(1745),
        VN2CN0_sign => VN_sign_out(1740),
        VN2CN1_sign => VN_sign_out(1741),
        VN2CN2_sign => VN_sign_out(1742),
        VN2CN3_sign => VN_sign_out(1743),
        VN2CN4_sign => VN_sign_out(1744),
        VN2CN5_sign => VN_sign_out(1745),
        codeword => codeword(290),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN291 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1751 downto 1746),
        Din0 => VN291_in0,
        Din1 => VN291_in1,
        Din2 => VN291_in2,
        Din3 => VN291_in3,
        Din4 => VN291_in4,
        Din5 => VN291_in5,
        VN2CN0_bit => VN_data_out(1746),
        VN2CN1_bit => VN_data_out(1747),
        VN2CN2_bit => VN_data_out(1748),
        VN2CN3_bit => VN_data_out(1749),
        VN2CN4_bit => VN_data_out(1750),
        VN2CN5_bit => VN_data_out(1751),
        VN2CN0_sign => VN_sign_out(1746),
        VN2CN1_sign => VN_sign_out(1747),
        VN2CN2_sign => VN_sign_out(1748),
        VN2CN3_sign => VN_sign_out(1749),
        VN2CN4_sign => VN_sign_out(1750),
        VN2CN5_sign => VN_sign_out(1751),
        codeword => codeword(291),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN292 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1757 downto 1752),
        Din0 => VN292_in0,
        Din1 => VN292_in1,
        Din2 => VN292_in2,
        Din3 => VN292_in3,
        Din4 => VN292_in4,
        Din5 => VN292_in5,
        VN2CN0_bit => VN_data_out(1752),
        VN2CN1_bit => VN_data_out(1753),
        VN2CN2_bit => VN_data_out(1754),
        VN2CN3_bit => VN_data_out(1755),
        VN2CN4_bit => VN_data_out(1756),
        VN2CN5_bit => VN_data_out(1757),
        VN2CN0_sign => VN_sign_out(1752),
        VN2CN1_sign => VN_sign_out(1753),
        VN2CN2_sign => VN_sign_out(1754),
        VN2CN3_sign => VN_sign_out(1755),
        VN2CN4_sign => VN_sign_out(1756),
        VN2CN5_sign => VN_sign_out(1757),
        codeword => codeword(292),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN293 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1763 downto 1758),
        Din0 => VN293_in0,
        Din1 => VN293_in1,
        Din2 => VN293_in2,
        Din3 => VN293_in3,
        Din4 => VN293_in4,
        Din5 => VN293_in5,
        VN2CN0_bit => VN_data_out(1758),
        VN2CN1_bit => VN_data_out(1759),
        VN2CN2_bit => VN_data_out(1760),
        VN2CN3_bit => VN_data_out(1761),
        VN2CN4_bit => VN_data_out(1762),
        VN2CN5_bit => VN_data_out(1763),
        VN2CN0_sign => VN_sign_out(1758),
        VN2CN1_sign => VN_sign_out(1759),
        VN2CN2_sign => VN_sign_out(1760),
        VN2CN3_sign => VN_sign_out(1761),
        VN2CN4_sign => VN_sign_out(1762),
        VN2CN5_sign => VN_sign_out(1763),
        codeword => codeword(293),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN294 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1769 downto 1764),
        Din0 => VN294_in0,
        Din1 => VN294_in1,
        Din2 => VN294_in2,
        Din3 => VN294_in3,
        Din4 => VN294_in4,
        Din5 => VN294_in5,
        VN2CN0_bit => VN_data_out(1764),
        VN2CN1_bit => VN_data_out(1765),
        VN2CN2_bit => VN_data_out(1766),
        VN2CN3_bit => VN_data_out(1767),
        VN2CN4_bit => VN_data_out(1768),
        VN2CN5_bit => VN_data_out(1769),
        VN2CN0_sign => VN_sign_out(1764),
        VN2CN1_sign => VN_sign_out(1765),
        VN2CN2_sign => VN_sign_out(1766),
        VN2CN3_sign => VN_sign_out(1767),
        VN2CN4_sign => VN_sign_out(1768),
        VN2CN5_sign => VN_sign_out(1769),
        codeword => codeword(294),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN295 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1775 downto 1770),
        Din0 => VN295_in0,
        Din1 => VN295_in1,
        Din2 => VN295_in2,
        Din3 => VN295_in3,
        Din4 => VN295_in4,
        Din5 => VN295_in5,
        VN2CN0_bit => VN_data_out(1770),
        VN2CN1_bit => VN_data_out(1771),
        VN2CN2_bit => VN_data_out(1772),
        VN2CN3_bit => VN_data_out(1773),
        VN2CN4_bit => VN_data_out(1774),
        VN2CN5_bit => VN_data_out(1775),
        VN2CN0_sign => VN_sign_out(1770),
        VN2CN1_sign => VN_sign_out(1771),
        VN2CN2_sign => VN_sign_out(1772),
        VN2CN3_sign => VN_sign_out(1773),
        VN2CN4_sign => VN_sign_out(1774),
        VN2CN5_sign => VN_sign_out(1775),
        codeword => codeword(295),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN296 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1781 downto 1776),
        Din0 => VN296_in0,
        Din1 => VN296_in1,
        Din2 => VN296_in2,
        Din3 => VN296_in3,
        Din4 => VN296_in4,
        Din5 => VN296_in5,
        VN2CN0_bit => VN_data_out(1776),
        VN2CN1_bit => VN_data_out(1777),
        VN2CN2_bit => VN_data_out(1778),
        VN2CN3_bit => VN_data_out(1779),
        VN2CN4_bit => VN_data_out(1780),
        VN2CN5_bit => VN_data_out(1781),
        VN2CN0_sign => VN_sign_out(1776),
        VN2CN1_sign => VN_sign_out(1777),
        VN2CN2_sign => VN_sign_out(1778),
        VN2CN3_sign => VN_sign_out(1779),
        VN2CN4_sign => VN_sign_out(1780),
        VN2CN5_sign => VN_sign_out(1781),
        codeword => codeword(296),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN297 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1787 downto 1782),
        Din0 => VN297_in0,
        Din1 => VN297_in1,
        Din2 => VN297_in2,
        Din3 => VN297_in3,
        Din4 => VN297_in4,
        Din5 => VN297_in5,
        VN2CN0_bit => VN_data_out(1782),
        VN2CN1_bit => VN_data_out(1783),
        VN2CN2_bit => VN_data_out(1784),
        VN2CN3_bit => VN_data_out(1785),
        VN2CN4_bit => VN_data_out(1786),
        VN2CN5_bit => VN_data_out(1787),
        VN2CN0_sign => VN_sign_out(1782),
        VN2CN1_sign => VN_sign_out(1783),
        VN2CN2_sign => VN_sign_out(1784),
        VN2CN3_sign => VN_sign_out(1785),
        VN2CN4_sign => VN_sign_out(1786),
        VN2CN5_sign => VN_sign_out(1787),
        codeword => codeword(297),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN298 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1793 downto 1788),
        Din0 => VN298_in0,
        Din1 => VN298_in1,
        Din2 => VN298_in2,
        Din3 => VN298_in3,
        Din4 => VN298_in4,
        Din5 => VN298_in5,
        VN2CN0_bit => VN_data_out(1788),
        VN2CN1_bit => VN_data_out(1789),
        VN2CN2_bit => VN_data_out(1790),
        VN2CN3_bit => VN_data_out(1791),
        VN2CN4_bit => VN_data_out(1792),
        VN2CN5_bit => VN_data_out(1793),
        VN2CN0_sign => VN_sign_out(1788),
        VN2CN1_sign => VN_sign_out(1789),
        VN2CN2_sign => VN_sign_out(1790),
        VN2CN3_sign => VN_sign_out(1791),
        VN2CN4_sign => VN_sign_out(1792),
        VN2CN5_sign => VN_sign_out(1793),
        codeword => codeword(298),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN299 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1799 downto 1794),
        Din0 => VN299_in0,
        Din1 => VN299_in1,
        Din2 => VN299_in2,
        Din3 => VN299_in3,
        Din4 => VN299_in4,
        Din5 => VN299_in5,
        VN2CN0_bit => VN_data_out(1794),
        VN2CN1_bit => VN_data_out(1795),
        VN2CN2_bit => VN_data_out(1796),
        VN2CN3_bit => VN_data_out(1797),
        VN2CN4_bit => VN_data_out(1798),
        VN2CN5_bit => VN_data_out(1799),
        VN2CN0_sign => VN_sign_out(1794),
        VN2CN1_sign => VN_sign_out(1795),
        VN2CN2_sign => VN_sign_out(1796),
        VN2CN3_sign => VN_sign_out(1797),
        VN2CN4_sign => VN_sign_out(1798),
        VN2CN5_sign => VN_sign_out(1799),
        codeword => codeword(299),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN300 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1805 downto 1800),
        Din0 => VN300_in0,
        Din1 => VN300_in1,
        Din2 => VN300_in2,
        Din3 => VN300_in3,
        Din4 => VN300_in4,
        Din5 => VN300_in5,
        VN2CN0_bit => VN_data_out(1800),
        VN2CN1_bit => VN_data_out(1801),
        VN2CN2_bit => VN_data_out(1802),
        VN2CN3_bit => VN_data_out(1803),
        VN2CN4_bit => VN_data_out(1804),
        VN2CN5_bit => VN_data_out(1805),
        VN2CN0_sign => VN_sign_out(1800),
        VN2CN1_sign => VN_sign_out(1801),
        VN2CN2_sign => VN_sign_out(1802),
        VN2CN3_sign => VN_sign_out(1803),
        VN2CN4_sign => VN_sign_out(1804),
        VN2CN5_sign => VN_sign_out(1805),
        codeword => codeword(300),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN301 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1811 downto 1806),
        Din0 => VN301_in0,
        Din1 => VN301_in1,
        Din2 => VN301_in2,
        Din3 => VN301_in3,
        Din4 => VN301_in4,
        Din5 => VN301_in5,
        VN2CN0_bit => VN_data_out(1806),
        VN2CN1_bit => VN_data_out(1807),
        VN2CN2_bit => VN_data_out(1808),
        VN2CN3_bit => VN_data_out(1809),
        VN2CN4_bit => VN_data_out(1810),
        VN2CN5_bit => VN_data_out(1811),
        VN2CN0_sign => VN_sign_out(1806),
        VN2CN1_sign => VN_sign_out(1807),
        VN2CN2_sign => VN_sign_out(1808),
        VN2CN3_sign => VN_sign_out(1809),
        VN2CN4_sign => VN_sign_out(1810),
        VN2CN5_sign => VN_sign_out(1811),
        codeword => codeword(301),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN302 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1817 downto 1812),
        Din0 => VN302_in0,
        Din1 => VN302_in1,
        Din2 => VN302_in2,
        Din3 => VN302_in3,
        Din4 => VN302_in4,
        Din5 => VN302_in5,
        VN2CN0_bit => VN_data_out(1812),
        VN2CN1_bit => VN_data_out(1813),
        VN2CN2_bit => VN_data_out(1814),
        VN2CN3_bit => VN_data_out(1815),
        VN2CN4_bit => VN_data_out(1816),
        VN2CN5_bit => VN_data_out(1817),
        VN2CN0_sign => VN_sign_out(1812),
        VN2CN1_sign => VN_sign_out(1813),
        VN2CN2_sign => VN_sign_out(1814),
        VN2CN3_sign => VN_sign_out(1815),
        VN2CN4_sign => VN_sign_out(1816),
        VN2CN5_sign => VN_sign_out(1817),
        codeword => codeword(302),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN303 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1823 downto 1818),
        Din0 => VN303_in0,
        Din1 => VN303_in1,
        Din2 => VN303_in2,
        Din3 => VN303_in3,
        Din4 => VN303_in4,
        Din5 => VN303_in5,
        VN2CN0_bit => VN_data_out(1818),
        VN2CN1_bit => VN_data_out(1819),
        VN2CN2_bit => VN_data_out(1820),
        VN2CN3_bit => VN_data_out(1821),
        VN2CN4_bit => VN_data_out(1822),
        VN2CN5_bit => VN_data_out(1823),
        VN2CN0_sign => VN_sign_out(1818),
        VN2CN1_sign => VN_sign_out(1819),
        VN2CN2_sign => VN_sign_out(1820),
        VN2CN3_sign => VN_sign_out(1821),
        VN2CN4_sign => VN_sign_out(1822),
        VN2CN5_sign => VN_sign_out(1823),
        codeword => codeword(303),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN304 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1829 downto 1824),
        Din0 => VN304_in0,
        Din1 => VN304_in1,
        Din2 => VN304_in2,
        Din3 => VN304_in3,
        Din4 => VN304_in4,
        Din5 => VN304_in5,
        VN2CN0_bit => VN_data_out(1824),
        VN2CN1_bit => VN_data_out(1825),
        VN2CN2_bit => VN_data_out(1826),
        VN2CN3_bit => VN_data_out(1827),
        VN2CN4_bit => VN_data_out(1828),
        VN2CN5_bit => VN_data_out(1829),
        VN2CN0_sign => VN_sign_out(1824),
        VN2CN1_sign => VN_sign_out(1825),
        VN2CN2_sign => VN_sign_out(1826),
        VN2CN3_sign => VN_sign_out(1827),
        VN2CN4_sign => VN_sign_out(1828),
        VN2CN5_sign => VN_sign_out(1829),
        codeword => codeword(304),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN305 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1835 downto 1830),
        Din0 => VN305_in0,
        Din1 => VN305_in1,
        Din2 => VN305_in2,
        Din3 => VN305_in3,
        Din4 => VN305_in4,
        Din5 => VN305_in5,
        VN2CN0_bit => VN_data_out(1830),
        VN2CN1_bit => VN_data_out(1831),
        VN2CN2_bit => VN_data_out(1832),
        VN2CN3_bit => VN_data_out(1833),
        VN2CN4_bit => VN_data_out(1834),
        VN2CN5_bit => VN_data_out(1835),
        VN2CN0_sign => VN_sign_out(1830),
        VN2CN1_sign => VN_sign_out(1831),
        VN2CN2_sign => VN_sign_out(1832),
        VN2CN3_sign => VN_sign_out(1833),
        VN2CN4_sign => VN_sign_out(1834),
        VN2CN5_sign => VN_sign_out(1835),
        codeword => codeword(305),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN306 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1841 downto 1836),
        Din0 => VN306_in0,
        Din1 => VN306_in1,
        Din2 => VN306_in2,
        Din3 => VN306_in3,
        Din4 => VN306_in4,
        Din5 => VN306_in5,
        VN2CN0_bit => VN_data_out(1836),
        VN2CN1_bit => VN_data_out(1837),
        VN2CN2_bit => VN_data_out(1838),
        VN2CN3_bit => VN_data_out(1839),
        VN2CN4_bit => VN_data_out(1840),
        VN2CN5_bit => VN_data_out(1841),
        VN2CN0_sign => VN_sign_out(1836),
        VN2CN1_sign => VN_sign_out(1837),
        VN2CN2_sign => VN_sign_out(1838),
        VN2CN3_sign => VN_sign_out(1839),
        VN2CN4_sign => VN_sign_out(1840),
        VN2CN5_sign => VN_sign_out(1841),
        codeword => codeword(306),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN307 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1847 downto 1842),
        Din0 => VN307_in0,
        Din1 => VN307_in1,
        Din2 => VN307_in2,
        Din3 => VN307_in3,
        Din4 => VN307_in4,
        Din5 => VN307_in5,
        VN2CN0_bit => VN_data_out(1842),
        VN2CN1_bit => VN_data_out(1843),
        VN2CN2_bit => VN_data_out(1844),
        VN2CN3_bit => VN_data_out(1845),
        VN2CN4_bit => VN_data_out(1846),
        VN2CN5_bit => VN_data_out(1847),
        VN2CN0_sign => VN_sign_out(1842),
        VN2CN1_sign => VN_sign_out(1843),
        VN2CN2_sign => VN_sign_out(1844),
        VN2CN3_sign => VN_sign_out(1845),
        VN2CN4_sign => VN_sign_out(1846),
        VN2CN5_sign => VN_sign_out(1847),
        codeword => codeword(307),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN308 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1853 downto 1848),
        Din0 => VN308_in0,
        Din1 => VN308_in1,
        Din2 => VN308_in2,
        Din3 => VN308_in3,
        Din4 => VN308_in4,
        Din5 => VN308_in5,
        VN2CN0_bit => VN_data_out(1848),
        VN2CN1_bit => VN_data_out(1849),
        VN2CN2_bit => VN_data_out(1850),
        VN2CN3_bit => VN_data_out(1851),
        VN2CN4_bit => VN_data_out(1852),
        VN2CN5_bit => VN_data_out(1853),
        VN2CN0_sign => VN_sign_out(1848),
        VN2CN1_sign => VN_sign_out(1849),
        VN2CN2_sign => VN_sign_out(1850),
        VN2CN3_sign => VN_sign_out(1851),
        VN2CN4_sign => VN_sign_out(1852),
        VN2CN5_sign => VN_sign_out(1853),
        codeword => codeword(308),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN309 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1859 downto 1854),
        Din0 => VN309_in0,
        Din1 => VN309_in1,
        Din2 => VN309_in2,
        Din3 => VN309_in3,
        Din4 => VN309_in4,
        Din5 => VN309_in5,
        VN2CN0_bit => VN_data_out(1854),
        VN2CN1_bit => VN_data_out(1855),
        VN2CN2_bit => VN_data_out(1856),
        VN2CN3_bit => VN_data_out(1857),
        VN2CN4_bit => VN_data_out(1858),
        VN2CN5_bit => VN_data_out(1859),
        VN2CN0_sign => VN_sign_out(1854),
        VN2CN1_sign => VN_sign_out(1855),
        VN2CN2_sign => VN_sign_out(1856),
        VN2CN3_sign => VN_sign_out(1857),
        VN2CN4_sign => VN_sign_out(1858),
        VN2CN5_sign => VN_sign_out(1859),
        codeword => codeword(309),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN310 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1865 downto 1860),
        Din0 => VN310_in0,
        Din1 => VN310_in1,
        Din2 => VN310_in2,
        Din3 => VN310_in3,
        Din4 => VN310_in4,
        Din5 => VN310_in5,
        VN2CN0_bit => VN_data_out(1860),
        VN2CN1_bit => VN_data_out(1861),
        VN2CN2_bit => VN_data_out(1862),
        VN2CN3_bit => VN_data_out(1863),
        VN2CN4_bit => VN_data_out(1864),
        VN2CN5_bit => VN_data_out(1865),
        VN2CN0_sign => VN_sign_out(1860),
        VN2CN1_sign => VN_sign_out(1861),
        VN2CN2_sign => VN_sign_out(1862),
        VN2CN3_sign => VN_sign_out(1863),
        VN2CN4_sign => VN_sign_out(1864),
        VN2CN5_sign => VN_sign_out(1865),
        codeword => codeword(310),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN311 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1871 downto 1866),
        Din0 => VN311_in0,
        Din1 => VN311_in1,
        Din2 => VN311_in2,
        Din3 => VN311_in3,
        Din4 => VN311_in4,
        Din5 => VN311_in5,
        VN2CN0_bit => VN_data_out(1866),
        VN2CN1_bit => VN_data_out(1867),
        VN2CN2_bit => VN_data_out(1868),
        VN2CN3_bit => VN_data_out(1869),
        VN2CN4_bit => VN_data_out(1870),
        VN2CN5_bit => VN_data_out(1871),
        VN2CN0_sign => VN_sign_out(1866),
        VN2CN1_sign => VN_sign_out(1867),
        VN2CN2_sign => VN_sign_out(1868),
        VN2CN3_sign => VN_sign_out(1869),
        VN2CN4_sign => VN_sign_out(1870),
        VN2CN5_sign => VN_sign_out(1871),
        codeword => codeword(311),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN312 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1877 downto 1872),
        Din0 => VN312_in0,
        Din1 => VN312_in1,
        Din2 => VN312_in2,
        Din3 => VN312_in3,
        Din4 => VN312_in4,
        Din5 => VN312_in5,
        VN2CN0_bit => VN_data_out(1872),
        VN2CN1_bit => VN_data_out(1873),
        VN2CN2_bit => VN_data_out(1874),
        VN2CN3_bit => VN_data_out(1875),
        VN2CN4_bit => VN_data_out(1876),
        VN2CN5_bit => VN_data_out(1877),
        VN2CN0_sign => VN_sign_out(1872),
        VN2CN1_sign => VN_sign_out(1873),
        VN2CN2_sign => VN_sign_out(1874),
        VN2CN3_sign => VN_sign_out(1875),
        VN2CN4_sign => VN_sign_out(1876),
        VN2CN5_sign => VN_sign_out(1877),
        codeword => codeword(312),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN313 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1883 downto 1878),
        Din0 => VN313_in0,
        Din1 => VN313_in1,
        Din2 => VN313_in2,
        Din3 => VN313_in3,
        Din4 => VN313_in4,
        Din5 => VN313_in5,
        VN2CN0_bit => VN_data_out(1878),
        VN2CN1_bit => VN_data_out(1879),
        VN2CN2_bit => VN_data_out(1880),
        VN2CN3_bit => VN_data_out(1881),
        VN2CN4_bit => VN_data_out(1882),
        VN2CN5_bit => VN_data_out(1883),
        VN2CN0_sign => VN_sign_out(1878),
        VN2CN1_sign => VN_sign_out(1879),
        VN2CN2_sign => VN_sign_out(1880),
        VN2CN3_sign => VN_sign_out(1881),
        VN2CN4_sign => VN_sign_out(1882),
        VN2CN5_sign => VN_sign_out(1883),
        codeword => codeword(313),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN314 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1889 downto 1884),
        Din0 => VN314_in0,
        Din1 => VN314_in1,
        Din2 => VN314_in2,
        Din3 => VN314_in3,
        Din4 => VN314_in4,
        Din5 => VN314_in5,
        VN2CN0_bit => VN_data_out(1884),
        VN2CN1_bit => VN_data_out(1885),
        VN2CN2_bit => VN_data_out(1886),
        VN2CN3_bit => VN_data_out(1887),
        VN2CN4_bit => VN_data_out(1888),
        VN2CN5_bit => VN_data_out(1889),
        VN2CN0_sign => VN_sign_out(1884),
        VN2CN1_sign => VN_sign_out(1885),
        VN2CN2_sign => VN_sign_out(1886),
        VN2CN3_sign => VN_sign_out(1887),
        VN2CN4_sign => VN_sign_out(1888),
        VN2CN5_sign => VN_sign_out(1889),
        codeword => codeword(314),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN315 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1895 downto 1890),
        Din0 => VN315_in0,
        Din1 => VN315_in1,
        Din2 => VN315_in2,
        Din3 => VN315_in3,
        Din4 => VN315_in4,
        Din5 => VN315_in5,
        VN2CN0_bit => VN_data_out(1890),
        VN2CN1_bit => VN_data_out(1891),
        VN2CN2_bit => VN_data_out(1892),
        VN2CN3_bit => VN_data_out(1893),
        VN2CN4_bit => VN_data_out(1894),
        VN2CN5_bit => VN_data_out(1895),
        VN2CN0_sign => VN_sign_out(1890),
        VN2CN1_sign => VN_sign_out(1891),
        VN2CN2_sign => VN_sign_out(1892),
        VN2CN3_sign => VN_sign_out(1893),
        VN2CN4_sign => VN_sign_out(1894),
        VN2CN5_sign => VN_sign_out(1895),
        codeword => codeword(315),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN316 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1901 downto 1896),
        Din0 => VN316_in0,
        Din1 => VN316_in1,
        Din2 => VN316_in2,
        Din3 => VN316_in3,
        Din4 => VN316_in4,
        Din5 => VN316_in5,
        VN2CN0_bit => VN_data_out(1896),
        VN2CN1_bit => VN_data_out(1897),
        VN2CN2_bit => VN_data_out(1898),
        VN2CN3_bit => VN_data_out(1899),
        VN2CN4_bit => VN_data_out(1900),
        VN2CN5_bit => VN_data_out(1901),
        VN2CN0_sign => VN_sign_out(1896),
        VN2CN1_sign => VN_sign_out(1897),
        VN2CN2_sign => VN_sign_out(1898),
        VN2CN3_sign => VN_sign_out(1899),
        VN2CN4_sign => VN_sign_out(1900),
        VN2CN5_sign => VN_sign_out(1901),
        codeword => codeword(316),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN317 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1907 downto 1902),
        Din0 => VN317_in0,
        Din1 => VN317_in1,
        Din2 => VN317_in2,
        Din3 => VN317_in3,
        Din4 => VN317_in4,
        Din5 => VN317_in5,
        VN2CN0_bit => VN_data_out(1902),
        VN2CN1_bit => VN_data_out(1903),
        VN2CN2_bit => VN_data_out(1904),
        VN2CN3_bit => VN_data_out(1905),
        VN2CN4_bit => VN_data_out(1906),
        VN2CN5_bit => VN_data_out(1907),
        VN2CN0_sign => VN_sign_out(1902),
        VN2CN1_sign => VN_sign_out(1903),
        VN2CN2_sign => VN_sign_out(1904),
        VN2CN3_sign => VN_sign_out(1905),
        VN2CN4_sign => VN_sign_out(1906),
        VN2CN5_sign => VN_sign_out(1907),
        codeword => codeword(317),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN318 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1913 downto 1908),
        Din0 => VN318_in0,
        Din1 => VN318_in1,
        Din2 => VN318_in2,
        Din3 => VN318_in3,
        Din4 => VN318_in4,
        Din5 => VN318_in5,
        VN2CN0_bit => VN_data_out(1908),
        VN2CN1_bit => VN_data_out(1909),
        VN2CN2_bit => VN_data_out(1910),
        VN2CN3_bit => VN_data_out(1911),
        VN2CN4_bit => VN_data_out(1912),
        VN2CN5_bit => VN_data_out(1913),
        VN2CN0_sign => VN_sign_out(1908),
        VN2CN1_sign => VN_sign_out(1909),
        VN2CN2_sign => VN_sign_out(1910),
        VN2CN3_sign => VN_sign_out(1911),
        VN2CN4_sign => VN_sign_out(1912),
        VN2CN5_sign => VN_sign_out(1913),
        codeword => codeword(318),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN319 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1919 downto 1914),
        Din0 => VN319_in0,
        Din1 => VN319_in1,
        Din2 => VN319_in2,
        Din3 => VN319_in3,
        Din4 => VN319_in4,
        Din5 => VN319_in5,
        VN2CN0_bit => VN_data_out(1914),
        VN2CN1_bit => VN_data_out(1915),
        VN2CN2_bit => VN_data_out(1916),
        VN2CN3_bit => VN_data_out(1917),
        VN2CN4_bit => VN_data_out(1918),
        VN2CN5_bit => VN_data_out(1919),
        VN2CN0_sign => VN_sign_out(1914),
        VN2CN1_sign => VN_sign_out(1915),
        VN2CN2_sign => VN_sign_out(1916),
        VN2CN3_sign => VN_sign_out(1917),
        VN2CN4_sign => VN_sign_out(1918),
        VN2CN5_sign => VN_sign_out(1919),
        codeword => codeword(319),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN320 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1925 downto 1920),
        Din0 => VN320_in0,
        Din1 => VN320_in1,
        Din2 => VN320_in2,
        Din3 => VN320_in3,
        Din4 => VN320_in4,
        Din5 => VN320_in5,
        VN2CN0_bit => VN_data_out(1920),
        VN2CN1_bit => VN_data_out(1921),
        VN2CN2_bit => VN_data_out(1922),
        VN2CN3_bit => VN_data_out(1923),
        VN2CN4_bit => VN_data_out(1924),
        VN2CN5_bit => VN_data_out(1925),
        VN2CN0_sign => VN_sign_out(1920),
        VN2CN1_sign => VN_sign_out(1921),
        VN2CN2_sign => VN_sign_out(1922),
        VN2CN3_sign => VN_sign_out(1923),
        VN2CN4_sign => VN_sign_out(1924),
        VN2CN5_sign => VN_sign_out(1925),
        codeword => codeword(320),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN321 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1931 downto 1926),
        Din0 => VN321_in0,
        Din1 => VN321_in1,
        Din2 => VN321_in2,
        Din3 => VN321_in3,
        Din4 => VN321_in4,
        Din5 => VN321_in5,
        VN2CN0_bit => VN_data_out(1926),
        VN2CN1_bit => VN_data_out(1927),
        VN2CN2_bit => VN_data_out(1928),
        VN2CN3_bit => VN_data_out(1929),
        VN2CN4_bit => VN_data_out(1930),
        VN2CN5_bit => VN_data_out(1931),
        VN2CN0_sign => VN_sign_out(1926),
        VN2CN1_sign => VN_sign_out(1927),
        VN2CN2_sign => VN_sign_out(1928),
        VN2CN3_sign => VN_sign_out(1929),
        VN2CN4_sign => VN_sign_out(1930),
        VN2CN5_sign => VN_sign_out(1931),
        codeword => codeword(321),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN322 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1937 downto 1932),
        Din0 => VN322_in0,
        Din1 => VN322_in1,
        Din2 => VN322_in2,
        Din3 => VN322_in3,
        Din4 => VN322_in4,
        Din5 => VN322_in5,
        VN2CN0_bit => VN_data_out(1932),
        VN2CN1_bit => VN_data_out(1933),
        VN2CN2_bit => VN_data_out(1934),
        VN2CN3_bit => VN_data_out(1935),
        VN2CN4_bit => VN_data_out(1936),
        VN2CN5_bit => VN_data_out(1937),
        VN2CN0_sign => VN_sign_out(1932),
        VN2CN1_sign => VN_sign_out(1933),
        VN2CN2_sign => VN_sign_out(1934),
        VN2CN3_sign => VN_sign_out(1935),
        VN2CN4_sign => VN_sign_out(1936),
        VN2CN5_sign => VN_sign_out(1937),
        codeword => codeword(322),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN323 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1943 downto 1938),
        Din0 => VN323_in0,
        Din1 => VN323_in1,
        Din2 => VN323_in2,
        Din3 => VN323_in3,
        Din4 => VN323_in4,
        Din5 => VN323_in5,
        VN2CN0_bit => VN_data_out(1938),
        VN2CN1_bit => VN_data_out(1939),
        VN2CN2_bit => VN_data_out(1940),
        VN2CN3_bit => VN_data_out(1941),
        VN2CN4_bit => VN_data_out(1942),
        VN2CN5_bit => VN_data_out(1943),
        VN2CN0_sign => VN_sign_out(1938),
        VN2CN1_sign => VN_sign_out(1939),
        VN2CN2_sign => VN_sign_out(1940),
        VN2CN3_sign => VN_sign_out(1941),
        VN2CN4_sign => VN_sign_out(1942),
        VN2CN5_sign => VN_sign_out(1943),
        codeword => codeword(323),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN324 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1949 downto 1944),
        Din0 => VN324_in0,
        Din1 => VN324_in1,
        Din2 => VN324_in2,
        Din3 => VN324_in3,
        Din4 => VN324_in4,
        Din5 => VN324_in5,
        VN2CN0_bit => VN_data_out(1944),
        VN2CN1_bit => VN_data_out(1945),
        VN2CN2_bit => VN_data_out(1946),
        VN2CN3_bit => VN_data_out(1947),
        VN2CN4_bit => VN_data_out(1948),
        VN2CN5_bit => VN_data_out(1949),
        VN2CN0_sign => VN_sign_out(1944),
        VN2CN1_sign => VN_sign_out(1945),
        VN2CN2_sign => VN_sign_out(1946),
        VN2CN3_sign => VN_sign_out(1947),
        VN2CN4_sign => VN_sign_out(1948),
        VN2CN5_sign => VN_sign_out(1949),
        codeword => codeword(324),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN325 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1955 downto 1950),
        Din0 => VN325_in0,
        Din1 => VN325_in1,
        Din2 => VN325_in2,
        Din3 => VN325_in3,
        Din4 => VN325_in4,
        Din5 => VN325_in5,
        VN2CN0_bit => VN_data_out(1950),
        VN2CN1_bit => VN_data_out(1951),
        VN2CN2_bit => VN_data_out(1952),
        VN2CN3_bit => VN_data_out(1953),
        VN2CN4_bit => VN_data_out(1954),
        VN2CN5_bit => VN_data_out(1955),
        VN2CN0_sign => VN_sign_out(1950),
        VN2CN1_sign => VN_sign_out(1951),
        VN2CN2_sign => VN_sign_out(1952),
        VN2CN3_sign => VN_sign_out(1953),
        VN2CN4_sign => VN_sign_out(1954),
        VN2CN5_sign => VN_sign_out(1955),
        codeword => codeword(325),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN326 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1961 downto 1956),
        Din0 => VN326_in0,
        Din1 => VN326_in1,
        Din2 => VN326_in2,
        Din3 => VN326_in3,
        Din4 => VN326_in4,
        Din5 => VN326_in5,
        VN2CN0_bit => VN_data_out(1956),
        VN2CN1_bit => VN_data_out(1957),
        VN2CN2_bit => VN_data_out(1958),
        VN2CN3_bit => VN_data_out(1959),
        VN2CN4_bit => VN_data_out(1960),
        VN2CN5_bit => VN_data_out(1961),
        VN2CN0_sign => VN_sign_out(1956),
        VN2CN1_sign => VN_sign_out(1957),
        VN2CN2_sign => VN_sign_out(1958),
        VN2CN3_sign => VN_sign_out(1959),
        VN2CN4_sign => VN_sign_out(1960),
        VN2CN5_sign => VN_sign_out(1961),
        codeword => codeword(326),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN327 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1967 downto 1962),
        Din0 => VN327_in0,
        Din1 => VN327_in1,
        Din2 => VN327_in2,
        Din3 => VN327_in3,
        Din4 => VN327_in4,
        Din5 => VN327_in5,
        VN2CN0_bit => VN_data_out(1962),
        VN2CN1_bit => VN_data_out(1963),
        VN2CN2_bit => VN_data_out(1964),
        VN2CN3_bit => VN_data_out(1965),
        VN2CN4_bit => VN_data_out(1966),
        VN2CN5_bit => VN_data_out(1967),
        VN2CN0_sign => VN_sign_out(1962),
        VN2CN1_sign => VN_sign_out(1963),
        VN2CN2_sign => VN_sign_out(1964),
        VN2CN3_sign => VN_sign_out(1965),
        VN2CN4_sign => VN_sign_out(1966),
        VN2CN5_sign => VN_sign_out(1967),
        codeword => codeword(327),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN328 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1973 downto 1968),
        Din0 => VN328_in0,
        Din1 => VN328_in1,
        Din2 => VN328_in2,
        Din3 => VN328_in3,
        Din4 => VN328_in4,
        Din5 => VN328_in5,
        VN2CN0_bit => VN_data_out(1968),
        VN2CN1_bit => VN_data_out(1969),
        VN2CN2_bit => VN_data_out(1970),
        VN2CN3_bit => VN_data_out(1971),
        VN2CN4_bit => VN_data_out(1972),
        VN2CN5_bit => VN_data_out(1973),
        VN2CN0_sign => VN_sign_out(1968),
        VN2CN1_sign => VN_sign_out(1969),
        VN2CN2_sign => VN_sign_out(1970),
        VN2CN3_sign => VN_sign_out(1971),
        VN2CN4_sign => VN_sign_out(1972),
        VN2CN5_sign => VN_sign_out(1973),
        codeword => codeword(328),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN329 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1979 downto 1974),
        Din0 => VN329_in0,
        Din1 => VN329_in1,
        Din2 => VN329_in2,
        Din3 => VN329_in3,
        Din4 => VN329_in4,
        Din5 => VN329_in5,
        VN2CN0_bit => VN_data_out(1974),
        VN2CN1_bit => VN_data_out(1975),
        VN2CN2_bit => VN_data_out(1976),
        VN2CN3_bit => VN_data_out(1977),
        VN2CN4_bit => VN_data_out(1978),
        VN2CN5_bit => VN_data_out(1979),
        VN2CN0_sign => VN_sign_out(1974),
        VN2CN1_sign => VN_sign_out(1975),
        VN2CN2_sign => VN_sign_out(1976),
        VN2CN3_sign => VN_sign_out(1977),
        VN2CN4_sign => VN_sign_out(1978),
        VN2CN5_sign => VN_sign_out(1979),
        codeword => codeword(329),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN330 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1985 downto 1980),
        Din0 => VN330_in0,
        Din1 => VN330_in1,
        Din2 => VN330_in2,
        Din3 => VN330_in3,
        Din4 => VN330_in4,
        Din5 => VN330_in5,
        VN2CN0_bit => VN_data_out(1980),
        VN2CN1_bit => VN_data_out(1981),
        VN2CN2_bit => VN_data_out(1982),
        VN2CN3_bit => VN_data_out(1983),
        VN2CN4_bit => VN_data_out(1984),
        VN2CN5_bit => VN_data_out(1985),
        VN2CN0_sign => VN_sign_out(1980),
        VN2CN1_sign => VN_sign_out(1981),
        VN2CN2_sign => VN_sign_out(1982),
        VN2CN3_sign => VN_sign_out(1983),
        VN2CN4_sign => VN_sign_out(1984),
        VN2CN5_sign => VN_sign_out(1985),
        codeword => codeword(330),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN331 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1991 downto 1986),
        Din0 => VN331_in0,
        Din1 => VN331_in1,
        Din2 => VN331_in2,
        Din3 => VN331_in3,
        Din4 => VN331_in4,
        Din5 => VN331_in5,
        VN2CN0_bit => VN_data_out(1986),
        VN2CN1_bit => VN_data_out(1987),
        VN2CN2_bit => VN_data_out(1988),
        VN2CN3_bit => VN_data_out(1989),
        VN2CN4_bit => VN_data_out(1990),
        VN2CN5_bit => VN_data_out(1991),
        VN2CN0_sign => VN_sign_out(1986),
        VN2CN1_sign => VN_sign_out(1987),
        VN2CN2_sign => VN_sign_out(1988),
        VN2CN3_sign => VN_sign_out(1989),
        VN2CN4_sign => VN_sign_out(1990),
        VN2CN5_sign => VN_sign_out(1991),
        codeword => codeword(331),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN332 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(1997 downto 1992),
        Din0 => VN332_in0,
        Din1 => VN332_in1,
        Din2 => VN332_in2,
        Din3 => VN332_in3,
        Din4 => VN332_in4,
        Din5 => VN332_in5,
        VN2CN0_bit => VN_data_out(1992),
        VN2CN1_bit => VN_data_out(1993),
        VN2CN2_bit => VN_data_out(1994),
        VN2CN3_bit => VN_data_out(1995),
        VN2CN4_bit => VN_data_out(1996),
        VN2CN5_bit => VN_data_out(1997),
        VN2CN0_sign => VN_sign_out(1992),
        VN2CN1_sign => VN_sign_out(1993),
        VN2CN2_sign => VN_sign_out(1994),
        VN2CN3_sign => VN_sign_out(1995),
        VN2CN4_sign => VN_sign_out(1996),
        VN2CN5_sign => VN_sign_out(1997),
        codeword => codeword(332),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN333 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2003 downto 1998),
        Din0 => VN333_in0,
        Din1 => VN333_in1,
        Din2 => VN333_in2,
        Din3 => VN333_in3,
        Din4 => VN333_in4,
        Din5 => VN333_in5,
        VN2CN0_bit => VN_data_out(1998),
        VN2CN1_bit => VN_data_out(1999),
        VN2CN2_bit => VN_data_out(2000),
        VN2CN3_bit => VN_data_out(2001),
        VN2CN4_bit => VN_data_out(2002),
        VN2CN5_bit => VN_data_out(2003),
        VN2CN0_sign => VN_sign_out(1998),
        VN2CN1_sign => VN_sign_out(1999),
        VN2CN2_sign => VN_sign_out(2000),
        VN2CN3_sign => VN_sign_out(2001),
        VN2CN4_sign => VN_sign_out(2002),
        VN2CN5_sign => VN_sign_out(2003),
        codeword => codeword(333),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN334 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2009 downto 2004),
        Din0 => VN334_in0,
        Din1 => VN334_in1,
        Din2 => VN334_in2,
        Din3 => VN334_in3,
        Din4 => VN334_in4,
        Din5 => VN334_in5,
        VN2CN0_bit => VN_data_out(2004),
        VN2CN1_bit => VN_data_out(2005),
        VN2CN2_bit => VN_data_out(2006),
        VN2CN3_bit => VN_data_out(2007),
        VN2CN4_bit => VN_data_out(2008),
        VN2CN5_bit => VN_data_out(2009),
        VN2CN0_sign => VN_sign_out(2004),
        VN2CN1_sign => VN_sign_out(2005),
        VN2CN2_sign => VN_sign_out(2006),
        VN2CN3_sign => VN_sign_out(2007),
        VN2CN4_sign => VN_sign_out(2008),
        VN2CN5_sign => VN_sign_out(2009),
        codeword => codeword(334),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN335 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2015 downto 2010),
        Din0 => VN335_in0,
        Din1 => VN335_in1,
        Din2 => VN335_in2,
        Din3 => VN335_in3,
        Din4 => VN335_in4,
        Din5 => VN335_in5,
        VN2CN0_bit => VN_data_out(2010),
        VN2CN1_bit => VN_data_out(2011),
        VN2CN2_bit => VN_data_out(2012),
        VN2CN3_bit => VN_data_out(2013),
        VN2CN4_bit => VN_data_out(2014),
        VN2CN5_bit => VN_data_out(2015),
        VN2CN0_sign => VN_sign_out(2010),
        VN2CN1_sign => VN_sign_out(2011),
        VN2CN2_sign => VN_sign_out(2012),
        VN2CN3_sign => VN_sign_out(2013),
        VN2CN4_sign => VN_sign_out(2014),
        VN2CN5_sign => VN_sign_out(2015),
        codeword => codeword(335),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN336 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2021 downto 2016),
        Din0 => VN336_in0,
        Din1 => VN336_in1,
        Din2 => VN336_in2,
        Din3 => VN336_in3,
        Din4 => VN336_in4,
        Din5 => VN336_in5,
        VN2CN0_bit => VN_data_out(2016),
        VN2CN1_bit => VN_data_out(2017),
        VN2CN2_bit => VN_data_out(2018),
        VN2CN3_bit => VN_data_out(2019),
        VN2CN4_bit => VN_data_out(2020),
        VN2CN5_bit => VN_data_out(2021),
        VN2CN0_sign => VN_sign_out(2016),
        VN2CN1_sign => VN_sign_out(2017),
        VN2CN2_sign => VN_sign_out(2018),
        VN2CN3_sign => VN_sign_out(2019),
        VN2CN4_sign => VN_sign_out(2020),
        VN2CN5_sign => VN_sign_out(2021),
        codeword => codeword(336),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN337 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2027 downto 2022),
        Din0 => VN337_in0,
        Din1 => VN337_in1,
        Din2 => VN337_in2,
        Din3 => VN337_in3,
        Din4 => VN337_in4,
        Din5 => VN337_in5,
        VN2CN0_bit => VN_data_out(2022),
        VN2CN1_bit => VN_data_out(2023),
        VN2CN2_bit => VN_data_out(2024),
        VN2CN3_bit => VN_data_out(2025),
        VN2CN4_bit => VN_data_out(2026),
        VN2CN5_bit => VN_data_out(2027),
        VN2CN0_sign => VN_sign_out(2022),
        VN2CN1_sign => VN_sign_out(2023),
        VN2CN2_sign => VN_sign_out(2024),
        VN2CN3_sign => VN_sign_out(2025),
        VN2CN4_sign => VN_sign_out(2026),
        VN2CN5_sign => VN_sign_out(2027),
        codeword => codeword(337),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN338 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2033 downto 2028),
        Din0 => VN338_in0,
        Din1 => VN338_in1,
        Din2 => VN338_in2,
        Din3 => VN338_in3,
        Din4 => VN338_in4,
        Din5 => VN338_in5,
        VN2CN0_bit => VN_data_out(2028),
        VN2CN1_bit => VN_data_out(2029),
        VN2CN2_bit => VN_data_out(2030),
        VN2CN3_bit => VN_data_out(2031),
        VN2CN4_bit => VN_data_out(2032),
        VN2CN5_bit => VN_data_out(2033),
        VN2CN0_sign => VN_sign_out(2028),
        VN2CN1_sign => VN_sign_out(2029),
        VN2CN2_sign => VN_sign_out(2030),
        VN2CN3_sign => VN_sign_out(2031),
        VN2CN4_sign => VN_sign_out(2032),
        VN2CN5_sign => VN_sign_out(2033),
        codeword => codeword(338),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN339 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2039 downto 2034),
        Din0 => VN339_in0,
        Din1 => VN339_in1,
        Din2 => VN339_in2,
        Din3 => VN339_in3,
        Din4 => VN339_in4,
        Din5 => VN339_in5,
        VN2CN0_bit => VN_data_out(2034),
        VN2CN1_bit => VN_data_out(2035),
        VN2CN2_bit => VN_data_out(2036),
        VN2CN3_bit => VN_data_out(2037),
        VN2CN4_bit => VN_data_out(2038),
        VN2CN5_bit => VN_data_out(2039),
        VN2CN0_sign => VN_sign_out(2034),
        VN2CN1_sign => VN_sign_out(2035),
        VN2CN2_sign => VN_sign_out(2036),
        VN2CN3_sign => VN_sign_out(2037),
        VN2CN4_sign => VN_sign_out(2038),
        VN2CN5_sign => VN_sign_out(2039),
        codeword => codeword(339),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN340 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2045 downto 2040),
        Din0 => VN340_in0,
        Din1 => VN340_in1,
        Din2 => VN340_in2,
        Din3 => VN340_in3,
        Din4 => VN340_in4,
        Din5 => VN340_in5,
        VN2CN0_bit => VN_data_out(2040),
        VN2CN1_bit => VN_data_out(2041),
        VN2CN2_bit => VN_data_out(2042),
        VN2CN3_bit => VN_data_out(2043),
        VN2CN4_bit => VN_data_out(2044),
        VN2CN5_bit => VN_data_out(2045),
        VN2CN0_sign => VN_sign_out(2040),
        VN2CN1_sign => VN_sign_out(2041),
        VN2CN2_sign => VN_sign_out(2042),
        VN2CN3_sign => VN_sign_out(2043),
        VN2CN4_sign => VN_sign_out(2044),
        VN2CN5_sign => VN_sign_out(2045),
        codeword => codeword(340),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN341 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2051 downto 2046),
        Din0 => VN341_in0,
        Din1 => VN341_in1,
        Din2 => VN341_in2,
        Din3 => VN341_in3,
        Din4 => VN341_in4,
        Din5 => VN341_in5,
        VN2CN0_bit => VN_data_out(2046),
        VN2CN1_bit => VN_data_out(2047),
        VN2CN2_bit => VN_data_out(2048),
        VN2CN3_bit => VN_data_out(2049),
        VN2CN4_bit => VN_data_out(2050),
        VN2CN5_bit => VN_data_out(2051),
        VN2CN0_sign => VN_sign_out(2046),
        VN2CN1_sign => VN_sign_out(2047),
        VN2CN2_sign => VN_sign_out(2048),
        VN2CN3_sign => VN_sign_out(2049),
        VN2CN4_sign => VN_sign_out(2050),
        VN2CN5_sign => VN_sign_out(2051),
        codeword => codeword(341),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN342 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2057 downto 2052),
        Din0 => VN342_in0,
        Din1 => VN342_in1,
        Din2 => VN342_in2,
        Din3 => VN342_in3,
        Din4 => VN342_in4,
        Din5 => VN342_in5,
        VN2CN0_bit => VN_data_out(2052),
        VN2CN1_bit => VN_data_out(2053),
        VN2CN2_bit => VN_data_out(2054),
        VN2CN3_bit => VN_data_out(2055),
        VN2CN4_bit => VN_data_out(2056),
        VN2CN5_bit => VN_data_out(2057),
        VN2CN0_sign => VN_sign_out(2052),
        VN2CN1_sign => VN_sign_out(2053),
        VN2CN2_sign => VN_sign_out(2054),
        VN2CN3_sign => VN_sign_out(2055),
        VN2CN4_sign => VN_sign_out(2056),
        VN2CN5_sign => VN_sign_out(2057),
        codeword => codeword(342),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN343 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2063 downto 2058),
        Din0 => VN343_in0,
        Din1 => VN343_in1,
        Din2 => VN343_in2,
        Din3 => VN343_in3,
        Din4 => VN343_in4,
        Din5 => VN343_in5,
        VN2CN0_bit => VN_data_out(2058),
        VN2CN1_bit => VN_data_out(2059),
        VN2CN2_bit => VN_data_out(2060),
        VN2CN3_bit => VN_data_out(2061),
        VN2CN4_bit => VN_data_out(2062),
        VN2CN5_bit => VN_data_out(2063),
        VN2CN0_sign => VN_sign_out(2058),
        VN2CN1_sign => VN_sign_out(2059),
        VN2CN2_sign => VN_sign_out(2060),
        VN2CN3_sign => VN_sign_out(2061),
        VN2CN4_sign => VN_sign_out(2062),
        VN2CN5_sign => VN_sign_out(2063),
        codeword => codeword(343),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN344 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2069 downto 2064),
        Din0 => VN344_in0,
        Din1 => VN344_in1,
        Din2 => VN344_in2,
        Din3 => VN344_in3,
        Din4 => VN344_in4,
        Din5 => VN344_in5,
        VN2CN0_bit => VN_data_out(2064),
        VN2CN1_bit => VN_data_out(2065),
        VN2CN2_bit => VN_data_out(2066),
        VN2CN3_bit => VN_data_out(2067),
        VN2CN4_bit => VN_data_out(2068),
        VN2CN5_bit => VN_data_out(2069),
        VN2CN0_sign => VN_sign_out(2064),
        VN2CN1_sign => VN_sign_out(2065),
        VN2CN2_sign => VN_sign_out(2066),
        VN2CN3_sign => VN_sign_out(2067),
        VN2CN4_sign => VN_sign_out(2068),
        VN2CN5_sign => VN_sign_out(2069),
        codeword => codeword(344),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN345 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2075 downto 2070),
        Din0 => VN345_in0,
        Din1 => VN345_in1,
        Din2 => VN345_in2,
        Din3 => VN345_in3,
        Din4 => VN345_in4,
        Din5 => VN345_in5,
        VN2CN0_bit => VN_data_out(2070),
        VN2CN1_bit => VN_data_out(2071),
        VN2CN2_bit => VN_data_out(2072),
        VN2CN3_bit => VN_data_out(2073),
        VN2CN4_bit => VN_data_out(2074),
        VN2CN5_bit => VN_data_out(2075),
        VN2CN0_sign => VN_sign_out(2070),
        VN2CN1_sign => VN_sign_out(2071),
        VN2CN2_sign => VN_sign_out(2072),
        VN2CN3_sign => VN_sign_out(2073),
        VN2CN4_sign => VN_sign_out(2074),
        VN2CN5_sign => VN_sign_out(2075),
        codeword => codeword(345),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN346 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2081 downto 2076),
        Din0 => VN346_in0,
        Din1 => VN346_in1,
        Din2 => VN346_in2,
        Din3 => VN346_in3,
        Din4 => VN346_in4,
        Din5 => VN346_in5,
        VN2CN0_bit => VN_data_out(2076),
        VN2CN1_bit => VN_data_out(2077),
        VN2CN2_bit => VN_data_out(2078),
        VN2CN3_bit => VN_data_out(2079),
        VN2CN4_bit => VN_data_out(2080),
        VN2CN5_bit => VN_data_out(2081),
        VN2CN0_sign => VN_sign_out(2076),
        VN2CN1_sign => VN_sign_out(2077),
        VN2CN2_sign => VN_sign_out(2078),
        VN2CN3_sign => VN_sign_out(2079),
        VN2CN4_sign => VN_sign_out(2080),
        VN2CN5_sign => VN_sign_out(2081),
        codeword => codeword(346),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN347 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2087 downto 2082),
        Din0 => VN347_in0,
        Din1 => VN347_in1,
        Din2 => VN347_in2,
        Din3 => VN347_in3,
        Din4 => VN347_in4,
        Din5 => VN347_in5,
        VN2CN0_bit => VN_data_out(2082),
        VN2CN1_bit => VN_data_out(2083),
        VN2CN2_bit => VN_data_out(2084),
        VN2CN3_bit => VN_data_out(2085),
        VN2CN4_bit => VN_data_out(2086),
        VN2CN5_bit => VN_data_out(2087),
        VN2CN0_sign => VN_sign_out(2082),
        VN2CN1_sign => VN_sign_out(2083),
        VN2CN2_sign => VN_sign_out(2084),
        VN2CN3_sign => VN_sign_out(2085),
        VN2CN4_sign => VN_sign_out(2086),
        VN2CN5_sign => VN_sign_out(2087),
        codeword => codeword(347),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN348 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2093 downto 2088),
        Din0 => VN348_in0,
        Din1 => VN348_in1,
        Din2 => VN348_in2,
        Din3 => VN348_in3,
        Din4 => VN348_in4,
        Din5 => VN348_in5,
        VN2CN0_bit => VN_data_out(2088),
        VN2CN1_bit => VN_data_out(2089),
        VN2CN2_bit => VN_data_out(2090),
        VN2CN3_bit => VN_data_out(2091),
        VN2CN4_bit => VN_data_out(2092),
        VN2CN5_bit => VN_data_out(2093),
        VN2CN0_sign => VN_sign_out(2088),
        VN2CN1_sign => VN_sign_out(2089),
        VN2CN2_sign => VN_sign_out(2090),
        VN2CN3_sign => VN_sign_out(2091),
        VN2CN4_sign => VN_sign_out(2092),
        VN2CN5_sign => VN_sign_out(2093),
        codeword => codeword(348),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN349 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2099 downto 2094),
        Din0 => VN349_in0,
        Din1 => VN349_in1,
        Din2 => VN349_in2,
        Din3 => VN349_in3,
        Din4 => VN349_in4,
        Din5 => VN349_in5,
        VN2CN0_bit => VN_data_out(2094),
        VN2CN1_bit => VN_data_out(2095),
        VN2CN2_bit => VN_data_out(2096),
        VN2CN3_bit => VN_data_out(2097),
        VN2CN4_bit => VN_data_out(2098),
        VN2CN5_bit => VN_data_out(2099),
        VN2CN0_sign => VN_sign_out(2094),
        VN2CN1_sign => VN_sign_out(2095),
        VN2CN2_sign => VN_sign_out(2096),
        VN2CN3_sign => VN_sign_out(2097),
        VN2CN4_sign => VN_sign_out(2098),
        VN2CN5_sign => VN_sign_out(2099),
        codeword => codeword(349),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN350 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2105 downto 2100),
        Din0 => VN350_in0,
        Din1 => VN350_in1,
        Din2 => VN350_in2,
        Din3 => VN350_in3,
        Din4 => VN350_in4,
        Din5 => VN350_in5,
        VN2CN0_bit => VN_data_out(2100),
        VN2CN1_bit => VN_data_out(2101),
        VN2CN2_bit => VN_data_out(2102),
        VN2CN3_bit => VN_data_out(2103),
        VN2CN4_bit => VN_data_out(2104),
        VN2CN5_bit => VN_data_out(2105),
        VN2CN0_sign => VN_sign_out(2100),
        VN2CN1_sign => VN_sign_out(2101),
        VN2CN2_sign => VN_sign_out(2102),
        VN2CN3_sign => VN_sign_out(2103),
        VN2CN4_sign => VN_sign_out(2104),
        VN2CN5_sign => VN_sign_out(2105),
        codeword => codeword(350),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN351 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2111 downto 2106),
        Din0 => VN351_in0,
        Din1 => VN351_in1,
        Din2 => VN351_in2,
        Din3 => VN351_in3,
        Din4 => VN351_in4,
        Din5 => VN351_in5,
        VN2CN0_bit => VN_data_out(2106),
        VN2CN1_bit => VN_data_out(2107),
        VN2CN2_bit => VN_data_out(2108),
        VN2CN3_bit => VN_data_out(2109),
        VN2CN4_bit => VN_data_out(2110),
        VN2CN5_bit => VN_data_out(2111),
        VN2CN0_sign => VN_sign_out(2106),
        VN2CN1_sign => VN_sign_out(2107),
        VN2CN2_sign => VN_sign_out(2108),
        VN2CN3_sign => VN_sign_out(2109),
        VN2CN4_sign => VN_sign_out(2110),
        VN2CN5_sign => VN_sign_out(2111),
        codeword => codeword(351),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN352 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2117 downto 2112),
        Din0 => VN352_in0,
        Din1 => VN352_in1,
        Din2 => VN352_in2,
        Din3 => VN352_in3,
        Din4 => VN352_in4,
        Din5 => VN352_in5,
        VN2CN0_bit => VN_data_out(2112),
        VN2CN1_bit => VN_data_out(2113),
        VN2CN2_bit => VN_data_out(2114),
        VN2CN3_bit => VN_data_out(2115),
        VN2CN4_bit => VN_data_out(2116),
        VN2CN5_bit => VN_data_out(2117),
        VN2CN0_sign => VN_sign_out(2112),
        VN2CN1_sign => VN_sign_out(2113),
        VN2CN2_sign => VN_sign_out(2114),
        VN2CN3_sign => VN_sign_out(2115),
        VN2CN4_sign => VN_sign_out(2116),
        VN2CN5_sign => VN_sign_out(2117),
        codeword => codeword(352),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN353 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2123 downto 2118),
        Din0 => VN353_in0,
        Din1 => VN353_in1,
        Din2 => VN353_in2,
        Din3 => VN353_in3,
        Din4 => VN353_in4,
        Din5 => VN353_in5,
        VN2CN0_bit => VN_data_out(2118),
        VN2CN1_bit => VN_data_out(2119),
        VN2CN2_bit => VN_data_out(2120),
        VN2CN3_bit => VN_data_out(2121),
        VN2CN4_bit => VN_data_out(2122),
        VN2CN5_bit => VN_data_out(2123),
        VN2CN0_sign => VN_sign_out(2118),
        VN2CN1_sign => VN_sign_out(2119),
        VN2CN2_sign => VN_sign_out(2120),
        VN2CN3_sign => VN_sign_out(2121),
        VN2CN4_sign => VN_sign_out(2122),
        VN2CN5_sign => VN_sign_out(2123),
        codeword => codeword(353),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN354 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2129 downto 2124),
        Din0 => VN354_in0,
        Din1 => VN354_in1,
        Din2 => VN354_in2,
        Din3 => VN354_in3,
        Din4 => VN354_in4,
        Din5 => VN354_in5,
        VN2CN0_bit => VN_data_out(2124),
        VN2CN1_bit => VN_data_out(2125),
        VN2CN2_bit => VN_data_out(2126),
        VN2CN3_bit => VN_data_out(2127),
        VN2CN4_bit => VN_data_out(2128),
        VN2CN5_bit => VN_data_out(2129),
        VN2CN0_sign => VN_sign_out(2124),
        VN2CN1_sign => VN_sign_out(2125),
        VN2CN2_sign => VN_sign_out(2126),
        VN2CN3_sign => VN_sign_out(2127),
        VN2CN4_sign => VN_sign_out(2128),
        VN2CN5_sign => VN_sign_out(2129),
        codeword => codeword(354),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN355 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2135 downto 2130),
        Din0 => VN355_in0,
        Din1 => VN355_in1,
        Din2 => VN355_in2,
        Din3 => VN355_in3,
        Din4 => VN355_in4,
        Din5 => VN355_in5,
        VN2CN0_bit => VN_data_out(2130),
        VN2CN1_bit => VN_data_out(2131),
        VN2CN2_bit => VN_data_out(2132),
        VN2CN3_bit => VN_data_out(2133),
        VN2CN4_bit => VN_data_out(2134),
        VN2CN5_bit => VN_data_out(2135),
        VN2CN0_sign => VN_sign_out(2130),
        VN2CN1_sign => VN_sign_out(2131),
        VN2CN2_sign => VN_sign_out(2132),
        VN2CN3_sign => VN_sign_out(2133),
        VN2CN4_sign => VN_sign_out(2134),
        VN2CN5_sign => VN_sign_out(2135),
        codeword => codeword(355),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN356 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2141 downto 2136),
        Din0 => VN356_in0,
        Din1 => VN356_in1,
        Din2 => VN356_in2,
        Din3 => VN356_in3,
        Din4 => VN356_in4,
        Din5 => VN356_in5,
        VN2CN0_bit => VN_data_out(2136),
        VN2CN1_bit => VN_data_out(2137),
        VN2CN2_bit => VN_data_out(2138),
        VN2CN3_bit => VN_data_out(2139),
        VN2CN4_bit => VN_data_out(2140),
        VN2CN5_bit => VN_data_out(2141),
        VN2CN0_sign => VN_sign_out(2136),
        VN2CN1_sign => VN_sign_out(2137),
        VN2CN2_sign => VN_sign_out(2138),
        VN2CN3_sign => VN_sign_out(2139),
        VN2CN4_sign => VN_sign_out(2140),
        VN2CN5_sign => VN_sign_out(2141),
        codeword => codeword(356),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN357 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2147 downto 2142),
        Din0 => VN357_in0,
        Din1 => VN357_in1,
        Din2 => VN357_in2,
        Din3 => VN357_in3,
        Din4 => VN357_in4,
        Din5 => VN357_in5,
        VN2CN0_bit => VN_data_out(2142),
        VN2CN1_bit => VN_data_out(2143),
        VN2CN2_bit => VN_data_out(2144),
        VN2CN3_bit => VN_data_out(2145),
        VN2CN4_bit => VN_data_out(2146),
        VN2CN5_bit => VN_data_out(2147),
        VN2CN0_sign => VN_sign_out(2142),
        VN2CN1_sign => VN_sign_out(2143),
        VN2CN2_sign => VN_sign_out(2144),
        VN2CN3_sign => VN_sign_out(2145),
        VN2CN4_sign => VN_sign_out(2146),
        VN2CN5_sign => VN_sign_out(2147),
        codeword => codeword(357),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN358 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2153 downto 2148),
        Din0 => VN358_in0,
        Din1 => VN358_in1,
        Din2 => VN358_in2,
        Din3 => VN358_in3,
        Din4 => VN358_in4,
        Din5 => VN358_in5,
        VN2CN0_bit => VN_data_out(2148),
        VN2CN1_bit => VN_data_out(2149),
        VN2CN2_bit => VN_data_out(2150),
        VN2CN3_bit => VN_data_out(2151),
        VN2CN4_bit => VN_data_out(2152),
        VN2CN5_bit => VN_data_out(2153),
        VN2CN0_sign => VN_sign_out(2148),
        VN2CN1_sign => VN_sign_out(2149),
        VN2CN2_sign => VN_sign_out(2150),
        VN2CN3_sign => VN_sign_out(2151),
        VN2CN4_sign => VN_sign_out(2152),
        VN2CN5_sign => VN_sign_out(2153),
        codeword => codeword(358),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN359 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2159 downto 2154),
        Din0 => VN359_in0,
        Din1 => VN359_in1,
        Din2 => VN359_in2,
        Din3 => VN359_in3,
        Din4 => VN359_in4,
        Din5 => VN359_in5,
        VN2CN0_bit => VN_data_out(2154),
        VN2CN1_bit => VN_data_out(2155),
        VN2CN2_bit => VN_data_out(2156),
        VN2CN3_bit => VN_data_out(2157),
        VN2CN4_bit => VN_data_out(2158),
        VN2CN5_bit => VN_data_out(2159),
        VN2CN0_sign => VN_sign_out(2154),
        VN2CN1_sign => VN_sign_out(2155),
        VN2CN2_sign => VN_sign_out(2156),
        VN2CN3_sign => VN_sign_out(2157),
        VN2CN4_sign => VN_sign_out(2158),
        VN2CN5_sign => VN_sign_out(2159),
        codeword => codeword(359),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN360 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2165 downto 2160),
        Din0 => VN360_in0,
        Din1 => VN360_in1,
        Din2 => VN360_in2,
        Din3 => VN360_in3,
        Din4 => VN360_in4,
        Din5 => VN360_in5,
        VN2CN0_bit => VN_data_out(2160),
        VN2CN1_bit => VN_data_out(2161),
        VN2CN2_bit => VN_data_out(2162),
        VN2CN3_bit => VN_data_out(2163),
        VN2CN4_bit => VN_data_out(2164),
        VN2CN5_bit => VN_data_out(2165),
        VN2CN0_sign => VN_sign_out(2160),
        VN2CN1_sign => VN_sign_out(2161),
        VN2CN2_sign => VN_sign_out(2162),
        VN2CN3_sign => VN_sign_out(2163),
        VN2CN4_sign => VN_sign_out(2164),
        VN2CN5_sign => VN_sign_out(2165),
        codeword => codeword(360),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN361 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2171 downto 2166),
        Din0 => VN361_in0,
        Din1 => VN361_in1,
        Din2 => VN361_in2,
        Din3 => VN361_in3,
        Din4 => VN361_in4,
        Din5 => VN361_in5,
        VN2CN0_bit => VN_data_out(2166),
        VN2CN1_bit => VN_data_out(2167),
        VN2CN2_bit => VN_data_out(2168),
        VN2CN3_bit => VN_data_out(2169),
        VN2CN4_bit => VN_data_out(2170),
        VN2CN5_bit => VN_data_out(2171),
        VN2CN0_sign => VN_sign_out(2166),
        VN2CN1_sign => VN_sign_out(2167),
        VN2CN2_sign => VN_sign_out(2168),
        VN2CN3_sign => VN_sign_out(2169),
        VN2CN4_sign => VN_sign_out(2170),
        VN2CN5_sign => VN_sign_out(2171),
        codeword => codeword(361),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN362 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2177 downto 2172),
        Din0 => VN362_in0,
        Din1 => VN362_in1,
        Din2 => VN362_in2,
        Din3 => VN362_in3,
        Din4 => VN362_in4,
        Din5 => VN362_in5,
        VN2CN0_bit => VN_data_out(2172),
        VN2CN1_bit => VN_data_out(2173),
        VN2CN2_bit => VN_data_out(2174),
        VN2CN3_bit => VN_data_out(2175),
        VN2CN4_bit => VN_data_out(2176),
        VN2CN5_bit => VN_data_out(2177),
        VN2CN0_sign => VN_sign_out(2172),
        VN2CN1_sign => VN_sign_out(2173),
        VN2CN2_sign => VN_sign_out(2174),
        VN2CN3_sign => VN_sign_out(2175),
        VN2CN4_sign => VN_sign_out(2176),
        VN2CN5_sign => VN_sign_out(2177),
        codeword => codeword(362),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN363 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2183 downto 2178),
        Din0 => VN363_in0,
        Din1 => VN363_in1,
        Din2 => VN363_in2,
        Din3 => VN363_in3,
        Din4 => VN363_in4,
        Din5 => VN363_in5,
        VN2CN0_bit => VN_data_out(2178),
        VN2CN1_bit => VN_data_out(2179),
        VN2CN2_bit => VN_data_out(2180),
        VN2CN3_bit => VN_data_out(2181),
        VN2CN4_bit => VN_data_out(2182),
        VN2CN5_bit => VN_data_out(2183),
        VN2CN0_sign => VN_sign_out(2178),
        VN2CN1_sign => VN_sign_out(2179),
        VN2CN2_sign => VN_sign_out(2180),
        VN2CN3_sign => VN_sign_out(2181),
        VN2CN4_sign => VN_sign_out(2182),
        VN2CN5_sign => VN_sign_out(2183),
        codeword => codeword(363),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN364 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2189 downto 2184),
        Din0 => VN364_in0,
        Din1 => VN364_in1,
        Din2 => VN364_in2,
        Din3 => VN364_in3,
        Din4 => VN364_in4,
        Din5 => VN364_in5,
        VN2CN0_bit => VN_data_out(2184),
        VN2CN1_bit => VN_data_out(2185),
        VN2CN2_bit => VN_data_out(2186),
        VN2CN3_bit => VN_data_out(2187),
        VN2CN4_bit => VN_data_out(2188),
        VN2CN5_bit => VN_data_out(2189),
        VN2CN0_sign => VN_sign_out(2184),
        VN2CN1_sign => VN_sign_out(2185),
        VN2CN2_sign => VN_sign_out(2186),
        VN2CN3_sign => VN_sign_out(2187),
        VN2CN4_sign => VN_sign_out(2188),
        VN2CN5_sign => VN_sign_out(2189),
        codeword => codeword(364),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN365 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2195 downto 2190),
        Din0 => VN365_in0,
        Din1 => VN365_in1,
        Din2 => VN365_in2,
        Din3 => VN365_in3,
        Din4 => VN365_in4,
        Din5 => VN365_in5,
        VN2CN0_bit => VN_data_out(2190),
        VN2CN1_bit => VN_data_out(2191),
        VN2CN2_bit => VN_data_out(2192),
        VN2CN3_bit => VN_data_out(2193),
        VN2CN4_bit => VN_data_out(2194),
        VN2CN5_bit => VN_data_out(2195),
        VN2CN0_sign => VN_sign_out(2190),
        VN2CN1_sign => VN_sign_out(2191),
        VN2CN2_sign => VN_sign_out(2192),
        VN2CN3_sign => VN_sign_out(2193),
        VN2CN4_sign => VN_sign_out(2194),
        VN2CN5_sign => VN_sign_out(2195),
        codeword => codeword(365),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN366 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2201 downto 2196),
        Din0 => VN366_in0,
        Din1 => VN366_in1,
        Din2 => VN366_in2,
        Din3 => VN366_in3,
        Din4 => VN366_in4,
        Din5 => VN366_in5,
        VN2CN0_bit => VN_data_out(2196),
        VN2CN1_bit => VN_data_out(2197),
        VN2CN2_bit => VN_data_out(2198),
        VN2CN3_bit => VN_data_out(2199),
        VN2CN4_bit => VN_data_out(2200),
        VN2CN5_bit => VN_data_out(2201),
        VN2CN0_sign => VN_sign_out(2196),
        VN2CN1_sign => VN_sign_out(2197),
        VN2CN2_sign => VN_sign_out(2198),
        VN2CN3_sign => VN_sign_out(2199),
        VN2CN4_sign => VN_sign_out(2200),
        VN2CN5_sign => VN_sign_out(2201),
        codeword => codeword(366),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN367 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2207 downto 2202),
        Din0 => VN367_in0,
        Din1 => VN367_in1,
        Din2 => VN367_in2,
        Din3 => VN367_in3,
        Din4 => VN367_in4,
        Din5 => VN367_in5,
        VN2CN0_bit => VN_data_out(2202),
        VN2CN1_bit => VN_data_out(2203),
        VN2CN2_bit => VN_data_out(2204),
        VN2CN3_bit => VN_data_out(2205),
        VN2CN4_bit => VN_data_out(2206),
        VN2CN5_bit => VN_data_out(2207),
        VN2CN0_sign => VN_sign_out(2202),
        VN2CN1_sign => VN_sign_out(2203),
        VN2CN2_sign => VN_sign_out(2204),
        VN2CN3_sign => VN_sign_out(2205),
        VN2CN4_sign => VN_sign_out(2206),
        VN2CN5_sign => VN_sign_out(2207),
        codeword => codeword(367),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN368 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2213 downto 2208),
        Din0 => VN368_in0,
        Din1 => VN368_in1,
        Din2 => VN368_in2,
        Din3 => VN368_in3,
        Din4 => VN368_in4,
        Din5 => VN368_in5,
        VN2CN0_bit => VN_data_out(2208),
        VN2CN1_bit => VN_data_out(2209),
        VN2CN2_bit => VN_data_out(2210),
        VN2CN3_bit => VN_data_out(2211),
        VN2CN4_bit => VN_data_out(2212),
        VN2CN5_bit => VN_data_out(2213),
        VN2CN0_sign => VN_sign_out(2208),
        VN2CN1_sign => VN_sign_out(2209),
        VN2CN2_sign => VN_sign_out(2210),
        VN2CN3_sign => VN_sign_out(2211),
        VN2CN4_sign => VN_sign_out(2212),
        VN2CN5_sign => VN_sign_out(2213),
        codeword => codeword(368),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN369 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2219 downto 2214),
        Din0 => VN369_in0,
        Din1 => VN369_in1,
        Din2 => VN369_in2,
        Din3 => VN369_in3,
        Din4 => VN369_in4,
        Din5 => VN369_in5,
        VN2CN0_bit => VN_data_out(2214),
        VN2CN1_bit => VN_data_out(2215),
        VN2CN2_bit => VN_data_out(2216),
        VN2CN3_bit => VN_data_out(2217),
        VN2CN4_bit => VN_data_out(2218),
        VN2CN5_bit => VN_data_out(2219),
        VN2CN0_sign => VN_sign_out(2214),
        VN2CN1_sign => VN_sign_out(2215),
        VN2CN2_sign => VN_sign_out(2216),
        VN2CN3_sign => VN_sign_out(2217),
        VN2CN4_sign => VN_sign_out(2218),
        VN2CN5_sign => VN_sign_out(2219),
        codeword => codeword(369),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN370 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2225 downto 2220),
        Din0 => VN370_in0,
        Din1 => VN370_in1,
        Din2 => VN370_in2,
        Din3 => VN370_in3,
        Din4 => VN370_in4,
        Din5 => VN370_in5,
        VN2CN0_bit => VN_data_out(2220),
        VN2CN1_bit => VN_data_out(2221),
        VN2CN2_bit => VN_data_out(2222),
        VN2CN3_bit => VN_data_out(2223),
        VN2CN4_bit => VN_data_out(2224),
        VN2CN5_bit => VN_data_out(2225),
        VN2CN0_sign => VN_sign_out(2220),
        VN2CN1_sign => VN_sign_out(2221),
        VN2CN2_sign => VN_sign_out(2222),
        VN2CN3_sign => VN_sign_out(2223),
        VN2CN4_sign => VN_sign_out(2224),
        VN2CN5_sign => VN_sign_out(2225),
        codeword => codeword(370),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN371 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2231 downto 2226),
        Din0 => VN371_in0,
        Din1 => VN371_in1,
        Din2 => VN371_in2,
        Din3 => VN371_in3,
        Din4 => VN371_in4,
        Din5 => VN371_in5,
        VN2CN0_bit => VN_data_out(2226),
        VN2CN1_bit => VN_data_out(2227),
        VN2CN2_bit => VN_data_out(2228),
        VN2CN3_bit => VN_data_out(2229),
        VN2CN4_bit => VN_data_out(2230),
        VN2CN5_bit => VN_data_out(2231),
        VN2CN0_sign => VN_sign_out(2226),
        VN2CN1_sign => VN_sign_out(2227),
        VN2CN2_sign => VN_sign_out(2228),
        VN2CN3_sign => VN_sign_out(2229),
        VN2CN4_sign => VN_sign_out(2230),
        VN2CN5_sign => VN_sign_out(2231),
        codeword => codeword(371),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN372 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2237 downto 2232),
        Din0 => VN372_in0,
        Din1 => VN372_in1,
        Din2 => VN372_in2,
        Din3 => VN372_in3,
        Din4 => VN372_in4,
        Din5 => VN372_in5,
        VN2CN0_bit => VN_data_out(2232),
        VN2CN1_bit => VN_data_out(2233),
        VN2CN2_bit => VN_data_out(2234),
        VN2CN3_bit => VN_data_out(2235),
        VN2CN4_bit => VN_data_out(2236),
        VN2CN5_bit => VN_data_out(2237),
        VN2CN0_sign => VN_sign_out(2232),
        VN2CN1_sign => VN_sign_out(2233),
        VN2CN2_sign => VN_sign_out(2234),
        VN2CN3_sign => VN_sign_out(2235),
        VN2CN4_sign => VN_sign_out(2236),
        VN2CN5_sign => VN_sign_out(2237),
        codeword => codeword(372),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN373 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2243 downto 2238),
        Din0 => VN373_in0,
        Din1 => VN373_in1,
        Din2 => VN373_in2,
        Din3 => VN373_in3,
        Din4 => VN373_in4,
        Din5 => VN373_in5,
        VN2CN0_bit => VN_data_out(2238),
        VN2CN1_bit => VN_data_out(2239),
        VN2CN2_bit => VN_data_out(2240),
        VN2CN3_bit => VN_data_out(2241),
        VN2CN4_bit => VN_data_out(2242),
        VN2CN5_bit => VN_data_out(2243),
        VN2CN0_sign => VN_sign_out(2238),
        VN2CN1_sign => VN_sign_out(2239),
        VN2CN2_sign => VN_sign_out(2240),
        VN2CN3_sign => VN_sign_out(2241),
        VN2CN4_sign => VN_sign_out(2242),
        VN2CN5_sign => VN_sign_out(2243),
        codeword => codeword(373),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN374 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2249 downto 2244),
        Din0 => VN374_in0,
        Din1 => VN374_in1,
        Din2 => VN374_in2,
        Din3 => VN374_in3,
        Din4 => VN374_in4,
        Din5 => VN374_in5,
        VN2CN0_bit => VN_data_out(2244),
        VN2CN1_bit => VN_data_out(2245),
        VN2CN2_bit => VN_data_out(2246),
        VN2CN3_bit => VN_data_out(2247),
        VN2CN4_bit => VN_data_out(2248),
        VN2CN5_bit => VN_data_out(2249),
        VN2CN0_sign => VN_sign_out(2244),
        VN2CN1_sign => VN_sign_out(2245),
        VN2CN2_sign => VN_sign_out(2246),
        VN2CN3_sign => VN_sign_out(2247),
        VN2CN4_sign => VN_sign_out(2248),
        VN2CN5_sign => VN_sign_out(2249),
        codeword => codeword(374),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN375 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2255 downto 2250),
        Din0 => VN375_in0,
        Din1 => VN375_in1,
        Din2 => VN375_in2,
        Din3 => VN375_in3,
        Din4 => VN375_in4,
        Din5 => VN375_in5,
        VN2CN0_bit => VN_data_out(2250),
        VN2CN1_bit => VN_data_out(2251),
        VN2CN2_bit => VN_data_out(2252),
        VN2CN3_bit => VN_data_out(2253),
        VN2CN4_bit => VN_data_out(2254),
        VN2CN5_bit => VN_data_out(2255),
        VN2CN0_sign => VN_sign_out(2250),
        VN2CN1_sign => VN_sign_out(2251),
        VN2CN2_sign => VN_sign_out(2252),
        VN2CN3_sign => VN_sign_out(2253),
        VN2CN4_sign => VN_sign_out(2254),
        VN2CN5_sign => VN_sign_out(2255),
        codeword => codeword(375),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN376 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2261 downto 2256),
        Din0 => VN376_in0,
        Din1 => VN376_in1,
        Din2 => VN376_in2,
        Din3 => VN376_in3,
        Din4 => VN376_in4,
        Din5 => VN376_in5,
        VN2CN0_bit => VN_data_out(2256),
        VN2CN1_bit => VN_data_out(2257),
        VN2CN2_bit => VN_data_out(2258),
        VN2CN3_bit => VN_data_out(2259),
        VN2CN4_bit => VN_data_out(2260),
        VN2CN5_bit => VN_data_out(2261),
        VN2CN0_sign => VN_sign_out(2256),
        VN2CN1_sign => VN_sign_out(2257),
        VN2CN2_sign => VN_sign_out(2258),
        VN2CN3_sign => VN_sign_out(2259),
        VN2CN4_sign => VN_sign_out(2260),
        VN2CN5_sign => VN_sign_out(2261),
        codeword => codeword(376),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN377 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2267 downto 2262),
        Din0 => VN377_in0,
        Din1 => VN377_in1,
        Din2 => VN377_in2,
        Din3 => VN377_in3,
        Din4 => VN377_in4,
        Din5 => VN377_in5,
        VN2CN0_bit => VN_data_out(2262),
        VN2CN1_bit => VN_data_out(2263),
        VN2CN2_bit => VN_data_out(2264),
        VN2CN3_bit => VN_data_out(2265),
        VN2CN4_bit => VN_data_out(2266),
        VN2CN5_bit => VN_data_out(2267),
        VN2CN0_sign => VN_sign_out(2262),
        VN2CN1_sign => VN_sign_out(2263),
        VN2CN2_sign => VN_sign_out(2264),
        VN2CN3_sign => VN_sign_out(2265),
        VN2CN4_sign => VN_sign_out(2266),
        VN2CN5_sign => VN_sign_out(2267),
        codeword => codeword(377),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN378 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2273 downto 2268),
        Din0 => VN378_in0,
        Din1 => VN378_in1,
        Din2 => VN378_in2,
        Din3 => VN378_in3,
        Din4 => VN378_in4,
        Din5 => VN378_in5,
        VN2CN0_bit => VN_data_out(2268),
        VN2CN1_bit => VN_data_out(2269),
        VN2CN2_bit => VN_data_out(2270),
        VN2CN3_bit => VN_data_out(2271),
        VN2CN4_bit => VN_data_out(2272),
        VN2CN5_bit => VN_data_out(2273),
        VN2CN0_sign => VN_sign_out(2268),
        VN2CN1_sign => VN_sign_out(2269),
        VN2CN2_sign => VN_sign_out(2270),
        VN2CN3_sign => VN_sign_out(2271),
        VN2CN4_sign => VN_sign_out(2272),
        VN2CN5_sign => VN_sign_out(2273),
        codeword => codeword(378),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN379 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2279 downto 2274),
        Din0 => VN379_in0,
        Din1 => VN379_in1,
        Din2 => VN379_in2,
        Din3 => VN379_in3,
        Din4 => VN379_in4,
        Din5 => VN379_in5,
        VN2CN0_bit => VN_data_out(2274),
        VN2CN1_bit => VN_data_out(2275),
        VN2CN2_bit => VN_data_out(2276),
        VN2CN3_bit => VN_data_out(2277),
        VN2CN4_bit => VN_data_out(2278),
        VN2CN5_bit => VN_data_out(2279),
        VN2CN0_sign => VN_sign_out(2274),
        VN2CN1_sign => VN_sign_out(2275),
        VN2CN2_sign => VN_sign_out(2276),
        VN2CN3_sign => VN_sign_out(2277),
        VN2CN4_sign => VN_sign_out(2278),
        VN2CN5_sign => VN_sign_out(2279),
        codeword => codeword(379),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN380 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2285 downto 2280),
        Din0 => VN380_in0,
        Din1 => VN380_in1,
        Din2 => VN380_in2,
        Din3 => VN380_in3,
        Din4 => VN380_in4,
        Din5 => VN380_in5,
        VN2CN0_bit => VN_data_out(2280),
        VN2CN1_bit => VN_data_out(2281),
        VN2CN2_bit => VN_data_out(2282),
        VN2CN3_bit => VN_data_out(2283),
        VN2CN4_bit => VN_data_out(2284),
        VN2CN5_bit => VN_data_out(2285),
        VN2CN0_sign => VN_sign_out(2280),
        VN2CN1_sign => VN_sign_out(2281),
        VN2CN2_sign => VN_sign_out(2282),
        VN2CN3_sign => VN_sign_out(2283),
        VN2CN4_sign => VN_sign_out(2284),
        VN2CN5_sign => VN_sign_out(2285),
        codeword => codeword(380),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN381 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2291 downto 2286),
        Din0 => VN381_in0,
        Din1 => VN381_in1,
        Din2 => VN381_in2,
        Din3 => VN381_in3,
        Din4 => VN381_in4,
        Din5 => VN381_in5,
        VN2CN0_bit => VN_data_out(2286),
        VN2CN1_bit => VN_data_out(2287),
        VN2CN2_bit => VN_data_out(2288),
        VN2CN3_bit => VN_data_out(2289),
        VN2CN4_bit => VN_data_out(2290),
        VN2CN5_bit => VN_data_out(2291),
        VN2CN0_sign => VN_sign_out(2286),
        VN2CN1_sign => VN_sign_out(2287),
        VN2CN2_sign => VN_sign_out(2288),
        VN2CN3_sign => VN_sign_out(2289),
        VN2CN4_sign => VN_sign_out(2290),
        VN2CN5_sign => VN_sign_out(2291),
        codeword => codeword(381),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN382 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2297 downto 2292),
        Din0 => VN382_in0,
        Din1 => VN382_in1,
        Din2 => VN382_in2,
        Din3 => VN382_in3,
        Din4 => VN382_in4,
        Din5 => VN382_in5,
        VN2CN0_bit => VN_data_out(2292),
        VN2CN1_bit => VN_data_out(2293),
        VN2CN2_bit => VN_data_out(2294),
        VN2CN3_bit => VN_data_out(2295),
        VN2CN4_bit => VN_data_out(2296),
        VN2CN5_bit => VN_data_out(2297),
        VN2CN0_sign => VN_sign_out(2292),
        VN2CN1_sign => VN_sign_out(2293),
        VN2CN2_sign => VN_sign_out(2294),
        VN2CN3_sign => VN_sign_out(2295),
        VN2CN4_sign => VN_sign_out(2296),
        VN2CN5_sign => VN_sign_out(2297),
        codeword => codeword(382),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN383 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2303 downto 2298),
        Din0 => VN383_in0,
        Din1 => VN383_in1,
        Din2 => VN383_in2,
        Din3 => VN383_in3,
        Din4 => VN383_in4,
        Din5 => VN383_in5,
        VN2CN0_bit => VN_data_out(2298),
        VN2CN1_bit => VN_data_out(2299),
        VN2CN2_bit => VN_data_out(2300),
        VN2CN3_bit => VN_data_out(2301),
        VN2CN4_bit => VN_data_out(2302),
        VN2CN5_bit => VN_data_out(2303),
        VN2CN0_sign => VN_sign_out(2298),
        VN2CN1_sign => VN_sign_out(2299),
        VN2CN2_sign => VN_sign_out(2300),
        VN2CN3_sign => VN_sign_out(2301),
        VN2CN4_sign => VN_sign_out(2302),
        VN2CN5_sign => VN_sign_out(2303),
        codeword => codeword(383),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN384 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2309 downto 2304),
        Din0 => VN384_in0,
        Din1 => VN384_in1,
        Din2 => VN384_in2,
        Din3 => VN384_in3,
        Din4 => VN384_in4,
        Din5 => VN384_in5,
        VN2CN0_bit => VN_data_out(2304),
        VN2CN1_bit => VN_data_out(2305),
        VN2CN2_bit => VN_data_out(2306),
        VN2CN3_bit => VN_data_out(2307),
        VN2CN4_bit => VN_data_out(2308),
        VN2CN5_bit => VN_data_out(2309),
        VN2CN0_sign => VN_sign_out(2304),
        VN2CN1_sign => VN_sign_out(2305),
        VN2CN2_sign => VN_sign_out(2306),
        VN2CN3_sign => VN_sign_out(2307),
        VN2CN4_sign => VN_sign_out(2308),
        VN2CN5_sign => VN_sign_out(2309),
        codeword => codeword(384),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN385 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2315 downto 2310),
        Din0 => VN385_in0,
        Din1 => VN385_in1,
        Din2 => VN385_in2,
        Din3 => VN385_in3,
        Din4 => VN385_in4,
        Din5 => VN385_in5,
        VN2CN0_bit => VN_data_out(2310),
        VN2CN1_bit => VN_data_out(2311),
        VN2CN2_bit => VN_data_out(2312),
        VN2CN3_bit => VN_data_out(2313),
        VN2CN4_bit => VN_data_out(2314),
        VN2CN5_bit => VN_data_out(2315),
        VN2CN0_sign => VN_sign_out(2310),
        VN2CN1_sign => VN_sign_out(2311),
        VN2CN2_sign => VN_sign_out(2312),
        VN2CN3_sign => VN_sign_out(2313),
        VN2CN4_sign => VN_sign_out(2314),
        VN2CN5_sign => VN_sign_out(2315),
        codeword => codeword(385),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN386 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2321 downto 2316),
        Din0 => VN386_in0,
        Din1 => VN386_in1,
        Din2 => VN386_in2,
        Din3 => VN386_in3,
        Din4 => VN386_in4,
        Din5 => VN386_in5,
        VN2CN0_bit => VN_data_out(2316),
        VN2CN1_bit => VN_data_out(2317),
        VN2CN2_bit => VN_data_out(2318),
        VN2CN3_bit => VN_data_out(2319),
        VN2CN4_bit => VN_data_out(2320),
        VN2CN5_bit => VN_data_out(2321),
        VN2CN0_sign => VN_sign_out(2316),
        VN2CN1_sign => VN_sign_out(2317),
        VN2CN2_sign => VN_sign_out(2318),
        VN2CN3_sign => VN_sign_out(2319),
        VN2CN4_sign => VN_sign_out(2320),
        VN2CN5_sign => VN_sign_out(2321),
        codeword => codeword(386),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN387 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2327 downto 2322),
        Din0 => VN387_in0,
        Din1 => VN387_in1,
        Din2 => VN387_in2,
        Din3 => VN387_in3,
        Din4 => VN387_in4,
        Din5 => VN387_in5,
        VN2CN0_bit => VN_data_out(2322),
        VN2CN1_bit => VN_data_out(2323),
        VN2CN2_bit => VN_data_out(2324),
        VN2CN3_bit => VN_data_out(2325),
        VN2CN4_bit => VN_data_out(2326),
        VN2CN5_bit => VN_data_out(2327),
        VN2CN0_sign => VN_sign_out(2322),
        VN2CN1_sign => VN_sign_out(2323),
        VN2CN2_sign => VN_sign_out(2324),
        VN2CN3_sign => VN_sign_out(2325),
        VN2CN4_sign => VN_sign_out(2326),
        VN2CN5_sign => VN_sign_out(2327),
        codeword => codeword(387),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN388 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2333 downto 2328),
        Din0 => VN388_in0,
        Din1 => VN388_in1,
        Din2 => VN388_in2,
        Din3 => VN388_in3,
        Din4 => VN388_in4,
        Din5 => VN388_in5,
        VN2CN0_bit => VN_data_out(2328),
        VN2CN1_bit => VN_data_out(2329),
        VN2CN2_bit => VN_data_out(2330),
        VN2CN3_bit => VN_data_out(2331),
        VN2CN4_bit => VN_data_out(2332),
        VN2CN5_bit => VN_data_out(2333),
        VN2CN0_sign => VN_sign_out(2328),
        VN2CN1_sign => VN_sign_out(2329),
        VN2CN2_sign => VN_sign_out(2330),
        VN2CN3_sign => VN_sign_out(2331),
        VN2CN4_sign => VN_sign_out(2332),
        VN2CN5_sign => VN_sign_out(2333),
        codeword => codeword(388),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN389 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2339 downto 2334),
        Din0 => VN389_in0,
        Din1 => VN389_in1,
        Din2 => VN389_in2,
        Din3 => VN389_in3,
        Din4 => VN389_in4,
        Din5 => VN389_in5,
        VN2CN0_bit => VN_data_out(2334),
        VN2CN1_bit => VN_data_out(2335),
        VN2CN2_bit => VN_data_out(2336),
        VN2CN3_bit => VN_data_out(2337),
        VN2CN4_bit => VN_data_out(2338),
        VN2CN5_bit => VN_data_out(2339),
        VN2CN0_sign => VN_sign_out(2334),
        VN2CN1_sign => VN_sign_out(2335),
        VN2CN2_sign => VN_sign_out(2336),
        VN2CN3_sign => VN_sign_out(2337),
        VN2CN4_sign => VN_sign_out(2338),
        VN2CN5_sign => VN_sign_out(2339),
        codeword => codeword(389),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN390 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2345 downto 2340),
        Din0 => VN390_in0,
        Din1 => VN390_in1,
        Din2 => VN390_in2,
        Din3 => VN390_in3,
        Din4 => VN390_in4,
        Din5 => VN390_in5,
        VN2CN0_bit => VN_data_out(2340),
        VN2CN1_bit => VN_data_out(2341),
        VN2CN2_bit => VN_data_out(2342),
        VN2CN3_bit => VN_data_out(2343),
        VN2CN4_bit => VN_data_out(2344),
        VN2CN5_bit => VN_data_out(2345),
        VN2CN0_sign => VN_sign_out(2340),
        VN2CN1_sign => VN_sign_out(2341),
        VN2CN2_sign => VN_sign_out(2342),
        VN2CN3_sign => VN_sign_out(2343),
        VN2CN4_sign => VN_sign_out(2344),
        VN2CN5_sign => VN_sign_out(2345),
        codeword => codeword(390),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN391 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2351 downto 2346),
        Din0 => VN391_in0,
        Din1 => VN391_in1,
        Din2 => VN391_in2,
        Din3 => VN391_in3,
        Din4 => VN391_in4,
        Din5 => VN391_in5,
        VN2CN0_bit => VN_data_out(2346),
        VN2CN1_bit => VN_data_out(2347),
        VN2CN2_bit => VN_data_out(2348),
        VN2CN3_bit => VN_data_out(2349),
        VN2CN4_bit => VN_data_out(2350),
        VN2CN5_bit => VN_data_out(2351),
        VN2CN0_sign => VN_sign_out(2346),
        VN2CN1_sign => VN_sign_out(2347),
        VN2CN2_sign => VN_sign_out(2348),
        VN2CN3_sign => VN_sign_out(2349),
        VN2CN4_sign => VN_sign_out(2350),
        VN2CN5_sign => VN_sign_out(2351),
        codeword => codeword(391),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN392 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2357 downto 2352),
        Din0 => VN392_in0,
        Din1 => VN392_in1,
        Din2 => VN392_in2,
        Din3 => VN392_in3,
        Din4 => VN392_in4,
        Din5 => VN392_in5,
        VN2CN0_bit => VN_data_out(2352),
        VN2CN1_bit => VN_data_out(2353),
        VN2CN2_bit => VN_data_out(2354),
        VN2CN3_bit => VN_data_out(2355),
        VN2CN4_bit => VN_data_out(2356),
        VN2CN5_bit => VN_data_out(2357),
        VN2CN0_sign => VN_sign_out(2352),
        VN2CN1_sign => VN_sign_out(2353),
        VN2CN2_sign => VN_sign_out(2354),
        VN2CN3_sign => VN_sign_out(2355),
        VN2CN4_sign => VN_sign_out(2356),
        VN2CN5_sign => VN_sign_out(2357),
        codeword => codeword(392),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN393 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2363 downto 2358),
        Din0 => VN393_in0,
        Din1 => VN393_in1,
        Din2 => VN393_in2,
        Din3 => VN393_in3,
        Din4 => VN393_in4,
        Din5 => VN393_in5,
        VN2CN0_bit => VN_data_out(2358),
        VN2CN1_bit => VN_data_out(2359),
        VN2CN2_bit => VN_data_out(2360),
        VN2CN3_bit => VN_data_out(2361),
        VN2CN4_bit => VN_data_out(2362),
        VN2CN5_bit => VN_data_out(2363),
        VN2CN0_sign => VN_sign_out(2358),
        VN2CN1_sign => VN_sign_out(2359),
        VN2CN2_sign => VN_sign_out(2360),
        VN2CN3_sign => VN_sign_out(2361),
        VN2CN4_sign => VN_sign_out(2362),
        VN2CN5_sign => VN_sign_out(2363),
        codeword => codeword(393),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN394 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2369 downto 2364),
        Din0 => VN394_in0,
        Din1 => VN394_in1,
        Din2 => VN394_in2,
        Din3 => VN394_in3,
        Din4 => VN394_in4,
        Din5 => VN394_in5,
        VN2CN0_bit => VN_data_out(2364),
        VN2CN1_bit => VN_data_out(2365),
        VN2CN2_bit => VN_data_out(2366),
        VN2CN3_bit => VN_data_out(2367),
        VN2CN4_bit => VN_data_out(2368),
        VN2CN5_bit => VN_data_out(2369),
        VN2CN0_sign => VN_sign_out(2364),
        VN2CN1_sign => VN_sign_out(2365),
        VN2CN2_sign => VN_sign_out(2366),
        VN2CN3_sign => VN_sign_out(2367),
        VN2CN4_sign => VN_sign_out(2368),
        VN2CN5_sign => VN_sign_out(2369),
        codeword => codeword(394),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN395 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2375 downto 2370),
        Din0 => VN395_in0,
        Din1 => VN395_in1,
        Din2 => VN395_in2,
        Din3 => VN395_in3,
        Din4 => VN395_in4,
        Din5 => VN395_in5,
        VN2CN0_bit => VN_data_out(2370),
        VN2CN1_bit => VN_data_out(2371),
        VN2CN2_bit => VN_data_out(2372),
        VN2CN3_bit => VN_data_out(2373),
        VN2CN4_bit => VN_data_out(2374),
        VN2CN5_bit => VN_data_out(2375),
        VN2CN0_sign => VN_sign_out(2370),
        VN2CN1_sign => VN_sign_out(2371),
        VN2CN2_sign => VN_sign_out(2372),
        VN2CN3_sign => VN_sign_out(2373),
        VN2CN4_sign => VN_sign_out(2374),
        VN2CN5_sign => VN_sign_out(2375),
        codeword => codeword(395),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN396 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2381 downto 2376),
        Din0 => VN396_in0,
        Din1 => VN396_in1,
        Din2 => VN396_in2,
        Din3 => VN396_in3,
        Din4 => VN396_in4,
        Din5 => VN396_in5,
        VN2CN0_bit => VN_data_out(2376),
        VN2CN1_bit => VN_data_out(2377),
        VN2CN2_bit => VN_data_out(2378),
        VN2CN3_bit => VN_data_out(2379),
        VN2CN4_bit => VN_data_out(2380),
        VN2CN5_bit => VN_data_out(2381),
        VN2CN0_sign => VN_sign_out(2376),
        VN2CN1_sign => VN_sign_out(2377),
        VN2CN2_sign => VN_sign_out(2378),
        VN2CN3_sign => VN_sign_out(2379),
        VN2CN4_sign => VN_sign_out(2380),
        VN2CN5_sign => VN_sign_out(2381),
        codeword => codeword(396),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN397 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2387 downto 2382),
        Din0 => VN397_in0,
        Din1 => VN397_in1,
        Din2 => VN397_in2,
        Din3 => VN397_in3,
        Din4 => VN397_in4,
        Din5 => VN397_in5,
        VN2CN0_bit => VN_data_out(2382),
        VN2CN1_bit => VN_data_out(2383),
        VN2CN2_bit => VN_data_out(2384),
        VN2CN3_bit => VN_data_out(2385),
        VN2CN4_bit => VN_data_out(2386),
        VN2CN5_bit => VN_data_out(2387),
        VN2CN0_sign => VN_sign_out(2382),
        VN2CN1_sign => VN_sign_out(2383),
        VN2CN2_sign => VN_sign_out(2384),
        VN2CN3_sign => VN_sign_out(2385),
        VN2CN4_sign => VN_sign_out(2386),
        VN2CN5_sign => VN_sign_out(2387),
        codeword => codeword(397),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN398 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2393 downto 2388),
        Din0 => VN398_in0,
        Din1 => VN398_in1,
        Din2 => VN398_in2,
        Din3 => VN398_in3,
        Din4 => VN398_in4,
        Din5 => VN398_in5,
        VN2CN0_bit => VN_data_out(2388),
        VN2CN1_bit => VN_data_out(2389),
        VN2CN2_bit => VN_data_out(2390),
        VN2CN3_bit => VN_data_out(2391),
        VN2CN4_bit => VN_data_out(2392),
        VN2CN5_bit => VN_data_out(2393),
        VN2CN0_sign => VN_sign_out(2388),
        VN2CN1_sign => VN_sign_out(2389),
        VN2CN2_sign => VN_sign_out(2390),
        VN2CN3_sign => VN_sign_out(2391),
        VN2CN4_sign => VN_sign_out(2392),
        VN2CN5_sign => VN_sign_out(2393),
        codeword => codeword(398),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN399 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2399 downto 2394),
        Din0 => VN399_in0,
        Din1 => VN399_in1,
        Din2 => VN399_in2,
        Din3 => VN399_in3,
        Din4 => VN399_in4,
        Din5 => VN399_in5,
        VN2CN0_bit => VN_data_out(2394),
        VN2CN1_bit => VN_data_out(2395),
        VN2CN2_bit => VN_data_out(2396),
        VN2CN3_bit => VN_data_out(2397),
        VN2CN4_bit => VN_data_out(2398),
        VN2CN5_bit => VN_data_out(2399),
        VN2CN0_sign => VN_sign_out(2394),
        VN2CN1_sign => VN_sign_out(2395),
        VN2CN2_sign => VN_sign_out(2396),
        VN2CN3_sign => VN_sign_out(2397),
        VN2CN4_sign => VN_sign_out(2398),
        VN2CN5_sign => VN_sign_out(2399),
        codeword => codeword(399),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN400 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2405 downto 2400),
        Din0 => VN400_in0,
        Din1 => VN400_in1,
        Din2 => VN400_in2,
        Din3 => VN400_in3,
        Din4 => VN400_in4,
        Din5 => VN400_in5,
        VN2CN0_bit => VN_data_out(2400),
        VN2CN1_bit => VN_data_out(2401),
        VN2CN2_bit => VN_data_out(2402),
        VN2CN3_bit => VN_data_out(2403),
        VN2CN4_bit => VN_data_out(2404),
        VN2CN5_bit => VN_data_out(2405),
        VN2CN0_sign => VN_sign_out(2400),
        VN2CN1_sign => VN_sign_out(2401),
        VN2CN2_sign => VN_sign_out(2402),
        VN2CN3_sign => VN_sign_out(2403),
        VN2CN4_sign => VN_sign_out(2404),
        VN2CN5_sign => VN_sign_out(2405),
        codeword => codeword(400),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN401 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2411 downto 2406),
        Din0 => VN401_in0,
        Din1 => VN401_in1,
        Din2 => VN401_in2,
        Din3 => VN401_in3,
        Din4 => VN401_in4,
        Din5 => VN401_in5,
        VN2CN0_bit => VN_data_out(2406),
        VN2CN1_bit => VN_data_out(2407),
        VN2CN2_bit => VN_data_out(2408),
        VN2CN3_bit => VN_data_out(2409),
        VN2CN4_bit => VN_data_out(2410),
        VN2CN5_bit => VN_data_out(2411),
        VN2CN0_sign => VN_sign_out(2406),
        VN2CN1_sign => VN_sign_out(2407),
        VN2CN2_sign => VN_sign_out(2408),
        VN2CN3_sign => VN_sign_out(2409),
        VN2CN4_sign => VN_sign_out(2410),
        VN2CN5_sign => VN_sign_out(2411),
        codeword => codeword(401),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN402 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2417 downto 2412),
        Din0 => VN402_in0,
        Din1 => VN402_in1,
        Din2 => VN402_in2,
        Din3 => VN402_in3,
        Din4 => VN402_in4,
        Din5 => VN402_in5,
        VN2CN0_bit => VN_data_out(2412),
        VN2CN1_bit => VN_data_out(2413),
        VN2CN2_bit => VN_data_out(2414),
        VN2CN3_bit => VN_data_out(2415),
        VN2CN4_bit => VN_data_out(2416),
        VN2CN5_bit => VN_data_out(2417),
        VN2CN0_sign => VN_sign_out(2412),
        VN2CN1_sign => VN_sign_out(2413),
        VN2CN2_sign => VN_sign_out(2414),
        VN2CN3_sign => VN_sign_out(2415),
        VN2CN4_sign => VN_sign_out(2416),
        VN2CN5_sign => VN_sign_out(2417),
        codeword => codeword(402),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN403 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2423 downto 2418),
        Din0 => VN403_in0,
        Din1 => VN403_in1,
        Din2 => VN403_in2,
        Din3 => VN403_in3,
        Din4 => VN403_in4,
        Din5 => VN403_in5,
        VN2CN0_bit => VN_data_out(2418),
        VN2CN1_bit => VN_data_out(2419),
        VN2CN2_bit => VN_data_out(2420),
        VN2CN3_bit => VN_data_out(2421),
        VN2CN4_bit => VN_data_out(2422),
        VN2CN5_bit => VN_data_out(2423),
        VN2CN0_sign => VN_sign_out(2418),
        VN2CN1_sign => VN_sign_out(2419),
        VN2CN2_sign => VN_sign_out(2420),
        VN2CN3_sign => VN_sign_out(2421),
        VN2CN4_sign => VN_sign_out(2422),
        VN2CN5_sign => VN_sign_out(2423),
        codeword => codeword(403),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN404 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2429 downto 2424),
        Din0 => VN404_in0,
        Din1 => VN404_in1,
        Din2 => VN404_in2,
        Din3 => VN404_in3,
        Din4 => VN404_in4,
        Din5 => VN404_in5,
        VN2CN0_bit => VN_data_out(2424),
        VN2CN1_bit => VN_data_out(2425),
        VN2CN2_bit => VN_data_out(2426),
        VN2CN3_bit => VN_data_out(2427),
        VN2CN4_bit => VN_data_out(2428),
        VN2CN5_bit => VN_data_out(2429),
        VN2CN0_sign => VN_sign_out(2424),
        VN2CN1_sign => VN_sign_out(2425),
        VN2CN2_sign => VN_sign_out(2426),
        VN2CN3_sign => VN_sign_out(2427),
        VN2CN4_sign => VN_sign_out(2428),
        VN2CN5_sign => VN_sign_out(2429),
        codeword => codeword(404),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN405 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2435 downto 2430),
        Din0 => VN405_in0,
        Din1 => VN405_in1,
        Din2 => VN405_in2,
        Din3 => VN405_in3,
        Din4 => VN405_in4,
        Din5 => VN405_in5,
        VN2CN0_bit => VN_data_out(2430),
        VN2CN1_bit => VN_data_out(2431),
        VN2CN2_bit => VN_data_out(2432),
        VN2CN3_bit => VN_data_out(2433),
        VN2CN4_bit => VN_data_out(2434),
        VN2CN5_bit => VN_data_out(2435),
        VN2CN0_sign => VN_sign_out(2430),
        VN2CN1_sign => VN_sign_out(2431),
        VN2CN2_sign => VN_sign_out(2432),
        VN2CN3_sign => VN_sign_out(2433),
        VN2CN4_sign => VN_sign_out(2434),
        VN2CN5_sign => VN_sign_out(2435),
        codeword => codeword(405),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN406 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2441 downto 2436),
        Din0 => VN406_in0,
        Din1 => VN406_in1,
        Din2 => VN406_in2,
        Din3 => VN406_in3,
        Din4 => VN406_in4,
        Din5 => VN406_in5,
        VN2CN0_bit => VN_data_out(2436),
        VN2CN1_bit => VN_data_out(2437),
        VN2CN2_bit => VN_data_out(2438),
        VN2CN3_bit => VN_data_out(2439),
        VN2CN4_bit => VN_data_out(2440),
        VN2CN5_bit => VN_data_out(2441),
        VN2CN0_sign => VN_sign_out(2436),
        VN2CN1_sign => VN_sign_out(2437),
        VN2CN2_sign => VN_sign_out(2438),
        VN2CN3_sign => VN_sign_out(2439),
        VN2CN4_sign => VN_sign_out(2440),
        VN2CN5_sign => VN_sign_out(2441),
        codeword => codeword(406),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN407 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2447 downto 2442),
        Din0 => VN407_in0,
        Din1 => VN407_in1,
        Din2 => VN407_in2,
        Din3 => VN407_in3,
        Din4 => VN407_in4,
        Din5 => VN407_in5,
        VN2CN0_bit => VN_data_out(2442),
        VN2CN1_bit => VN_data_out(2443),
        VN2CN2_bit => VN_data_out(2444),
        VN2CN3_bit => VN_data_out(2445),
        VN2CN4_bit => VN_data_out(2446),
        VN2CN5_bit => VN_data_out(2447),
        VN2CN0_sign => VN_sign_out(2442),
        VN2CN1_sign => VN_sign_out(2443),
        VN2CN2_sign => VN_sign_out(2444),
        VN2CN3_sign => VN_sign_out(2445),
        VN2CN4_sign => VN_sign_out(2446),
        VN2CN5_sign => VN_sign_out(2447),
        codeword => codeword(407),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN408 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2453 downto 2448),
        Din0 => VN408_in0,
        Din1 => VN408_in1,
        Din2 => VN408_in2,
        Din3 => VN408_in3,
        Din4 => VN408_in4,
        Din5 => VN408_in5,
        VN2CN0_bit => VN_data_out(2448),
        VN2CN1_bit => VN_data_out(2449),
        VN2CN2_bit => VN_data_out(2450),
        VN2CN3_bit => VN_data_out(2451),
        VN2CN4_bit => VN_data_out(2452),
        VN2CN5_bit => VN_data_out(2453),
        VN2CN0_sign => VN_sign_out(2448),
        VN2CN1_sign => VN_sign_out(2449),
        VN2CN2_sign => VN_sign_out(2450),
        VN2CN3_sign => VN_sign_out(2451),
        VN2CN4_sign => VN_sign_out(2452),
        VN2CN5_sign => VN_sign_out(2453),
        codeword => codeword(408),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN409 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2459 downto 2454),
        Din0 => VN409_in0,
        Din1 => VN409_in1,
        Din2 => VN409_in2,
        Din3 => VN409_in3,
        Din4 => VN409_in4,
        Din5 => VN409_in5,
        VN2CN0_bit => VN_data_out(2454),
        VN2CN1_bit => VN_data_out(2455),
        VN2CN2_bit => VN_data_out(2456),
        VN2CN3_bit => VN_data_out(2457),
        VN2CN4_bit => VN_data_out(2458),
        VN2CN5_bit => VN_data_out(2459),
        VN2CN0_sign => VN_sign_out(2454),
        VN2CN1_sign => VN_sign_out(2455),
        VN2CN2_sign => VN_sign_out(2456),
        VN2CN3_sign => VN_sign_out(2457),
        VN2CN4_sign => VN_sign_out(2458),
        VN2CN5_sign => VN_sign_out(2459),
        codeword => codeword(409),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN410 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2465 downto 2460),
        Din0 => VN410_in0,
        Din1 => VN410_in1,
        Din2 => VN410_in2,
        Din3 => VN410_in3,
        Din4 => VN410_in4,
        Din5 => VN410_in5,
        VN2CN0_bit => VN_data_out(2460),
        VN2CN1_bit => VN_data_out(2461),
        VN2CN2_bit => VN_data_out(2462),
        VN2CN3_bit => VN_data_out(2463),
        VN2CN4_bit => VN_data_out(2464),
        VN2CN5_bit => VN_data_out(2465),
        VN2CN0_sign => VN_sign_out(2460),
        VN2CN1_sign => VN_sign_out(2461),
        VN2CN2_sign => VN_sign_out(2462),
        VN2CN3_sign => VN_sign_out(2463),
        VN2CN4_sign => VN_sign_out(2464),
        VN2CN5_sign => VN_sign_out(2465),
        codeword => codeword(410),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN411 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2471 downto 2466),
        Din0 => VN411_in0,
        Din1 => VN411_in1,
        Din2 => VN411_in2,
        Din3 => VN411_in3,
        Din4 => VN411_in4,
        Din5 => VN411_in5,
        VN2CN0_bit => VN_data_out(2466),
        VN2CN1_bit => VN_data_out(2467),
        VN2CN2_bit => VN_data_out(2468),
        VN2CN3_bit => VN_data_out(2469),
        VN2CN4_bit => VN_data_out(2470),
        VN2CN5_bit => VN_data_out(2471),
        VN2CN0_sign => VN_sign_out(2466),
        VN2CN1_sign => VN_sign_out(2467),
        VN2CN2_sign => VN_sign_out(2468),
        VN2CN3_sign => VN_sign_out(2469),
        VN2CN4_sign => VN_sign_out(2470),
        VN2CN5_sign => VN_sign_out(2471),
        codeword => codeword(411),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN412 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2477 downto 2472),
        Din0 => VN412_in0,
        Din1 => VN412_in1,
        Din2 => VN412_in2,
        Din3 => VN412_in3,
        Din4 => VN412_in4,
        Din5 => VN412_in5,
        VN2CN0_bit => VN_data_out(2472),
        VN2CN1_bit => VN_data_out(2473),
        VN2CN2_bit => VN_data_out(2474),
        VN2CN3_bit => VN_data_out(2475),
        VN2CN4_bit => VN_data_out(2476),
        VN2CN5_bit => VN_data_out(2477),
        VN2CN0_sign => VN_sign_out(2472),
        VN2CN1_sign => VN_sign_out(2473),
        VN2CN2_sign => VN_sign_out(2474),
        VN2CN3_sign => VN_sign_out(2475),
        VN2CN4_sign => VN_sign_out(2476),
        VN2CN5_sign => VN_sign_out(2477),
        codeword => codeword(412),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN413 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2483 downto 2478),
        Din0 => VN413_in0,
        Din1 => VN413_in1,
        Din2 => VN413_in2,
        Din3 => VN413_in3,
        Din4 => VN413_in4,
        Din5 => VN413_in5,
        VN2CN0_bit => VN_data_out(2478),
        VN2CN1_bit => VN_data_out(2479),
        VN2CN2_bit => VN_data_out(2480),
        VN2CN3_bit => VN_data_out(2481),
        VN2CN4_bit => VN_data_out(2482),
        VN2CN5_bit => VN_data_out(2483),
        VN2CN0_sign => VN_sign_out(2478),
        VN2CN1_sign => VN_sign_out(2479),
        VN2CN2_sign => VN_sign_out(2480),
        VN2CN3_sign => VN_sign_out(2481),
        VN2CN4_sign => VN_sign_out(2482),
        VN2CN5_sign => VN_sign_out(2483),
        codeword => codeword(413),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN414 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2489 downto 2484),
        Din0 => VN414_in0,
        Din1 => VN414_in1,
        Din2 => VN414_in2,
        Din3 => VN414_in3,
        Din4 => VN414_in4,
        Din5 => VN414_in5,
        VN2CN0_bit => VN_data_out(2484),
        VN2CN1_bit => VN_data_out(2485),
        VN2CN2_bit => VN_data_out(2486),
        VN2CN3_bit => VN_data_out(2487),
        VN2CN4_bit => VN_data_out(2488),
        VN2CN5_bit => VN_data_out(2489),
        VN2CN0_sign => VN_sign_out(2484),
        VN2CN1_sign => VN_sign_out(2485),
        VN2CN2_sign => VN_sign_out(2486),
        VN2CN3_sign => VN_sign_out(2487),
        VN2CN4_sign => VN_sign_out(2488),
        VN2CN5_sign => VN_sign_out(2489),
        codeword => codeword(414),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN415 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2495 downto 2490),
        Din0 => VN415_in0,
        Din1 => VN415_in1,
        Din2 => VN415_in2,
        Din3 => VN415_in3,
        Din4 => VN415_in4,
        Din5 => VN415_in5,
        VN2CN0_bit => VN_data_out(2490),
        VN2CN1_bit => VN_data_out(2491),
        VN2CN2_bit => VN_data_out(2492),
        VN2CN3_bit => VN_data_out(2493),
        VN2CN4_bit => VN_data_out(2494),
        VN2CN5_bit => VN_data_out(2495),
        VN2CN0_sign => VN_sign_out(2490),
        VN2CN1_sign => VN_sign_out(2491),
        VN2CN2_sign => VN_sign_out(2492),
        VN2CN3_sign => VN_sign_out(2493),
        VN2CN4_sign => VN_sign_out(2494),
        VN2CN5_sign => VN_sign_out(2495),
        codeword => codeword(415),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN416 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2501 downto 2496),
        Din0 => VN416_in0,
        Din1 => VN416_in1,
        Din2 => VN416_in2,
        Din3 => VN416_in3,
        Din4 => VN416_in4,
        Din5 => VN416_in5,
        VN2CN0_bit => VN_data_out(2496),
        VN2CN1_bit => VN_data_out(2497),
        VN2CN2_bit => VN_data_out(2498),
        VN2CN3_bit => VN_data_out(2499),
        VN2CN4_bit => VN_data_out(2500),
        VN2CN5_bit => VN_data_out(2501),
        VN2CN0_sign => VN_sign_out(2496),
        VN2CN1_sign => VN_sign_out(2497),
        VN2CN2_sign => VN_sign_out(2498),
        VN2CN3_sign => VN_sign_out(2499),
        VN2CN4_sign => VN_sign_out(2500),
        VN2CN5_sign => VN_sign_out(2501),
        codeword => codeword(416),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN417 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2507 downto 2502),
        Din0 => VN417_in0,
        Din1 => VN417_in1,
        Din2 => VN417_in2,
        Din3 => VN417_in3,
        Din4 => VN417_in4,
        Din5 => VN417_in5,
        VN2CN0_bit => VN_data_out(2502),
        VN2CN1_bit => VN_data_out(2503),
        VN2CN2_bit => VN_data_out(2504),
        VN2CN3_bit => VN_data_out(2505),
        VN2CN4_bit => VN_data_out(2506),
        VN2CN5_bit => VN_data_out(2507),
        VN2CN0_sign => VN_sign_out(2502),
        VN2CN1_sign => VN_sign_out(2503),
        VN2CN2_sign => VN_sign_out(2504),
        VN2CN3_sign => VN_sign_out(2505),
        VN2CN4_sign => VN_sign_out(2506),
        VN2CN5_sign => VN_sign_out(2507),
        codeword => codeword(417),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN418 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2513 downto 2508),
        Din0 => VN418_in0,
        Din1 => VN418_in1,
        Din2 => VN418_in2,
        Din3 => VN418_in3,
        Din4 => VN418_in4,
        Din5 => VN418_in5,
        VN2CN0_bit => VN_data_out(2508),
        VN2CN1_bit => VN_data_out(2509),
        VN2CN2_bit => VN_data_out(2510),
        VN2CN3_bit => VN_data_out(2511),
        VN2CN4_bit => VN_data_out(2512),
        VN2CN5_bit => VN_data_out(2513),
        VN2CN0_sign => VN_sign_out(2508),
        VN2CN1_sign => VN_sign_out(2509),
        VN2CN2_sign => VN_sign_out(2510),
        VN2CN3_sign => VN_sign_out(2511),
        VN2CN4_sign => VN_sign_out(2512),
        VN2CN5_sign => VN_sign_out(2513),
        codeword => codeword(418),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN419 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2519 downto 2514),
        Din0 => VN419_in0,
        Din1 => VN419_in1,
        Din2 => VN419_in2,
        Din3 => VN419_in3,
        Din4 => VN419_in4,
        Din5 => VN419_in5,
        VN2CN0_bit => VN_data_out(2514),
        VN2CN1_bit => VN_data_out(2515),
        VN2CN2_bit => VN_data_out(2516),
        VN2CN3_bit => VN_data_out(2517),
        VN2CN4_bit => VN_data_out(2518),
        VN2CN5_bit => VN_data_out(2519),
        VN2CN0_sign => VN_sign_out(2514),
        VN2CN1_sign => VN_sign_out(2515),
        VN2CN2_sign => VN_sign_out(2516),
        VN2CN3_sign => VN_sign_out(2517),
        VN2CN4_sign => VN_sign_out(2518),
        VN2CN5_sign => VN_sign_out(2519),
        codeword => codeword(419),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN420 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2525 downto 2520),
        Din0 => VN420_in0,
        Din1 => VN420_in1,
        Din2 => VN420_in2,
        Din3 => VN420_in3,
        Din4 => VN420_in4,
        Din5 => VN420_in5,
        VN2CN0_bit => VN_data_out(2520),
        VN2CN1_bit => VN_data_out(2521),
        VN2CN2_bit => VN_data_out(2522),
        VN2CN3_bit => VN_data_out(2523),
        VN2CN4_bit => VN_data_out(2524),
        VN2CN5_bit => VN_data_out(2525),
        VN2CN0_sign => VN_sign_out(2520),
        VN2CN1_sign => VN_sign_out(2521),
        VN2CN2_sign => VN_sign_out(2522),
        VN2CN3_sign => VN_sign_out(2523),
        VN2CN4_sign => VN_sign_out(2524),
        VN2CN5_sign => VN_sign_out(2525),
        codeword => codeword(420),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN421 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2531 downto 2526),
        Din0 => VN421_in0,
        Din1 => VN421_in1,
        Din2 => VN421_in2,
        Din3 => VN421_in3,
        Din4 => VN421_in4,
        Din5 => VN421_in5,
        VN2CN0_bit => VN_data_out(2526),
        VN2CN1_bit => VN_data_out(2527),
        VN2CN2_bit => VN_data_out(2528),
        VN2CN3_bit => VN_data_out(2529),
        VN2CN4_bit => VN_data_out(2530),
        VN2CN5_bit => VN_data_out(2531),
        VN2CN0_sign => VN_sign_out(2526),
        VN2CN1_sign => VN_sign_out(2527),
        VN2CN2_sign => VN_sign_out(2528),
        VN2CN3_sign => VN_sign_out(2529),
        VN2CN4_sign => VN_sign_out(2530),
        VN2CN5_sign => VN_sign_out(2531),
        codeword => codeword(421),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN422 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2537 downto 2532),
        Din0 => VN422_in0,
        Din1 => VN422_in1,
        Din2 => VN422_in2,
        Din3 => VN422_in3,
        Din4 => VN422_in4,
        Din5 => VN422_in5,
        VN2CN0_bit => VN_data_out(2532),
        VN2CN1_bit => VN_data_out(2533),
        VN2CN2_bit => VN_data_out(2534),
        VN2CN3_bit => VN_data_out(2535),
        VN2CN4_bit => VN_data_out(2536),
        VN2CN5_bit => VN_data_out(2537),
        VN2CN0_sign => VN_sign_out(2532),
        VN2CN1_sign => VN_sign_out(2533),
        VN2CN2_sign => VN_sign_out(2534),
        VN2CN3_sign => VN_sign_out(2535),
        VN2CN4_sign => VN_sign_out(2536),
        VN2CN5_sign => VN_sign_out(2537),
        codeword => codeword(422),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN423 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2543 downto 2538),
        Din0 => VN423_in0,
        Din1 => VN423_in1,
        Din2 => VN423_in2,
        Din3 => VN423_in3,
        Din4 => VN423_in4,
        Din5 => VN423_in5,
        VN2CN0_bit => VN_data_out(2538),
        VN2CN1_bit => VN_data_out(2539),
        VN2CN2_bit => VN_data_out(2540),
        VN2CN3_bit => VN_data_out(2541),
        VN2CN4_bit => VN_data_out(2542),
        VN2CN5_bit => VN_data_out(2543),
        VN2CN0_sign => VN_sign_out(2538),
        VN2CN1_sign => VN_sign_out(2539),
        VN2CN2_sign => VN_sign_out(2540),
        VN2CN3_sign => VN_sign_out(2541),
        VN2CN4_sign => VN_sign_out(2542),
        VN2CN5_sign => VN_sign_out(2543),
        codeword => codeword(423),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN424 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2549 downto 2544),
        Din0 => VN424_in0,
        Din1 => VN424_in1,
        Din2 => VN424_in2,
        Din3 => VN424_in3,
        Din4 => VN424_in4,
        Din5 => VN424_in5,
        VN2CN0_bit => VN_data_out(2544),
        VN2CN1_bit => VN_data_out(2545),
        VN2CN2_bit => VN_data_out(2546),
        VN2CN3_bit => VN_data_out(2547),
        VN2CN4_bit => VN_data_out(2548),
        VN2CN5_bit => VN_data_out(2549),
        VN2CN0_sign => VN_sign_out(2544),
        VN2CN1_sign => VN_sign_out(2545),
        VN2CN2_sign => VN_sign_out(2546),
        VN2CN3_sign => VN_sign_out(2547),
        VN2CN4_sign => VN_sign_out(2548),
        VN2CN5_sign => VN_sign_out(2549),
        codeword => codeword(424),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN425 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2555 downto 2550),
        Din0 => VN425_in0,
        Din1 => VN425_in1,
        Din2 => VN425_in2,
        Din3 => VN425_in3,
        Din4 => VN425_in4,
        Din5 => VN425_in5,
        VN2CN0_bit => VN_data_out(2550),
        VN2CN1_bit => VN_data_out(2551),
        VN2CN2_bit => VN_data_out(2552),
        VN2CN3_bit => VN_data_out(2553),
        VN2CN4_bit => VN_data_out(2554),
        VN2CN5_bit => VN_data_out(2555),
        VN2CN0_sign => VN_sign_out(2550),
        VN2CN1_sign => VN_sign_out(2551),
        VN2CN2_sign => VN_sign_out(2552),
        VN2CN3_sign => VN_sign_out(2553),
        VN2CN4_sign => VN_sign_out(2554),
        VN2CN5_sign => VN_sign_out(2555),
        codeword => codeword(425),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN426 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2561 downto 2556),
        Din0 => VN426_in0,
        Din1 => VN426_in1,
        Din2 => VN426_in2,
        Din3 => VN426_in3,
        Din4 => VN426_in4,
        Din5 => VN426_in5,
        VN2CN0_bit => VN_data_out(2556),
        VN2CN1_bit => VN_data_out(2557),
        VN2CN2_bit => VN_data_out(2558),
        VN2CN3_bit => VN_data_out(2559),
        VN2CN4_bit => VN_data_out(2560),
        VN2CN5_bit => VN_data_out(2561),
        VN2CN0_sign => VN_sign_out(2556),
        VN2CN1_sign => VN_sign_out(2557),
        VN2CN2_sign => VN_sign_out(2558),
        VN2CN3_sign => VN_sign_out(2559),
        VN2CN4_sign => VN_sign_out(2560),
        VN2CN5_sign => VN_sign_out(2561),
        codeword => codeword(426),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN427 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2567 downto 2562),
        Din0 => VN427_in0,
        Din1 => VN427_in1,
        Din2 => VN427_in2,
        Din3 => VN427_in3,
        Din4 => VN427_in4,
        Din5 => VN427_in5,
        VN2CN0_bit => VN_data_out(2562),
        VN2CN1_bit => VN_data_out(2563),
        VN2CN2_bit => VN_data_out(2564),
        VN2CN3_bit => VN_data_out(2565),
        VN2CN4_bit => VN_data_out(2566),
        VN2CN5_bit => VN_data_out(2567),
        VN2CN0_sign => VN_sign_out(2562),
        VN2CN1_sign => VN_sign_out(2563),
        VN2CN2_sign => VN_sign_out(2564),
        VN2CN3_sign => VN_sign_out(2565),
        VN2CN4_sign => VN_sign_out(2566),
        VN2CN5_sign => VN_sign_out(2567),
        codeword => codeword(427),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN428 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2573 downto 2568),
        Din0 => VN428_in0,
        Din1 => VN428_in1,
        Din2 => VN428_in2,
        Din3 => VN428_in3,
        Din4 => VN428_in4,
        Din5 => VN428_in5,
        VN2CN0_bit => VN_data_out(2568),
        VN2CN1_bit => VN_data_out(2569),
        VN2CN2_bit => VN_data_out(2570),
        VN2CN3_bit => VN_data_out(2571),
        VN2CN4_bit => VN_data_out(2572),
        VN2CN5_bit => VN_data_out(2573),
        VN2CN0_sign => VN_sign_out(2568),
        VN2CN1_sign => VN_sign_out(2569),
        VN2CN2_sign => VN_sign_out(2570),
        VN2CN3_sign => VN_sign_out(2571),
        VN2CN4_sign => VN_sign_out(2572),
        VN2CN5_sign => VN_sign_out(2573),
        codeword => codeword(428),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN429 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2579 downto 2574),
        Din0 => VN429_in0,
        Din1 => VN429_in1,
        Din2 => VN429_in2,
        Din3 => VN429_in3,
        Din4 => VN429_in4,
        Din5 => VN429_in5,
        VN2CN0_bit => VN_data_out(2574),
        VN2CN1_bit => VN_data_out(2575),
        VN2CN2_bit => VN_data_out(2576),
        VN2CN3_bit => VN_data_out(2577),
        VN2CN4_bit => VN_data_out(2578),
        VN2CN5_bit => VN_data_out(2579),
        VN2CN0_sign => VN_sign_out(2574),
        VN2CN1_sign => VN_sign_out(2575),
        VN2CN2_sign => VN_sign_out(2576),
        VN2CN3_sign => VN_sign_out(2577),
        VN2CN4_sign => VN_sign_out(2578),
        VN2CN5_sign => VN_sign_out(2579),
        codeword => codeword(429),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN430 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2585 downto 2580),
        Din0 => VN430_in0,
        Din1 => VN430_in1,
        Din2 => VN430_in2,
        Din3 => VN430_in3,
        Din4 => VN430_in4,
        Din5 => VN430_in5,
        VN2CN0_bit => VN_data_out(2580),
        VN2CN1_bit => VN_data_out(2581),
        VN2CN2_bit => VN_data_out(2582),
        VN2CN3_bit => VN_data_out(2583),
        VN2CN4_bit => VN_data_out(2584),
        VN2CN5_bit => VN_data_out(2585),
        VN2CN0_sign => VN_sign_out(2580),
        VN2CN1_sign => VN_sign_out(2581),
        VN2CN2_sign => VN_sign_out(2582),
        VN2CN3_sign => VN_sign_out(2583),
        VN2CN4_sign => VN_sign_out(2584),
        VN2CN5_sign => VN_sign_out(2585),
        codeword => codeword(430),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN431 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2591 downto 2586),
        Din0 => VN431_in0,
        Din1 => VN431_in1,
        Din2 => VN431_in2,
        Din3 => VN431_in3,
        Din4 => VN431_in4,
        Din5 => VN431_in5,
        VN2CN0_bit => VN_data_out(2586),
        VN2CN1_bit => VN_data_out(2587),
        VN2CN2_bit => VN_data_out(2588),
        VN2CN3_bit => VN_data_out(2589),
        VN2CN4_bit => VN_data_out(2590),
        VN2CN5_bit => VN_data_out(2591),
        VN2CN0_sign => VN_sign_out(2586),
        VN2CN1_sign => VN_sign_out(2587),
        VN2CN2_sign => VN_sign_out(2588),
        VN2CN3_sign => VN_sign_out(2589),
        VN2CN4_sign => VN_sign_out(2590),
        VN2CN5_sign => VN_sign_out(2591),
        codeword => codeword(431),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN432 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2597 downto 2592),
        Din0 => VN432_in0,
        Din1 => VN432_in1,
        Din2 => VN432_in2,
        Din3 => VN432_in3,
        Din4 => VN432_in4,
        Din5 => VN432_in5,
        VN2CN0_bit => VN_data_out(2592),
        VN2CN1_bit => VN_data_out(2593),
        VN2CN2_bit => VN_data_out(2594),
        VN2CN3_bit => VN_data_out(2595),
        VN2CN4_bit => VN_data_out(2596),
        VN2CN5_bit => VN_data_out(2597),
        VN2CN0_sign => VN_sign_out(2592),
        VN2CN1_sign => VN_sign_out(2593),
        VN2CN2_sign => VN_sign_out(2594),
        VN2CN3_sign => VN_sign_out(2595),
        VN2CN4_sign => VN_sign_out(2596),
        VN2CN5_sign => VN_sign_out(2597),
        codeword => codeword(432),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN433 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2603 downto 2598),
        Din0 => VN433_in0,
        Din1 => VN433_in1,
        Din2 => VN433_in2,
        Din3 => VN433_in3,
        Din4 => VN433_in4,
        Din5 => VN433_in5,
        VN2CN0_bit => VN_data_out(2598),
        VN2CN1_bit => VN_data_out(2599),
        VN2CN2_bit => VN_data_out(2600),
        VN2CN3_bit => VN_data_out(2601),
        VN2CN4_bit => VN_data_out(2602),
        VN2CN5_bit => VN_data_out(2603),
        VN2CN0_sign => VN_sign_out(2598),
        VN2CN1_sign => VN_sign_out(2599),
        VN2CN2_sign => VN_sign_out(2600),
        VN2CN3_sign => VN_sign_out(2601),
        VN2CN4_sign => VN_sign_out(2602),
        VN2CN5_sign => VN_sign_out(2603),
        codeword => codeword(433),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN434 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2609 downto 2604),
        Din0 => VN434_in0,
        Din1 => VN434_in1,
        Din2 => VN434_in2,
        Din3 => VN434_in3,
        Din4 => VN434_in4,
        Din5 => VN434_in5,
        VN2CN0_bit => VN_data_out(2604),
        VN2CN1_bit => VN_data_out(2605),
        VN2CN2_bit => VN_data_out(2606),
        VN2CN3_bit => VN_data_out(2607),
        VN2CN4_bit => VN_data_out(2608),
        VN2CN5_bit => VN_data_out(2609),
        VN2CN0_sign => VN_sign_out(2604),
        VN2CN1_sign => VN_sign_out(2605),
        VN2CN2_sign => VN_sign_out(2606),
        VN2CN3_sign => VN_sign_out(2607),
        VN2CN4_sign => VN_sign_out(2608),
        VN2CN5_sign => VN_sign_out(2609),
        codeword => codeword(434),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN435 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2615 downto 2610),
        Din0 => VN435_in0,
        Din1 => VN435_in1,
        Din2 => VN435_in2,
        Din3 => VN435_in3,
        Din4 => VN435_in4,
        Din5 => VN435_in5,
        VN2CN0_bit => VN_data_out(2610),
        VN2CN1_bit => VN_data_out(2611),
        VN2CN2_bit => VN_data_out(2612),
        VN2CN3_bit => VN_data_out(2613),
        VN2CN4_bit => VN_data_out(2614),
        VN2CN5_bit => VN_data_out(2615),
        VN2CN0_sign => VN_sign_out(2610),
        VN2CN1_sign => VN_sign_out(2611),
        VN2CN2_sign => VN_sign_out(2612),
        VN2CN3_sign => VN_sign_out(2613),
        VN2CN4_sign => VN_sign_out(2614),
        VN2CN5_sign => VN_sign_out(2615),
        codeword => codeword(435),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN436 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2621 downto 2616),
        Din0 => VN436_in0,
        Din1 => VN436_in1,
        Din2 => VN436_in2,
        Din3 => VN436_in3,
        Din4 => VN436_in4,
        Din5 => VN436_in5,
        VN2CN0_bit => VN_data_out(2616),
        VN2CN1_bit => VN_data_out(2617),
        VN2CN2_bit => VN_data_out(2618),
        VN2CN3_bit => VN_data_out(2619),
        VN2CN4_bit => VN_data_out(2620),
        VN2CN5_bit => VN_data_out(2621),
        VN2CN0_sign => VN_sign_out(2616),
        VN2CN1_sign => VN_sign_out(2617),
        VN2CN2_sign => VN_sign_out(2618),
        VN2CN3_sign => VN_sign_out(2619),
        VN2CN4_sign => VN_sign_out(2620),
        VN2CN5_sign => VN_sign_out(2621),
        codeword => codeword(436),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN437 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2627 downto 2622),
        Din0 => VN437_in0,
        Din1 => VN437_in1,
        Din2 => VN437_in2,
        Din3 => VN437_in3,
        Din4 => VN437_in4,
        Din5 => VN437_in5,
        VN2CN0_bit => VN_data_out(2622),
        VN2CN1_bit => VN_data_out(2623),
        VN2CN2_bit => VN_data_out(2624),
        VN2CN3_bit => VN_data_out(2625),
        VN2CN4_bit => VN_data_out(2626),
        VN2CN5_bit => VN_data_out(2627),
        VN2CN0_sign => VN_sign_out(2622),
        VN2CN1_sign => VN_sign_out(2623),
        VN2CN2_sign => VN_sign_out(2624),
        VN2CN3_sign => VN_sign_out(2625),
        VN2CN4_sign => VN_sign_out(2626),
        VN2CN5_sign => VN_sign_out(2627),
        codeword => codeword(437),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN438 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2633 downto 2628),
        Din0 => VN438_in0,
        Din1 => VN438_in1,
        Din2 => VN438_in2,
        Din3 => VN438_in3,
        Din4 => VN438_in4,
        Din5 => VN438_in5,
        VN2CN0_bit => VN_data_out(2628),
        VN2CN1_bit => VN_data_out(2629),
        VN2CN2_bit => VN_data_out(2630),
        VN2CN3_bit => VN_data_out(2631),
        VN2CN4_bit => VN_data_out(2632),
        VN2CN5_bit => VN_data_out(2633),
        VN2CN0_sign => VN_sign_out(2628),
        VN2CN1_sign => VN_sign_out(2629),
        VN2CN2_sign => VN_sign_out(2630),
        VN2CN3_sign => VN_sign_out(2631),
        VN2CN4_sign => VN_sign_out(2632),
        VN2CN5_sign => VN_sign_out(2633),
        codeword => codeword(438),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN439 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2639 downto 2634),
        Din0 => VN439_in0,
        Din1 => VN439_in1,
        Din2 => VN439_in2,
        Din3 => VN439_in3,
        Din4 => VN439_in4,
        Din5 => VN439_in5,
        VN2CN0_bit => VN_data_out(2634),
        VN2CN1_bit => VN_data_out(2635),
        VN2CN2_bit => VN_data_out(2636),
        VN2CN3_bit => VN_data_out(2637),
        VN2CN4_bit => VN_data_out(2638),
        VN2CN5_bit => VN_data_out(2639),
        VN2CN0_sign => VN_sign_out(2634),
        VN2CN1_sign => VN_sign_out(2635),
        VN2CN2_sign => VN_sign_out(2636),
        VN2CN3_sign => VN_sign_out(2637),
        VN2CN4_sign => VN_sign_out(2638),
        VN2CN5_sign => VN_sign_out(2639),
        codeword => codeword(439),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN440 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2645 downto 2640),
        Din0 => VN440_in0,
        Din1 => VN440_in1,
        Din2 => VN440_in2,
        Din3 => VN440_in3,
        Din4 => VN440_in4,
        Din5 => VN440_in5,
        VN2CN0_bit => VN_data_out(2640),
        VN2CN1_bit => VN_data_out(2641),
        VN2CN2_bit => VN_data_out(2642),
        VN2CN3_bit => VN_data_out(2643),
        VN2CN4_bit => VN_data_out(2644),
        VN2CN5_bit => VN_data_out(2645),
        VN2CN0_sign => VN_sign_out(2640),
        VN2CN1_sign => VN_sign_out(2641),
        VN2CN2_sign => VN_sign_out(2642),
        VN2CN3_sign => VN_sign_out(2643),
        VN2CN4_sign => VN_sign_out(2644),
        VN2CN5_sign => VN_sign_out(2645),
        codeword => codeword(440),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN441 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2651 downto 2646),
        Din0 => VN441_in0,
        Din1 => VN441_in1,
        Din2 => VN441_in2,
        Din3 => VN441_in3,
        Din4 => VN441_in4,
        Din5 => VN441_in5,
        VN2CN0_bit => VN_data_out(2646),
        VN2CN1_bit => VN_data_out(2647),
        VN2CN2_bit => VN_data_out(2648),
        VN2CN3_bit => VN_data_out(2649),
        VN2CN4_bit => VN_data_out(2650),
        VN2CN5_bit => VN_data_out(2651),
        VN2CN0_sign => VN_sign_out(2646),
        VN2CN1_sign => VN_sign_out(2647),
        VN2CN2_sign => VN_sign_out(2648),
        VN2CN3_sign => VN_sign_out(2649),
        VN2CN4_sign => VN_sign_out(2650),
        VN2CN5_sign => VN_sign_out(2651),
        codeword => codeword(441),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN442 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2657 downto 2652),
        Din0 => VN442_in0,
        Din1 => VN442_in1,
        Din2 => VN442_in2,
        Din3 => VN442_in3,
        Din4 => VN442_in4,
        Din5 => VN442_in5,
        VN2CN0_bit => VN_data_out(2652),
        VN2CN1_bit => VN_data_out(2653),
        VN2CN2_bit => VN_data_out(2654),
        VN2CN3_bit => VN_data_out(2655),
        VN2CN4_bit => VN_data_out(2656),
        VN2CN5_bit => VN_data_out(2657),
        VN2CN0_sign => VN_sign_out(2652),
        VN2CN1_sign => VN_sign_out(2653),
        VN2CN2_sign => VN_sign_out(2654),
        VN2CN3_sign => VN_sign_out(2655),
        VN2CN4_sign => VN_sign_out(2656),
        VN2CN5_sign => VN_sign_out(2657),
        codeword => codeword(442),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN443 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2663 downto 2658),
        Din0 => VN443_in0,
        Din1 => VN443_in1,
        Din2 => VN443_in2,
        Din3 => VN443_in3,
        Din4 => VN443_in4,
        Din5 => VN443_in5,
        VN2CN0_bit => VN_data_out(2658),
        VN2CN1_bit => VN_data_out(2659),
        VN2CN2_bit => VN_data_out(2660),
        VN2CN3_bit => VN_data_out(2661),
        VN2CN4_bit => VN_data_out(2662),
        VN2CN5_bit => VN_data_out(2663),
        VN2CN0_sign => VN_sign_out(2658),
        VN2CN1_sign => VN_sign_out(2659),
        VN2CN2_sign => VN_sign_out(2660),
        VN2CN3_sign => VN_sign_out(2661),
        VN2CN4_sign => VN_sign_out(2662),
        VN2CN5_sign => VN_sign_out(2663),
        codeword => codeword(443),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN444 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2669 downto 2664),
        Din0 => VN444_in0,
        Din1 => VN444_in1,
        Din2 => VN444_in2,
        Din3 => VN444_in3,
        Din4 => VN444_in4,
        Din5 => VN444_in5,
        VN2CN0_bit => VN_data_out(2664),
        VN2CN1_bit => VN_data_out(2665),
        VN2CN2_bit => VN_data_out(2666),
        VN2CN3_bit => VN_data_out(2667),
        VN2CN4_bit => VN_data_out(2668),
        VN2CN5_bit => VN_data_out(2669),
        VN2CN0_sign => VN_sign_out(2664),
        VN2CN1_sign => VN_sign_out(2665),
        VN2CN2_sign => VN_sign_out(2666),
        VN2CN3_sign => VN_sign_out(2667),
        VN2CN4_sign => VN_sign_out(2668),
        VN2CN5_sign => VN_sign_out(2669),
        codeword => codeword(444),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN445 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2675 downto 2670),
        Din0 => VN445_in0,
        Din1 => VN445_in1,
        Din2 => VN445_in2,
        Din3 => VN445_in3,
        Din4 => VN445_in4,
        Din5 => VN445_in5,
        VN2CN0_bit => VN_data_out(2670),
        VN2CN1_bit => VN_data_out(2671),
        VN2CN2_bit => VN_data_out(2672),
        VN2CN3_bit => VN_data_out(2673),
        VN2CN4_bit => VN_data_out(2674),
        VN2CN5_bit => VN_data_out(2675),
        VN2CN0_sign => VN_sign_out(2670),
        VN2CN1_sign => VN_sign_out(2671),
        VN2CN2_sign => VN_sign_out(2672),
        VN2CN3_sign => VN_sign_out(2673),
        VN2CN4_sign => VN_sign_out(2674),
        VN2CN5_sign => VN_sign_out(2675),
        codeword => codeword(445),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN446 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2681 downto 2676),
        Din0 => VN446_in0,
        Din1 => VN446_in1,
        Din2 => VN446_in2,
        Din3 => VN446_in3,
        Din4 => VN446_in4,
        Din5 => VN446_in5,
        VN2CN0_bit => VN_data_out(2676),
        VN2CN1_bit => VN_data_out(2677),
        VN2CN2_bit => VN_data_out(2678),
        VN2CN3_bit => VN_data_out(2679),
        VN2CN4_bit => VN_data_out(2680),
        VN2CN5_bit => VN_data_out(2681),
        VN2CN0_sign => VN_sign_out(2676),
        VN2CN1_sign => VN_sign_out(2677),
        VN2CN2_sign => VN_sign_out(2678),
        VN2CN3_sign => VN_sign_out(2679),
        VN2CN4_sign => VN_sign_out(2680),
        VN2CN5_sign => VN_sign_out(2681),
        codeword => codeword(446),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN447 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2687 downto 2682),
        Din0 => VN447_in0,
        Din1 => VN447_in1,
        Din2 => VN447_in2,
        Din3 => VN447_in3,
        Din4 => VN447_in4,
        Din5 => VN447_in5,
        VN2CN0_bit => VN_data_out(2682),
        VN2CN1_bit => VN_data_out(2683),
        VN2CN2_bit => VN_data_out(2684),
        VN2CN3_bit => VN_data_out(2685),
        VN2CN4_bit => VN_data_out(2686),
        VN2CN5_bit => VN_data_out(2687),
        VN2CN0_sign => VN_sign_out(2682),
        VN2CN1_sign => VN_sign_out(2683),
        VN2CN2_sign => VN_sign_out(2684),
        VN2CN3_sign => VN_sign_out(2685),
        VN2CN4_sign => VN_sign_out(2686),
        VN2CN5_sign => VN_sign_out(2687),
        codeword => codeword(447),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN448 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2693 downto 2688),
        Din0 => VN448_in0,
        Din1 => VN448_in1,
        Din2 => VN448_in2,
        Din3 => VN448_in3,
        Din4 => VN448_in4,
        Din5 => VN448_in5,
        VN2CN0_bit => VN_data_out(2688),
        VN2CN1_bit => VN_data_out(2689),
        VN2CN2_bit => VN_data_out(2690),
        VN2CN3_bit => VN_data_out(2691),
        VN2CN4_bit => VN_data_out(2692),
        VN2CN5_bit => VN_data_out(2693),
        VN2CN0_sign => VN_sign_out(2688),
        VN2CN1_sign => VN_sign_out(2689),
        VN2CN2_sign => VN_sign_out(2690),
        VN2CN3_sign => VN_sign_out(2691),
        VN2CN4_sign => VN_sign_out(2692),
        VN2CN5_sign => VN_sign_out(2693),
        codeword => codeword(448),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN449 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2699 downto 2694),
        Din0 => VN449_in0,
        Din1 => VN449_in1,
        Din2 => VN449_in2,
        Din3 => VN449_in3,
        Din4 => VN449_in4,
        Din5 => VN449_in5,
        VN2CN0_bit => VN_data_out(2694),
        VN2CN1_bit => VN_data_out(2695),
        VN2CN2_bit => VN_data_out(2696),
        VN2CN3_bit => VN_data_out(2697),
        VN2CN4_bit => VN_data_out(2698),
        VN2CN5_bit => VN_data_out(2699),
        VN2CN0_sign => VN_sign_out(2694),
        VN2CN1_sign => VN_sign_out(2695),
        VN2CN2_sign => VN_sign_out(2696),
        VN2CN3_sign => VN_sign_out(2697),
        VN2CN4_sign => VN_sign_out(2698),
        VN2CN5_sign => VN_sign_out(2699),
        codeword => codeword(449),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN450 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2705 downto 2700),
        Din0 => VN450_in0,
        Din1 => VN450_in1,
        Din2 => VN450_in2,
        Din3 => VN450_in3,
        Din4 => VN450_in4,
        Din5 => VN450_in5,
        VN2CN0_bit => VN_data_out(2700),
        VN2CN1_bit => VN_data_out(2701),
        VN2CN2_bit => VN_data_out(2702),
        VN2CN3_bit => VN_data_out(2703),
        VN2CN4_bit => VN_data_out(2704),
        VN2CN5_bit => VN_data_out(2705),
        VN2CN0_sign => VN_sign_out(2700),
        VN2CN1_sign => VN_sign_out(2701),
        VN2CN2_sign => VN_sign_out(2702),
        VN2CN3_sign => VN_sign_out(2703),
        VN2CN4_sign => VN_sign_out(2704),
        VN2CN5_sign => VN_sign_out(2705),
        codeword => codeword(450),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN451 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2711 downto 2706),
        Din0 => VN451_in0,
        Din1 => VN451_in1,
        Din2 => VN451_in2,
        Din3 => VN451_in3,
        Din4 => VN451_in4,
        Din5 => VN451_in5,
        VN2CN0_bit => VN_data_out(2706),
        VN2CN1_bit => VN_data_out(2707),
        VN2CN2_bit => VN_data_out(2708),
        VN2CN3_bit => VN_data_out(2709),
        VN2CN4_bit => VN_data_out(2710),
        VN2CN5_bit => VN_data_out(2711),
        VN2CN0_sign => VN_sign_out(2706),
        VN2CN1_sign => VN_sign_out(2707),
        VN2CN2_sign => VN_sign_out(2708),
        VN2CN3_sign => VN_sign_out(2709),
        VN2CN4_sign => VN_sign_out(2710),
        VN2CN5_sign => VN_sign_out(2711),
        codeword => codeword(451),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN452 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2717 downto 2712),
        Din0 => VN452_in0,
        Din1 => VN452_in1,
        Din2 => VN452_in2,
        Din3 => VN452_in3,
        Din4 => VN452_in4,
        Din5 => VN452_in5,
        VN2CN0_bit => VN_data_out(2712),
        VN2CN1_bit => VN_data_out(2713),
        VN2CN2_bit => VN_data_out(2714),
        VN2CN3_bit => VN_data_out(2715),
        VN2CN4_bit => VN_data_out(2716),
        VN2CN5_bit => VN_data_out(2717),
        VN2CN0_sign => VN_sign_out(2712),
        VN2CN1_sign => VN_sign_out(2713),
        VN2CN2_sign => VN_sign_out(2714),
        VN2CN3_sign => VN_sign_out(2715),
        VN2CN4_sign => VN_sign_out(2716),
        VN2CN5_sign => VN_sign_out(2717),
        codeword => codeword(452),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN453 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2723 downto 2718),
        Din0 => VN453_in0,
        Din1 => VN453_in1,
        Din2 => VN453_in2,
        Din3 => VN453_in3,
        Din4 => VN453_in4,
        Din5 => VN453_in5,
        VN2CN0_bit => VN_data_out(2718),
        VN2CN1_bit => VN_data_out(2719),
        VN2CN2_bit => VN_data_out(2720),
        VN2CN3_bit => VN_data_out(2721),
        VN2CN4_bit => VN_data_out(2722),
        VN2CN5_bit => VN_data_out(2723),
        VN2CN0_sign => VN_sign_out(2718),
        VN2CN1_sign => VN_sign_out(2719),
        VN2CN2_sign => VN_sign_out(2720),
        VN2CN3_sign => VN_sign_out(2721),
        VN2CN4_sign => VN_sign_out(2722),
        VN2CN5_sign => VN_sign_out(2723),
        codeword => codeword(453),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN454 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2729 downto 2724),
        Din0 => VN454_in0,
        Din1 => VN454_in1,
        Din2 => VN454_in2,
        Din3 => VN454_in3,
        Din4 => VN454_in4,
        Din5 => VN454_in5,
        VN2CN0_bit => VN_data_out(2724),
        VN2CN1_bit => VN_data_out(2725),
        VN2CN2_bit => VN_data_out(2726),
        VN2CN3_bit => VN_data_out(2727),
        VN2CN4_bit => VN_data_out(2728),
        VN2CN5_bit => VN_data_out(2729),
        VN2CN0_sign => VN_sign_out(2724),
        VN2CN1_sign => VN_sign_out(2725),
        VN2CN2_sign => VN_sign_out(2726),
        VN2CN3_sign => VN_sign_out(2727),
        VN2CN4_sign => VN_sign_out(2728),
        VN2CN5_sign => VN_sign_out(2729),
        codeword => codeword(454),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN455 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2735 downto 2730),
        Din0 => VN455_in0,
        Din1 => VN455_in1,
        Din2 => VN455_in2,
        Din3 => VN455_in3,
        Din4 => VN455_in4,
        Din5 => VN455_in5,
        VN2CN0_bit => VN_data_out(2730),
        VN2CN1_bit => VN_data_out(2731),
        VN2CN2_bit => VN_data_out(2732),
        VN2CN3_bit => VN_data_out(2733),
        VN2CN4_bit => VN_data_out(2734),
        VN2CN5_bit => VN_data_out(2735),
        VN2CN0_sign => VN_sign_out(2730),
        VN2CN1_sign => VN_sign_out(2731),
        VN2CN2_sign => VN_sign_out(2732),
        VN2CN3_sign => VN_sign_out(2733),
        VN2CN4_sign => VN_sign_out(2734),
        VN2CN5_sign => VN_sign_out(2735),
        codeword => codeword(455),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN456 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2741 downto 2736),
        Din0 => VN456_in0,
        Din1 => VN456_in1,
        Din2 => VN456_in2,
        Din3 => VN456_in3,
        Din4 => VN456_in4,
        Din5 => VN456_in5,
        VN2CN0_bit => VN_data_out(2736),
        VN2CN1_bit => VN_data_out(2737),
        VN2CN2_bit => VN_data_out(2738),
        VN2CN3_bit => VN_data_out(2739),
        VN2CN4_bit => VN_data_out(2740),
        VN2CN5_bit => VN_data_out(2741),
        VN2CN0_sign => VN_sign_out(2736),
        VN2CN1_sign => VN_sign_out(2737),
        VN2CN2_sign => VN_sign_out(2738),
        VN2CN3_sign => VN_sign_out(2739),
        VN2CN4_sign => VN_sign_out(2740),
        VN2CN5_sign => VN_sign_out(2741),
        codeword => codeword(456),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN457 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2747 downto 2742),
        Din0 => VN457_in0,
        Din1 => VN457_in1,
        Din2 => VN457_in2,
        Din3 => VN457_in3,
        Din4 => VN457_in4,
        Din5 => VN457_in5,
        VN2CN0_bit => VN_data_out(2742),
        VN2CN1_bit => VN_data_out(2743),
        VN2CN2_bit => VN_data_out(2744),
        VN2CN3_bit => VN_data_out(2745),
        VN2CN4_bit => VN_data_out(2746),
        VN2CN5_bit => VN_data_out(2747),
        VN2CN0_sign => VN_sign_out(2742),
        VN2CN1_sign => VN_sign_out(2743),
        VN2CN2_sign => VN_sign_out(2744),
        VN2CN3_sign => VN_sign_out(2745),
        VN2CN4_sign => VN_sign_out(2746),
        VN2CN5_sign => VN_sign_out(2747),
        codeword => codeword(457),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN458 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2753 downto 2748),
        Din0 => VN458_in0,
        Din1 => VN458_in1,
        Din2 => VN458_in2,
        Din3 => VN458_in3,
        Din4 => VN458_in4,
        Din5 => VN458_in5,
        VN2CN0_bit => VN_data_out(2748),
        VN2CN1_bit => VN_data_out(2749),
        VN2CN2_bit => VN_data_out(2750),
        VN2CN3_bit => VN_data_out(2751),
        VN2CN4_bit => VN_data_out(2752),
        VN2CN5_bit => VN_data_out(2753),
        VN2CN0_sign => VN_sign_out(2748),
        VN2CN1_sign => VN_sign_out(2749),
        VN2CN2_sign => VN_sign_out(2750),
        VN2CN3_sign => VN_sign_out(2751),
        VN2CN4_sign => VN_sign_out(2752),
        VN2CN5_sign => VN_sign_out(2753),
        codeword => codeword(458),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN459 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2759 downto 2754),
        Din0 => VN459_in0,
        Din1 => VN459_in1,
        Din2 => VN459_in2,
        Din3 => VN459_in3,
        Din4 => VN459_in4,
        Din5 => VN459_in5,
        VN2CN0_bit => VN_data_out(2754),
        VN2CN1_bit => VN_data_out(2755),
        VN2CN2_bit => VN_data_out(2756),
        VN2CN3_bit => VN_data_out(2757),
        VN2CN4_bit => VN_data_out(2758),
        VN2CN5_bit => VN_data_out(2759),
        VN2CN0_sign => VN_sign_out(2754),
        VN2CN1_sign => VN_sign_out(2755),
        VN2CN2_sign => VN_sign_out(2756),
        VN2CN3_sign => VN_sign_out(2757),
        VN2CN4_sign => VN_sign_out(2758),
        VN2CN5_sign => VN_sign_out(2759),
        codeword => codeword(459),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN460 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2765 downto 2760),
        Din0 => VN460_in0,
        Din1 => VN460_in1,
        Din2 => VN460_in2,
        Din3 => VN460_in3,
        Din4 => VN460_in4,
        Din5 => VN460_in5,
        VN2CN0_bit => VN_data_out(2760),
        VN2CN1_bit => VN_data_out(2761),
        VN2CN2_bit => VN_data_out(2762),
        VN2CN3_bit => VN_data_out(2763),
        VN2CN4_bit => VN_data_out(2764),
        VN2CN5_bit => VN_data_out(2765),
        VN2CN0_sign => VN_sign_out(2760),
        VN2CN1_sign => VN_sign_out(2761),
        VN2CN2_sign => VN_sign_out(2762),
        VN2CN3_sign => VN_sign_out(2763),
        VN2CN4_sign => VN_sign_out(2764),
        VN2CN5_sign => VN_sign_out(2765),
        codeword => codeword(460),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN461 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2771 downto 2766),
        Din0 => VN461_in0,
        Din1 => VN461_in1,
        Din2 => VN461_in2,
        Din3 => VN461_in3,
        Din4 => VN461_in4,
        Din5 => VN461_in5,
        VN2CN0_bit => VN_data_out(2766),
        VN2CN1_bit => VN_data_out(2767),
        VN2CN2_bit => VN_data_out(2768),
        VN2CN3_bit => VN_data_out(2769),
        VN2CN4_bit => VN_data_out(2770),
        VN2CN5_bit => VN_data_out(2771),
        VN2CN0_sign => VN_sign_out(2766),
        VN2CN1_sign => VN_sign_out(2767),
        VN2CN2_sign => VN_sign_out(2768),
        VN2CN3_sign => VN_sign_out(2769),
        VN2CN4_sign => VN_sign_out(2770),
        VN2CN5_sign => VN_sign_out(2771),
        codeword => codeword(461),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN462 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2777 downto 2772),
        Din0 => VN462_in0,
        Din1 => VN462_in1,
        Din2 => VN462_in2,
        Din3 => VN462_in3,
        Din4 => VN462_in4,
        Din5 => VN462_in5,
        VN2CN0_bit => VN_data_out(2772),
        VN2CN1_bit => VN_data_out(2773),
        VN2CN2_bit => VN_data_out(2774),
        VN2CN3_bit => VN_data_out(2775),
        VN2CN4_bit => VN_data_out(2776),
        VN2CN5_bit => VN_data_out(2777),
        VN2CN0_sign => VN_sign_out(2772),
        VN2CN1_sign => VN_sign_out(2773),
        VN2CN2_sign => VN_sign_out(2774),
        VN2CN3_sign => VN_sign_out(2775),
        VN2CN4_sign => VN_sign_out(2776),
        VN2CN5_sign => VN_sign_out(2777),
        codeword => codeword(462),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN463 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2783 downto 2778),
        Din0 => VN463_in0,
        Din1 => VN463_in1,
        Din2 => VN463_in2,
        Din3 => VN463_in3,
        Din4 => VN463_in4,
        Din5 => VN463_in5,
        VN2CN0_bit => VN_data_out(2778),
        VN2CN1_bit => VN_data_out(2779),
        VN2CN2_bit => VN_data_out(2780),
        VN2CN3_bit => VN_data_out(2781),
        VN2CN4_bit => VN_data_out(2782),
        VN2CN5_bit => VN_data_out(2783),
        VN2CN0_sign => VN_sign_out(2778),
        VN2CN1_sign => VN_sign_out(2779),
        VN2CN2_sign => VN_sign_out(2780),
        VN2CN3_sign => VN_sign_out(2781),
        VN2CN4_sign => VN_sign_out(2782),
        VN2CN5_sign => VN_sign_out(2783),
        codeword => codeword(463),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN464 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2789 downto 2784),
        Din0 => VN464_in0,
        Din1 => VN464_in1,
        Din2 => VN464_in2,
        Din3 => VN464_in3,
        Din4 => VN464_in4,
        Din5 => VN464_in5,
        VN2CN0_bit => VN_data_out(2784),
        VN2CN1_bit => VN_data_out(2785),
        VN2CN2_bit => VN_data_out(2786),
        VN2CN3_bit => VN_data_out(2787),
        VN2CN4_bit => VN_data_out(2788),
        VN2CN5_bit => VN_data_out(2789),
        VN2CN0_sign => VN_sign_out(2784),
        VN2CN1_sign => VN_sign_out(2785),
        VN2CN2_sign => VN_sign_out(2786),
        VN2CN3_sign => VN_sign_out(2787),
        VN2CN4_sign => VN_sign_out(2788),
        VN2CN5_sign => VN_sign_out(2789),
        codeword => codeword(464),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN465 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2795 downto 2790),
        Din0 => VN465_in0,
        Din1 => VN465_in1,
        Din2 => VN465_in2,
        Din3 => VN465_in3,
        Din4 => VN465_in4,
        Din5 => VN465_in5,
        VN2CN0_bit => VN_data_out(2790),
        VN2CN1_bit => VN_data_out(2791),
        VN2CN2_bit => VN_data_out(2792),
        VN2CN3_bit => VN_data_out(2793),
        VN2CN4_bit => VN_data_out(2794),
        VN2CN5_bit => VN_data_out(2795),
        VN2CN0_sign => VN_sign_out(2790),
        VN2CN1_sign => VN_sign_out(2791),
        VN2CN2_sign => VN_sign_out(2792),
        VN2CN3_sign => VN_sign_out(2793),
        VN2CN4_sign => VN_sign_out(2794),
        VN2CN5_sign => VN_sign_out(2795),
        codeword => codeword(465),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN466 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2801 downto 2796),
        Din0 => VN466_in0,
        Din1 => VN466_in1,
        Din2 => VN466_in2,
        Din3 => VN466_in3,
        Din4 => VN466_in4,
        Din5 => VN466_in5,
        VN2CN0_bit => VN_data_out(2796),
        VN2CN1_bit => VN_data_out(2797),
        VN2CN2_bit => VN_data_out(2798),
        VN2CN3_bit => VN_data_out(2799),
        VN2CN4_bit => VN_data_out(2800),
        VN2CN5_bit => VN_data_out(2801),
        VN2CN0_sign => VN_sign_out(2796),
        VN2CN1_sign => VN_sign_out(2797),
        VN2CN2_sign => VN_sign_out(2798),
        VN2CN3_sign => VN_sign_out(2799),
        VN2CN4_sign => VN_sign_out(2800),
        VN2CN5_sign => VN_sign_out(2801),
        codeword => codeword(466),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN467 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2807 downto 2802),
        Din0 => VN467_in0,
        Din1 => VN467_in1,
        Din2 => VN467_in2,
        Din3 => VN467_in3,
        Din4 => VN467_in4,
        Din5 => VN467_in5,
        VN2CN0_bit => VN_data_out(2802),
        VN2CN1_bit => VN_data_out(2803),
        VN2CN2_bit => VN_data_out(2804),
        VN2CN3_bit => VN_data_out(2805),
        VN2CN4_bit => VN_data_out(2806),
        VN2CN5_bit => VN_data_out(2807),
        VN2CN0_sign => VN_sign_out(2802),
        VN2CN1_sign => VN_sign_out(2803),
        VN2CN2_sign => VN_sign_out(2804),
        VN2CN3_sign => VN_sign_out(2805),
        VN2CN4_sign => VN_sign_out(2806),
        VN2CN5_sign => VN_sign_out(2807),
        codeword => codeword(467),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN468 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2813 downto 2808),
        Din0 => VN468_in0,
        Din1 => VN468_in1,
        Din2 => VN468_in2,
        Din3 => VN468_in3,
        Din4 => VN468_in4,
        Din5 => VN468_in5,
        VN2CN0_bit => VN_data_out(2808),
        VN2CN1_bit => VN_data_out(2809),
        VN2CN2_bit => VN_data_out(2810),
        VN2CN3_bit => VN_data_out(2811),
        VN2CN4_bit => VN_data_out(2812),
        VN2CN5_bit => VN_data_out(2813),
        VN2CN0_sign => VN_sign_out(2808),
        VN2CN1_sign => VN_sign_out(2809),
        VN2CN2_sign => VN_sign_out(2810),
        VN2CN3_sign => VN_sign_out(2811),
        VN2CN4_sign => VN_sign_out(2812),
        VN2CN5_sign => VN_sign_out(2813),
        codeword => codeword(468),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN469 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2819 downto 2814),
        Din0 => VN469_in0,
        Din1 => VN469_in1,
        Din2 => VN469_in2,
        Din3 => VN469_in3,
        Din4 => VN469_in4,
        Din5 => VN469_in5,
        VN2CN0_bit => VN_data_out(2814),
        VN2CN1_bit => VN_data_out(2815),
        VN2CN2_bit => VN_data_out(2816),
        VN2CN3_bit => VN_data_out(2817),
        VN2CN4_bit => VN_data_out(2818),
        VN2CN5_bit => VN_data_out(2819),
        VN2CN0_sign => VN_sign_out(2814),
        VN2CN1_sign => VN_sign_out(2815),
        VN2CN2_sign => VN_sign_out(2816),
        VN2CN3_sign => VN_sign_out(2817),
        VN2CN4_sign => VN_sign_out(2818),
        VN2CN5_sign => VN_sign_out(2819),
        codeword => codeword(469),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN470 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2825 downto 2820),
        Din0 => VN470_in0,
        Din1 => VN470_in1,
        Din2 => VN470_in2,
        Din3 => VN470_in3,
        Din4 => VN470_in4,
        Din5 => VN470_in5,
        VN2CN0_bit => VN_data_out(2820),
        VN2CN1_bit => VN_data_out(2821),
        VN2CN2_bit => VN_data_out(2822),
        VN2CN3_bit => VN_data_out(2823),
        VN2CN4_bit => VN_data_out(2824),
        VN2CN5_bit => VN_data_out(2825),
        VN2CN0_sign => VN_sign_out(2820),
        VN2CN1_sign => VN_sign_out(2821),
        VN2CN2_sign => VN_sign_out(2822),
        VN2CN3_sign => VN_sign_out(2823),
        VN2CN4_sign => VN_sign_out(2824),
        VN2CN5_sign => VN_sign_out(2825),
        codeword => codeword(470),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN471 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2831 downto 2826),
        Din0 => VN471_in0,
        Din1 => VN471_in1,
        Din2 => VN471_in2,
        Din3 => VN471_in3,
        Din4 => VN471_in4,
        Din5 => VN471_in5,
        VN2CN0_bit => VN_data_out(2826),
        VN2CN1_bit => VN_data_out(2827),
        VN2CN2_bit => VN_data_out(2828),
        VN2CN3_bit => VN_data_out(2829),
        VN2CN4_bit => VN_data_out(2830),
        VN2CN5_bit => VN_data_out(2831),
        VN2CN0_sign => VN_sign_out(2826),
        VN2CN1_sign => VN_sign_out(2827),
        VN2CN2_sign => VN_sign_out(2828),
        VN2CN3_sign => VN_sign_out(2829),
        VN2CN4_sign => VN_sign_out(2830),
        VN2CN5_sign => VN_sign_out(2831),
        codeword => codeword(471),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN472 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2837 downto 2832),
        Din0 => VN472_in0,
        Din1 => VN472_in1,
        Din2 => VN472_in2,
        Din3 => VN472_in3,
        Din4 => VN472_in4,
        Din5 => VN472_in5,
        VN2CN0_bit => VN_data_out(2832),
        VN2CN1_bit => VN_data_out(2833),
        VN2CN2_bit => VN_data_out(2834),
        VN2CN3_bit => VN_data_out(2835),
        VN2CN4_bit => VN_data_out(2836),
        VN2CN5_bit => VN_data_out(2837),
        VN2CN0_sign => VN_sign_out(2832),
        VN2CN1_sign => VN_sign_out(2833),
        VN2CN2_sign => VN_sign_out(2834),
        VN2CN3_sign => VN_sign_out(2835),
        VN2CN4_sign => VN_sign_out(2836),
        VN2CN5_sign => VN_sign_out(2837),
        codeword => codeword(472),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN473 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2843 downto 2838),
        Din0 => VN473_in0,
        Din1 => VN473_in1,
        Din2 => VN473_in2,
        Din3 => VN473_in3,
        Din4 => VN473_in4,
        Din5 => VN473_in5,
        VN2CN0_bit => VN_data_out(2838),
        VN2CN1_bit => VN_data_out(2839),
        VN2CN2_bit => VN_data_out(2840),
        VN2CN3_bit => VN_data_out(2841),
        VN2CN4_bit => VN_data_out(2842),
        VN2CN5_bit => VN_data_out(2843),
        VN2CN0_sign => VN_sign_out(2838),
        VN2CN1_sign => VN_sign_out(2839),
        VN2CN2_sign => VN_sign_out(2840),
        VN2CN3_sign => VN_sign_out(2841),
        VN2CN4_sign => VN_sign_out(2842),
        VN2CN5_sign => VN_sign_out(2843),
        codeword => codeword(473),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN474 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2849 downto 2844),
        Din0 => VN474_in0,
        Din1 => VN474_in1,
        Din2 => VN474_in2,
        Din3 => VN474_in3,
        Din4 => VN474_in4,
        Din5 => VN474_in5,
        VN2CN0_bit => VN_data_out(2844),
        VN2CN1_bit => VN_data_out(2845),
        VN2CN2_bit => VN_data_out(2846),
        VN2CN3_bit => VN_data_out(2847),
        VN2CN4_bit => VN_data_out(2848),
        VN2CN5_bit => VN_data_out(2849),
        VN2CN0_sign => VN_sign_out(2844),
        VN2CN1_sign => VN_sign_out(2845),
        VN2CN2_sign => VN_sign_out(2846),
        VN2CN3_sign => VN_sign_out(2847),
        VN2CN4_sign => VN_sign_out(2848),
        VN2CN5_sign => VN_sign_out(2849),
        codeword => codeword(474),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN475 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2855 downto 2850),
        Din0 => VN475_in0,
        Din1 => VN475_in1,
        Din2 => VN475_in2,
        Din3 => VN475_in3,
        Din4 => VN475_in4,
        Din5 => VN475_in5,
        VN2CN0_bit => VN_data_out(2850),
        VN2CN1_bit => VN_data_out(2851),
        VN2CN2_bit => VN_data_out(2852),
        VN2CN3_bit => VN_data_out(2853),
        VN2CN4_bit => VN_data_out(2854),
        VN2CN5_bit => VN_data_out(2855),
        VN2CN0_sign => VN_sign_out(2850),
        VN2CN1_sign => VN_sign_out(2851),
        VN2CN2_sign => VN_sign_out(2852),
        VN2CN3_sign => VN_sign_out(2853),
        VN2CN4_sign => VN_sign_out(2854),
        VN2CN5_sign => VN_sign_out(2855),
        codeword => codeword(475),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN476 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2861 downto 2856),
        Din0 => VN476_in0,
        Din1 => VN476_in1,
        Din2 => VN476_in2,
        Din3 => VN476_in3,
        Din4 => VN476_in4,
        Din5 => VN476_in5,
        VN2CN0_bit => VN_data_out(2856),
        VN2CN1_bit => VN_data_out(2857),
        VN2CN2_bit => VN_data_out(2858),
        VN2CN3_bit => VN_data_out(2859),
        VN2CN4_bit => VN_data_out(2860),
        VN2CN5_bit => VN_data_out(2861),
        VN2CN0_sign => VN_sign_out(2856),
        VN2CN1_sign => VN_sign_out(2857),
        VN2CN2_sign => VN_sign_out(2858),
        VN2CN3_sign => VN_sign_out(2859),
        VN2CN4_sign => VN_sign_out(2860),
        VN2CN5_sign => VN_sign_out(2861),
        codeword => codeword(476),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN477 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2867 downto 2862),
        Din0 => VN477_in0,
        Din1 => VN477_in1,
        Din2 => VN477_in2,
        Din3 => VN477_in3,
        Din4 => VN477_in4,
        Din5 => VN477_in5,
        VN2CN0_bit => VN_data_out(2862),
        VN2CN1_bit => VN_data_out(2863),
        VN2CN2_bit => VN_data_out(2864),
        VN2CN3_bit => VN_data_out(2865),
        VN2CN4_bit => VN_data_out(2866),
        VN2CN5_bit => VN_data_out(2867),
        VN2CN0_sign => VN_sign_out(2862),
        VN2CN1_sign => VN_sign_out(2863),
        VN2CN2_sign => VN_sign_out(2864),
        VN2CN3_sign => VN_sign_out(2865),
        VN2CN4_sign => VN_sign_out(2866),
        VN2CN5_sign => VN_sign_out(2867),
        codeword => codeword(477),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN478 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2873 downto 2868),
        Din0 => VN478_in0,
        Din1 => VN478_in1,
        Din2 => VN478_in2,
        Din3 => VN478_in3,
        Din4 => VN478_in4,
        Din5 => VN478_in5,
        VN2CN0_bit => VN_data_out(2868),
        VN2CN1_bit => VN_data_out(2869),
        VN2CN2_bit => VN_data_out(2870),
        VN2CN3_bit => VN_data_out(2871),
        VN2CN4_bit => VN_data_out(2872),
        VN2CN5_bit => VN_data_out(2873),
        VN2CN0_sign => VN_sign_out(2868),
        VN2CN1_sign => VN_sign_out(2869),
        VN2CN2_sign => VN_sign_out(2870),
        VN2CN3_sign => VN_sign_out(2871),
        VN2CN4_sign => VN_sign_out(2872),
        VN2CN5_sign => VN_sign_out(2873),
        codeword => codeword(478),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN479 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2879 downto 2874),
        Din0 => VN479_in0,
        Din1 => VN479_in1,
        Din2 => VN479_in2,
        Din3 => VN479_in3,
        Din4 => VN479_in4,
        Din5 => VN479_in5,
        VN2CN0_bit => VN_data_out(2874),
        VN2CN1_bit => VN_data_out(2875),
        VN2CN2_bit => VN_data_out(2876),
        VN2CN3_bit => VN_data_out(2877),
        VN2CN4_bit => VN_data_out(2878),
        VN2CN5_bit => VN_data_out(2879),
        VN2CN0_sign => VN_sign_out(2874),
        VN2CN1_sign => VN_sign_out(2875),
        VN2CN2_sign => VN_sign_out(2876),
        VN2CN3_sign => VN_sign_out(2877),
        VN2CN4_sign => VN_sign_out(2878),
        VN2CN5_sign => VN_sign_out(2879),
        codeword => codeword(479),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN480 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2885 downto 2880),
        Din0 => VN480_in0,
        Din1 => VN480_in1,
        Din2 => VN480_in2,
        Din3 => VN480_in3,
        Din4 => VN480_in4,
        Din5 => VN480_in5,
        VN2CN0_bit => VN_data_out(2880),
        VN2CN1_bit => VN_data_out(2881),
        VN2CN2_bit => VN_data_out(2882),
        VN2CN3_bit => VN_data_out(2883),
        VN2CN4_bit => VN_data_out(2884),
        VN2CN5_bit => VN_data_out(2885),
        VN2CN0_sign => VN_sign_out(2880),
        VN2CN1_sign => VN_sign_out(2881),
        VN2CN2_sign => VN_sign_out(2882),
        VN2CN3_sign => VN_sign_out(2883),
        VN2CN4_sign => VN_sign_out(2884),
        VN2CN5_sign => VN_sign_out(2885),
        codeword => codeword(480),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN481 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2891 downto 2886),
        Din0 => VN481_in0,
        Din1 => VN481_in1,
        Din2 => VN481_in2,
        Din3 => VN481_in3,
        Din4 => VN481_in4,
        Din5 => VN481_in5,
        VN2CN0_bit => VN_data_out(2886),
        VN2CN1_bit => VN_data_out(2887),
        VN2CN2_bit => VN_data_out(2888),
        VN2CN3_bit => VN_data_out(2889),
        VN2CN4_bit => VN_data_out(2890),
        VN2CN5_bit => VN_data_out(2891),
        VN2CN0_sign => VN_sign_out(2886),
        VN2CN1_sign => VN_sign_out(2887),
        VN2CN2_sign => VN_sign_out(2888),
        VN2CN3_sign => VN_sign_out(2889),
        VN2CN4_sign => VN_sign_out(2890),
        VN2CN5_sign => VN_sign_out(2891),
        codeword => codeword(481),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN482 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2897 downto 2892),
        Din0 => VN482_in0,
        Din1 => VN482_in1,
        Din2 => VN482_in2,
        Din3 => VN482_in3,
        Din4 => VN482_in4,
        Din5 => VN482_in5,
        VN2CN0_bit => VN_data_out(2892),
        VN2CN1_bit => VN_data_out(2893),
        VN2CN2_bit => VN_data_out(2894),
        VN2CN3_bit => VN_data_out(2895),
        VN2CN4_bit => VN_data_out(2896),
        VN2CN5_bit => VN_data_out(2897),
        VN2CN0_sign => VN_sign_out(2892),
        VN2CN1_sign => VN_sign_out(2893),
        VN2CN2_sign => VN_sign_out(2894),
        VN2CN3_sign => VN_sign_out(2895),
        VN2CN4_sign => VN_sign_out(2896),
        VN2CN5_sign => VN_sign_out(2897),
        codeword => codeword(482),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN483 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2903 downto 2898),
        Din0 => VN483_in0,
        Din1 => VN483_in1,
        Din2 => VN483_in2,
        Din3 => VN483_in3,
        Din4 => VN483_in4,
        Din5 => VN483_in5,
        VN2CN0_bit => VN_data_out(2898),
        VN2CN1_bit => VN_data_out(2899),
        VN2CN2_bit => VN_data_out(2900),
        VN2CN3_bit => VN_data_out(2901),
        VN2CN4_bit => VN_data_out(2902),
        VN2CN5_bit => VN_data_out(2903),
        VN2CN0_sign => VN_sign_out(2898),
        VN2CN1_sign => VN_sign_out(2899),
        VN2CN2_sign => VN_sign_out(2900),
        VN2CN3_sign => VN_sign_out(2901),
        VN2CN4_sign => VN_sign_out(2902),
        VN2CN5_sign => VN_sign_out(2903),
        codeword => codeword(483),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN484 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2909 downto 2904),
        Din0 => VN484_in0,
        Din1 => VN484_in1,
        Din2 => VN484_in2,
        Din3 => VN484_in3,
        Din4 => VN484_in4,
        Din5 => VN484_in5,
        VN2CN0_bit => VN_data_out(2904),
        VN2CN1_bit => VN_data_out(2905),
        VN2CN2_bit => VN_data_out(2906),
        VN2CN3_bit => VN_data_out(2907),
        VN2CN4_bit => VN_data_out(2908),
        VN2CN5_bit => VN_data_out(2909),
        VN2CN0_sign => VN_sign_out(2904),
        VN2CN1_sign => VN_sign_out(2905),
        VN2CN2_sign => VN_sign_out(2906),
        VN2CN3_sign => VN_sign_out(2907),
        VN2CN4_sign => VN_sign_out(2908),
        VN2CN5_sign => VN_sign_out(2909),
        codeword => codeword(484),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN485 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2915 downto 2910),
        Din0 => VN485_in0,
        Din1 => VN485_in1,
        Din2 => VN485_in2,
        Din3 => VN485_in3,
        Din4 => VN485_in4,
        Din5 => VN485_in5,
        VN2CN0_bit => VN_data_out(2910),
        VN2CN1_bit => VN_data_out(2911),
        VN2CN2_bit => VN_data_out(2912),
        VN2CN3_bit => VN_data_out(2913),
        VN2CN4_bit => VN_data_out(2914),
        VN2CN5_bit => VN_data_out(2915),
        VN2CN0_sign => VN_sign_out(2910),
        VN2CN1_sign => VN_sign_out(2911),
        VN2CN2_sign => VN_sign_out(2912),
        VN2CN3_sign => VN_sign_out(2913),
        VN2CN4_sign => VN_sign_out(2914),
        VN2CN5_sign => VN_sign_out(2915),
        codeword => codeword(485),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN486 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2921 downto 2916),
        Din0 => VN486_in0,
        Din1 => VN486_in1,
        Din2 => VN486_in2,
        Din3 => VN486_in3,
        Din4 => VN486_in4,
        Din5 => VN486_in5,
        VN2CN0_bit => VN_data_out(2916),
        VN2CN1_bit => VN_data_out(2917),
        VN2CN2_bit => VN_data_out(2918),
        VN2CN3_bit => VN_data_out(2919),
        VN2CN4_bit => VN_data_out(2920),
        VN2CN5_bit => VN_data_out(2921),
        VN2CN0_sign => VN_sign_out(2916),
        VN2CN1_sign => VN_sign_out(2917),
        VN2CN2_sign => VN_sign_out(2918),
        VN2CN3_sign => VN_sign_out(2919),
        VN2CN4_sign => VN_sign_out(2920),
        VN2CN5_sign => VN_sign_out(2921),
        codeword => codeword(486),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN487 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2927 downto 2922),
        Din0 => VN487_in0,
        Din1 => VN487_in1,
        Din2 => VN487_in2,
        Din3 => VN487_in3,
        Din4 => VN487_in4,
        Din5 => VN487_in5,
        VN2CN0_bit => VN_data_out(2922),
        VN2CN1_bit => VN_data_out(2923),
        VN2CN2_bit => VN_data_out(2924),
        VN2CN3_bit => VN_data_out(2925),
        VN2CN4_bit => VN_data_out(2926),
        VN2CN5_bit => VN_data_out(2927),
        VN2CN0_sign => VN_sign_out(2922),
        VN2CN1_sign => VN_sign_out(2923),
        VN2CN2_sign => VN_sign_out(2924),
        VN2CN3_sign => VN_sign_out(2925),
        VN2CN4_sign => VN_sign_out(2926),
        VN2CN5_sign => VN_sign_out(2927),
        codeword => codeword(487),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN488 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2933 downto 2928),
        Din0 => VN488_in0,
        Din1 => VN488_in1,
        Din2 => VN488_in2,
        Din3 => VN488_in3,
        Din4 => VN488_in4,
        Din5 => VN488_in5,
        VN2CN0_bit => VN_data_out(2928),
        VN2CN1_bit => VN_data_out(2929),
        VN2CN2_bit => VN_data_out(2930),
        VN2CN3_bit => VN_data_out(2931),
        VN2CN4_bit => VN_data_out(2932),
        VN2CN5_bit => VN_data_out(2933),
        VN2CN0_sign => VN_sign_out(2928),
        VN2CN1_sign => VN_sign_out(2929),
        VN2CN2_sign => VN_sign_out(2930),
        VN2CN3_sign => VN_sign_out(2931),
        VN2CN4_sign => VN_sign_out(2932),
        VN2CN5_sign => VN_sign_out(2933),
        codeword => codeword(488),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN489 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2939 downto 2934),
        Din0 => VN489_in0,
        Din1 => VN489_in1,
        Din2 => VN489_in2,
        Din3 => VN489_in3,
        Din4 => VN489_in4,
        Din5 => VN489_in5,
        VN2CN0_bit => VN_data_out(2934),
        VN2CN1_bit => VN_data_out(2935),
        VN2CN2_bit => VN_data_out(2936),
        VN2CN3_bit => VN_data_out(2937),
        VN2CN4_bit => VN_data_out(2938),
        VN2CN5_bit => VN_data_out(2939),
        VN2CN0_sign => VN_sign_out(2934),
        VN2CN1_sign => VN_sign_out(2935),
        VN2CN2_sign => VN_sign_out(2936),
        VN2CN3_sign => VN_sign_out(2937),
        VN2CN4_sign => VN_sign_out(2938),
        VN2CN5_sign => VN_sign_out(2939),
        codeword => codeword(489),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN490 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2945 downto 2940),
        Din0 => VN490_in0,
        Din1 => VN490_in1,
        Din2 => VN490_in2,
        Din3 => VN490_in3,
        Din4 => VN490_in4,
        Din5 => VN490_in5,
        VN2CN0_bit => VN_data_out(2940),
        VN2CN1_bit => VN_data_out(2941),
        VN2CN2_bit => VN_data_out(2942),
        VN2CN3_bit => VN_data_out(2943),
        VN2CN4_bit => VN_data_out(2944),
        VN2CN5_bit => VN_data_out(2945),
        VN2CN0_sign => VN_sign_out(2940),
        VN2CN1_sign => VN_sign_out(2941),
        VN2CN2_sign => VN_sign_out(2942),
        VN2CN3_sign => VN_sign_out(2943),
        VN2CN4_sign => VN_sign_out(2944),
        VN2CN5_sign => VN_sign_out(2945),
        codeword => codeword(490),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN491 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2951 downto 2946),
        Din0 => VN491_in0,
        Din1 => VN491_in1,
        Din2 => VN491_in2,
        Din3 => VN491_in3,
        Din4 => VN491_in4,
        Din5 => VN491_in5,
        VN2CN0_bit => VN_data_out(2946),
        VN2CN1_bit => VN_data_out(2947),
        VN2CN2_bit => VN_data_out(2948),
        VN2CN3_bit => VN_data_out(2949),
        VN2CN4_bit => VN_data_out(2950),
        VN2CN5_bit => VN_data_out(2951),
        VN2CN0_sign => VN_sign_out(2946),
        VN2CN1_sign => VN_sign_out(2947),
        VN2CN2_sign => VN_sign_out(2948),
        VN2CN3_sign => VN_sign_out(2949),
        VN2CN4_sign => VN_sign_out(2950),
        VN2CN5_sign => VN_sign_out(2951),
        codeword => codeword(491),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN492 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2957 downto 2952),
        Din0 => VN492_in0,
        Din1 => VN492_in1,
        Din2 => VN492_in2,
        Din3 => VN492_in3,
        Din4 => VN492_in4,
        Din5 => VN492_in5,
        VN2CN0_bit => VN_data_out(2952),
        VN2CN1_bit => VN_data_out(2953),
        VN2CN2_bit => VN_data_out(2954),
        VN2CN3_bit => VN_data_out(2955),
        VN2CN4_bit => VN_data_out(2956),
        VN2CN5_bit => VN_data_out(2957),
        VN2CN0_sign => VN_sign_out(2952),
        VN2CN1_sign => VN_sign_out(2953),
        VN2CN2_sign => VN_sign_out(2954),
        VN2CN3_sign => VN_sign_out(2955),
        VN2CN4_sign => VN_sign_out(2956),
        VN2CN5_sign => VN_sign_out(2957),
        codeword => codeword(492),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN493 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2963 downto 2958),
        Din0 => VN493_in0,
        Din1 => VN493_in1,
        Din2 => VN493_in2,
        Din3 => VN493_in3,
        Din4 => VN493_in4,
        Din5 => VN493_in5,
        VN2CN0_bit => VN_data_out(2958),
        VN2CN1_bit => VN_data_out(2959),
        VN2CN2_bit => VN_data_out(2960),
        VN2CN3_bit => VN_data_out(2961),
        VN2CN4_bit => VN_data_out(2962),
        VN2CN5_bit => VN_data_out(2963),
        VN2CN0_sign => VN_sign_out(2958),
        VN2CN1_sign => VN_sign_out(2959),
        VN2CN2_sign => VN_sign_out(2960),
        VN2CN3_sign => VN_sign_out(2961),
        VN2CN4_sign => VN_sign_out(2962),
        VN2CN5_sign => VN_sign_out(2963),
        codeword => codeword(493),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN494 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2969 downto 2964),
        Din0 => VN494_in0,
        Din1 => VN494_in1,
        Din2 => VN494_in2,
        Din3 => VN494_in3,
        Din4 => VN494_in4,
        Din5 => VN494_in5,
        VN2CN0_bit => VN_data_out(2964),
        VN2CN1_bit => VN_data_out(2965),
        VN2CN2_bit => VN_data_out(2966),
        VN2CN3_bit => VN_data_out(2967),
        VN2CN4_bit => VN_data_out(2968),
        VN2CN5_bit => VN_data_out(2969),
        VN2CN0_sign => VN_sign_out(2964),
        VN2CN1_sign => VN_sign_out(2965),
        VN2CN2_sign => VN_sign_out(2966),
        VN2CN3_sign => VN_sign_out(2967),
        VN2CN4_sign => VN_sign_out(2968),
        VN2CN5_sign => VN_sign_out(2969),
        codeword => codeword(494),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN495 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2975 downto 2970),
        Din0 => VN495_in0,
        Din1 => VN495_in1,
        Din2 => VN495_in2,
        Din3 => VN495_in3,
        Din4 => VN495_in4,
        Din5 => VN495_in5,
        VN2CN0_bit => VN_data_out(2970),
        VN2CN1_bit => VN_data_out(2971),
        VN2CN2_bit => VN_data_out(2972),
        VN2CN3_bit => VN_data_out(2973),
        VN2CN4_bit => VN_data_out(2974),
        VN2CN5_bit => VN_data_out(2975),
        VN2CN0_sign => VN_sign_out(2970),
        VN2CN1_sign => VN_sign_out(2971),
        VN2CN2_sign => VN_sign_out(2972),
        VN2CN3_sign => VN_sign_out(2973),
        VN2CN4_sign => VN_sign_out(2974),
        VN2CN5_sign => VN_sign_out(2975),
        codeword => codeword(495),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN496 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2981 downto 2976),
        Din0 => VN496_in0,
        Din1 => VN496_in1,
        Din2 => VN496_in2,
        Din3 => VN496_in3,
        Din4 => VN496_in4,
        Din5 => VN496_in5,
        VN2CN0_bit => VN_data_out(2976),
        VN2CN1_bit => VN_data_out(2977),
        VN2CN2_bit => VN_data_out(2978),
        VN2CN3_bit => VN_data_out(2979),
        VN2CN4_bit => VN_data_out(2980),
        VN2CN5_bit => VN_data_out(2981),
        VN2CN0_sign => VN_sign_out(2976),
        VN2CN1_sign => VN_sign_out(2977),
        VN2CN2_sign => VN_sign_out(2978),
        VN2CN3_sign => VN_sign_out(2979),
        VN2CN4_sign => VN_sign_out(2980),
        VN2CN5_sign => VN_sign_out(2981),
        codeword => codeword(496),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN497 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2987 downto 2982),
        Din0 => VN497_in0,
        Din1 => VN497_in1,
        Din2 => VN497_in2,
        Din3 => VN497_in3,
        Din4 => VN497_in4,
        Din5 => VN497_in5,
        VN2CN0_bit => VN_data_out(2982),
        VN2CN1_bit => VN_data_out(2983),
        VN2CN2_bit => VN_data_out(2984),
        VN2CN3_bit => VN_data_out(2985),
        VN2CN4_bit => VN_data_out(2986),
        VN2CN5_bit => VN_data_out(2987),
        VN2CN0_sign => VN_sign_out(2982),
        VN2CN1_sign => VN_sign_out(2983),
        VN2CN2_sign => VN_sign_out(2984),
        VN2CN3_sign => VN_sign_out(2985),
        VN2CN4_sign => VN_sign_out(2986),
        VN2CN5_sign => VN_sign_out(2987),
        codeword => codeword(497),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN498 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2993 downto 2988),
        Din0 => VN498_in0,
        Din1 => VN498_in1,
        Din2 => VN498_in2,
        Din3 => VN498_in3,
        Din4 => VN498_in4,
        Din5 => VN498_in5,
        VN2CN0_bit => VN_data_out(2988),
        VN2CN1_bit => VN_data_out(2989),
        VN2CN2_bit => VN_data_out(2990),
        VN2CN3_bit => VN_data_out(2991),
        VN2CN4_bit => VN_data_out(2992),
        VN2CN5_bit => VN_data_out(2993),
        VN2CN0_sign => VN_sign_out(2988),
        VN2CN1_sign => VN_sign_out(2989),
        VN2CN2_sign => VN_sign_out(2990),
        VN2CN3_sign => VN_sign_out(2991),
        VN2CN4_sign => VN_sign_out(2992),
        VN2CN5_sign => VN_sign_out(2993),
        codeword => codeword(498),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN499 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(2999 downto 2994),
        Din0 => VN499_in0,
        Din1 => VN499_in1,
        Din2 => VN499_in2,
        Din3 => VN499_in3,
        Din4 => VN499_in4,
        Din5 => VN499_in5,
        VN2CN0_bit => VN_data_out(2994),
        VN2CN1_bit => VN_data_out(2995),
        VN2CN2_bit => VN_data_out(2996),
        VN2CN3_bit => VN_data_out(2997),
        VN2CN4_bit => VN_data_out(2998),
        VN2CN5_bit => VN_data_out(2999),
        VN2CN0_sign => VN_sign_out(2994),
        VN2CN1_sign => VN_sign_out(2995),
        VN2CN2_sign => VN_sign_out(2996),
        VN2CN3_sign => VN_sign_out(2997),
        VN2CN4_sign => VN_sign_out(2998),
        VN2CN5_sign => VN_sign_out(2999),
        codeword => codeword(499),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN500 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3005 downto 3000),
        Din0 => VN500_in0,
        Din1 => VN500_in1,
        Din2 => VN500_in2,
        Din3 => VN500_in3,
        Din4 => VN500_in4,
        Din5 => VN500_in5,
        VN2CN0_bit => VN_data_out(3000),
        VN2CN1_bit => VN_data_out(3001),
        VN2CN2_bit => VN_data_out(3002),
        VN2CN3_bit => VN_data_out(3003),
        VN2CN4_bit => VN_data_out(3004),
        VN2CN5_bit => VN_data_out(3005),
        VN2CN0_sign => VN_sign_out(3000),
        VN2CN1_sign => VN_sign_out(3001),
        VN2CN2_sign => VN_sign_out(3002),
        VN2CN3_sign => VN_sign_out(3003),
        VN2CN4_sign => VN_sign_out(3004),
        VN2CN5_sign => VN_sign_out(3005),
        codeword => codeword(500),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN501 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3011 downto 3006),
        Din0 => VN501_in0,
        Din1 => VN501_in1,
        Din2 => VN501_in2,
        Din3 => VN501_in3,
        Din4 => VN501_in4,
        Din5 => VN501_in5,
        VN2CN0_bit => VN_data_out(3006),
        VN2CN1_bit => VN_data_out(3007),
        VN2CN2_bit => VN_data_out(3008),
        VN2CN3_bit => VN_data_out(3009),
        VN2CN4_bit => VN_data_out(3010),
        VN2CN5_bit => VN_data_out(3011),
        VN2CN0_sign => VN_sign_out(3006),
        VN2CN1_sign => VN_sign_out(3007),
        VN2CN2_sign => VN_sign_out(3008),
        VN2CN3_sign => VN_sign_out(3009),
        VN2CN4_sign => VN_sign_out(3010),
        VN2CN5_sign => VN_sign_out(3011),
        codeword => codeword(501),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN502 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3017 downto 3012),
        Din0 => VN502_in0,
        Din1 => VN502_in1,
        Din2 => VN502_in2,
        Din3 => VN502_in3,
        Din4 => VN502_in4,
        Din5 => VN502_in5,
        VN2CN0_bit => VN_data_out(3012),
        VN2CN1_bit => VN_data_out(3013),
        VN2CN2_bit => VN_data_out(3014),
        VN2CN3_bit => VN_data_out(3015),
        VN2CN4_bit => VN_data_out(3016),
        VN2CN5_bit => VN_data_out(3017),
        VN2CN0_sign => VN_sign_out(3012),
        VN2CN1_sign => VN_sign_out(3013),
        VN2CN2_sign => VN_sign_out(3014),
        VN2CN3_sign => VN_sign_out(3015),
        VN2CN4_sign => VN_sign_out(3016),
        VN2CN5_sign => VN_sign_out(3017),
        codeword => codeword(502),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN503 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3023 downto 3018),
        Din0 => VN503_in0,
        Din1 => VN503_in1,
        Din2 => VN503_in2,
        Din3 => VN503_in3,
        Din4 => VN503_in4,
        Din5 => VN503_in5,
        VN2CN0_bit => VN_data_out(3018),
        VN2CN1_bit => VN_data_out(3019),
        VN2CN2_bit => VN_data_out(3020),
        VN2CN3_bit => VN_data_out(3021),
        VN2CN4_bit => VN_data_out(3022),
        VN2CN5_bit => VN_data_out(3023),
        VN2CN0_sign => VN_sign_out(3018),
        VN2CN1_sign => VN_sign_out(3019),
        VN2CN2_sign => VN_sign_out(3020),
        VN2CN3_sign => VN_sign_out(3021),
        VN2CN4_sign => VN_sign_out(3022),
        VN2CN5_sign => VN_sign_out(3023),
        codeword => codeword(503),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN504 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3029 downto 3024),
        Din0 => VN504_in0,
        Din1 => VN504_in1,
        Din2 => VN504_in2,
        Din3 => VN504_in3,
        Din4 => VN504_in4,
        Din5 => VN504_in5,
        VN2CN0_bit => VN_data_out(3024),
        VN2CN1_bit => VN_data_out(3025),
        VN2CN2_bit => VN_data_out(3026),
        VN2CN3_bit => VN_data_out(3027),
        VN2CN4_bit => VN_data_out(3028),
        VN2CN5_bit => VN_data_out(3029),
        VN2CN0_sign => VN_sign_out(3024),
        VN2CN1_sign => VN_sign_out(3025),
        VN2CN2_sign => VN_sign_out(3026),
        VN2CN3_sign => VN_sign_out(3027),
        VN2CN4_sign => VN_sign_out(3028),
        VN2CN5_sign => VN_sign_out(3029),
        codeword => codeword(504),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN505 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3035 downto 3030),
        Din0 => VN505_in0,
        Din1 => VN505_in1,
        Din2 => VN505_in2,
        Din3 => VN505_in3,
        Din4 => VN505_in4,
        Din5 => VN505_in5,
        VN2CN0_bit => VN_data_out(3030),
        VN2CN1_bit => VN_data_out(3031),
        VN2CN2_bit => VN_data_out(3032),
        VN2CN3_bit => VN_data_out(3033),
        VN2CN4_bit => VN_data_out(3034),
        VN2CN5_bit => VN_data_out(3035),
        VN2CN0_sign => VN_sign_out(3030),
        VN2CN1_sign => VN_sign_out(3031),
        VN2CN2_sign => VN_sign_out(3032),
        VN2CN3_sign => VN_sign_out(3033),
        VN2CN4_sign => VN_sign_out(3034),
        VN2CN5_sign => VN_sign_out(3035),
        codeword => codeword(505),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN506 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3041 downto 3036),
        Din0 => VN506_in0,
        Din1 => VN506_in1,
        Din2 => VN506_in2,
        Din3 => VN506_in3,
        Din4 => VN506_in4,
        Din5 => VN506_in5,
        VN2CN0_bit => VN_data_out(3036),
        VN2CN1_bit => VN_data_out(3037),
        VN2CN2_bit => VN_data_out(3038),
        VN2CN3_bit => VN_data_out(3039),
        VN2CN4_bit => VN_data_out(3040),
        VN2CN5_bit => VN_data_out(3041),
        VN2CN0_sign => VN_sign_out(3036),
        VN2CN1_sign => VN_sign_out(3037),
        VN2CN2_sign => VN_sign_out(3038),
        VN2CN3_sign => VN_sign_out(3039),
        VN2CN4_sign => VN_sign_out(3040),
        VN2CN5_sign => VN_sign_out(3041),
        codeword => codeword(506),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN507 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3047 downto 3042),
        Din0 => VN507_in0,
        Din1 => VN507_in1,
        Din2 => VN507_in2,
        Din3 => VN507_in3,
        Din4 => VN507_in4,
        Din5 => VN507_in5,
        VN2CN0_bit => VN_data_out(3042),
        VN2CN1_bit => VN_data_out(3043),
        VN2CN2_bit => VN_data_out(3044),
        VN2CN3_bit => VN_data_out(3045),
        VN2CN4_bit => VN_data_out(3046),
        VN2CN5_bit => VN_data_out(3047),
        VN2CN0_sign => VN_sign_out(3042),
        VN2CN1_sign => VN_sign_out(3043),
        VN2CN2_sign => VN_sign_out(3044),
        VN2CN3_sign => VN_sign_out(3045),
        VN2CN4_sign => VN_sign_out(3046),
        VN2CN5_sign => VN_sign_out(3047),
        codeword => codeword(507),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN508 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3053 downto 3048),
        Din0 => VN508_in0,
        Din1 => VN508_in1,
        Din2 => VN508_in2,
        Din3 => VN508_in3,
        Din4 => VN508_in4,
        Din5 => VN508_in5,
        VN2CN0_bit => VN_data_out(3048),
        VN2CN1_bit => VN_data_out(3049),
        VN2CN2_bit => VN_data_out(3050),
        VN2CN3_bit => VN_data_out(3051),
        VN2CN4_bit => VN_data_out(3052),
        VN2CN5_bit => VN_data_out(3053),
        VN2CN0_sign => VN_sign_out(3048),
        VN2CN1_sign => VN_sign_out(3049),
        VN2CN2_sign => VN_sign_out(3050),
        VN2CN3_sign => VN_sign_out(3051),
        VN2CN4_sign => VN_sign_out(3052),
        VN2CN5_sign => VN_sign_out(3053),
        codeword => codeword(508),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN509 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3059 downto 3054),
        Din0 => VN509_in0,
        Din1 => VN509_in1,
        Din2 => VN509_in2,
        Din3 => VN509_in3,
        Din4 => VN509_in4,
        Din5 => VN509_in5,
        VN2CN0_bit => VN_data_out(3054),
        VN2CN1_bit => VN_data_out(3055),
        VN2CN2_bit => VN_data_out(3056),
        VN2CN3_bit => VN_data_out(3057),
        VN2CN4_bit => VN_data_out(3058),
        VN2CN5_bit => VN_data_out(3059),
        VN2CN0_sign => VN_sign_out(3054),
        VN2CN1_sign => VN_sign_out(3055),
        VN2CN2_sign => VN_sign_out(3056),
        VN2CN3_sign => VN_sign_out(3057),
        VN2CN4_sign => VN_sign_out(3058),
        VN2CN5_sign => VN_sign_out(3059),
        codeword => codeword(509),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN510 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3065 downto 3060),
        Din0 => VN510_in0,
        Din1 => VN510_in1,
        Din2 => VN510_in2,
        Din3 => VN510_in3,
        Din4 => VN510_in4,
        Din5 => VN510_in5,
        VN2CN0_bit => VN_data_out(3060),
        VN2CN1_bit => VN_data_out(3061),
        VN2CN2_bit => VN_data_out(3062),
        VN2CN3_bit => VN_data_out(3063),
        VN2CN4_bit => VN_data_out(3064),
        VN2CN5_bit => VN_data_out(3065),
        VN2CN0_sign => VN_sign_out(3060),
        VN2CN1_sign => VN_sign_out(3061),
        VN2CN2_sign => VN_sign_out(3062),
        VN2CN3_sign => VN_sign_out(3063),
        VN2CN4_sign => VN_sign_out(3064),
        VN2CN5_sign => VN_sign_out(3065),
        codeword => codeword(510),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN511 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3071 downto 3066),
        Din0 => VN511_in0,
        Din1 => VN511_in1,
        Din2 => VN511_in2,
        Din3 => VN511_in3,
        Din4 => VN511_in4,
        Din5 => VN511_in5,
        VN2CN0_bit => VN_data_out(3066),
        VN2CN1_bit => VN_data_out(3067),
        VN2CN2_bit => VN_data_out(3068),
        VN2CN3_bit => VN_data_out(3069),
        VN2CN4_bit => VN_data_out(3070),
        VN2CN5_bit => VN_data_out(3071),
        VN2CN0_sign => VN_sign_out(3066),
        VN2CN1_sign => VN_sign_out(3067),
        VN2CN2_sign => VN_sign_out(3068),
        VN2CN3_sign => VN_sign_out(3069),
        VN2CN4_sign => VN_sign_out(3070),
        VN2CN5_sign => VN_sign_out(3071),
        codeword => codeword(511),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN512 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3077 downto 3072),
        Din0 => VN512_in0,
        Din1 => VN512_in1,
        Din2 => VN512_in2,
        Din3 => VN512_in3,
        Din4 => VN512_in4,
        Din5 => VN512_in5,
        VN2CN0_bit => VN_data_out(3072),
        VN2CN1_bit => VN_data_out(3073),
        VN2CN2_bit => VN_data_out(3074),
        VN2CN3_bit => VN_data_out(3075),
        VN2CN4_bit => VN_data_out(3076),
        VN2CN5_bit => VN_data_out(3077),
        VN2CN0_sign => VN_sign_out(3072),
        VN2CN1_sign => VN_sign_out(3073),
        VN2CN2_sign => VN_sign_out(3074),
        VN2CN3_sign => VN_sign_out(3075),
        VN2CN4_sign => VN_sign_out(3076),
        VN2CN5_sign => VN_sign_out(3077),
        codeword => codeword(512),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN513 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3083 downto 3078),
        Din0 => VN513_in0,
        Din1 => VN513_in1,
        Din2 => VN513_in2,
        Din3 => VN513_in3,
        Din4 => VN513_in4,
        Din5 => VN513_in5,
        VN2CN0_bit => VN_data_out(3078),
        VN2CN1_bit => VN_data_out(3079),
        VN2CN2_bit => VN_data_out(3080),
        VN2CN3_bit => VN_data_out(3081),
        VN2CN4_bit => VN_data_out(3082),
        VN2CN5_bit => VN_data_out(3083),
        VN2CN0_sign => VN_sign_out(3078),
        VN2CN1_sign => VN_sign_out(3079),
        VN2CN2_sign => VN_sign_out(3080),
        VN2CN3_sign => VN_sign_out(3081),
        VN2CN4_sign => VN_sign_out(3082),
        VN2CN5_sign => VN_sign_out(3083),
        codeword => codeword(513),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN514 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3089 downto 3084),
        Din0 => VN514_in0,
        Din1 => VN514_in1,
        Din2 => VN514_in2,
        Din3 => VN514_in3,
        Din4 => VN514_in4,
        Din5 => VN514_in5,
        VN2CN0_bit => VN_data_out(3084),
        VN2CN1_bit => VN_data_out(3085),
        VN2CN2_bit => VN_data_out(3086),
        VN2CN3_bit => VN_data_out(3087),
        VN2CN4_bit => VN_data_out(3088),
        VN2CN5_bit => VN_data_out(3089),
        VN2CN0_sign => VN_sign_out(3084),
        VN2CN1_sign => VN_sign_out(3085),
        VN2CN2_sign => VN_sign_out(3086),
        VN2CN3_sign => VN_sign_out(3087),
        VN2CN4_sign => VN_sign_out(3088),
        VN2CN5_sign => VN_sign_out(3089),
        codeword => codeword(514),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN515 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3095 downto 3090),
        Din0 => VN515_in0,
        Din1 => VN515_in1,
        Din2 => VN515_in2,
        Din3 => VN515_in3,
        Din4 => VN515_in4,
        Din5 => VN515_in5,
        VN2CN0_bit => VN_data_out(3090),
        VN2CN1_bit => VN_data_out(3091),
        VN2CN2_bit => VN_data_out(3092),
        VN2CN3_bit => VN_data_out(3093),
        VN2CN4_bit => VN_data_out(3094),
        VN2CN5_bit => VN_data_out(3095),
        VN2CN0_sign => VN_sign_out(3090),
        VN2CN1_sign => VN_sign_out(3091),
        VN2CN2_sign => VN_sign_out(3092),
        VN2CN3_sign => VN_sign_out(3093),
        VN2CN4_sign => VN_sign_out(3094),
        VN2CN5_sign => VN_sign_out(3095),
        codeword => codeword(515),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN516 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3101 downto 3096),
        Din0 => VN516_in0,
        Din1 => VN516_in1,
        Din2 => VN516_in2,
        Din3 => VN516_in3,
        Din4 => VN516_in4,
        Din5 => VN516_in5,
        VN2CN0_bit => VN_data_out(3096),
        VN2CN1_bit => VN_data_out(3097),
        VN2CN2_bit => VN_data_out(3098),
        VN2CN3_bit => VN_data_out(3099),
        VN2CN4_bit => VN_data_out(3100),
        VN2CN5_bit => VN_data_out(3101),
        VN2CN0_sign => VN_sign_out(3096),
        VN2CN1_sign => VN_sign_out(3097),
        VN2CN2_sign => VN_sign_out(3098),
        VN2CN3_sign => VN_sign_out(3099),
        VN2CN4_sign => VN_sign_out(3100),
        VN2CN5_sign => VN_sign_out(3101),
        codeword => codeword(516),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN517 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3107 downto 3102),
        Din0 => VN517_in0,
        Din1 => VN517_in1,
        Din2 => VN517_in2,
        Din3 => VN517_in3,
        Din4 => VN517_in4,
        Din5 => VN517_in5,
        VN2CN0_bit => VN_data_out(3102),
        VN2CN1_bit => VN_data_out(3103),
        VN2CN2_bit => VN_data_out(3104),
        VN2CN3_bit => VN_data_out(3105),
        VN2CN4_bit => VN_data_out(3106),
        VN2CN5_bit => VN_data_out(3107),
        VN2CN0_sign => VN_sign_out(3102),
        VN2CN1_sign => VN_sign_out(3103),
        VN2CN2_sign => VN_sign_out(3104),
        VN2CN3_sign => VN_sign_out(3105),
        VN2CN4_sign => VN_sign_out(3106),
        VN2CN5_sign => VN_sign_out(3107),
        codeword => codeword(517),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN518 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3113 downto 3108),
        Din0 => VN518_in0,
        Din1 => VN518_in1,
        Din2 => VN518_in2,
        Din3 => VN518_in3,
        Din4 => VN518_in4,
        Din5 => VN518_in5,
        VN2CN0_bit => VN_data_out(3108),
        VN2CN1_bit => VN_data_out(3109),
        VN2CN2_bit => VN_data_out(3110),
        VN2CN3_bit => VN_data_out(3111),
        VN2CN4_bit => VN_data_out(3112),
        VN2CN5_bit => VN_data_out(3113),
        VN2CN0_sign => VN_sign_out(3108),
        VN2CN1_sign => VN_sign_out(3109),
        VN2CN2_sign => VN_sign_out(3110),
        VN2CN3_sign => VN_sign_out(3111),
        VN2CN4_sign => VN_sign_out(3112),
        VN2CN5_sign => VN_sign_out(3113),
        codeword => codeword(518),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN519 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3119 downto 3114),
        Din0 => VN519_in0,
        Din1 => VN519_in1,
        Din2 => VN519_in2,
        Din3 => VN519_in3,
        Din4 => VN519_in4,
        Din5 => VN519_in5,
        VN2CN0_bit => VN_data_out(3114),
        VN2CN1_bit => VN_data_out(3115),
        VN2CN2_bit => VN_data_out(3116),
        VN2CN3_bit => VN_data_out(3117),
        VN2CN4_bit => VN_data_out(3118),
        VN2CN5_bit => VN_data_out(3119),
        VN2CN0_sign => VN_sign_out(3114),
        VN2CN1_sign => VN_sign_out(3115),
        VN2CN2_sign => VN_sign_out(3116),
        VN2CN3_sign => VN_sign_out(3117),
        VN2CN4_sign => VN_sign_out(3118),
        VN2CN5_sign => VN_sign_out(3119),
        codeword => codeword(519),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN520 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3125 downto 3120),
        Din0 => VN520_in0,
        Din1 => VN520_in1,
        Din2 => VN520_in2,
        Din3 => VN520_in3,
        Din4 => VN520_in4,
        Din5 => VN520_in5,
        VN2CN0_bit => VN_data_out(3120),
        VN2CN1_bit => VN_data_out(3121),
        VN2CN2_bit => VN_data_out(3122),
        VN2CN3_bit => VN_data_out(3123),
        VN2CN4_bit => VN_data_out(3124),
        VN2CN5_bit => VN_data_out(3125),
        VN2CN0_sign => VN_sign_out(3120),
        VN2CN1_sign => VN_sign_out(3121),
        VN2CN2_sign => VN_sign_out(3122),
        VN2CN3_sign => VN_sign_out(3123),
        VN2CN4_sign => VN_sign_out(3124),
        VN2CN5_sign => VN_sign_out(3125),
        codeword => codeword(520),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN521 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3131 downto 3126),
        Din0 => VN521_in0,
        Din1 => VN521_in1,
        Din2 => VN521_in2,
        Din3 => VN521_in3,
        Din4 => VN521_in4,
        Din5 => VN521_in5,
        VN2CN0_bit => VN_data_out(3126),
        VN2CN1_bit => VN_data_out(3127),
        VN2CN2_bit => VN_data_out(3128),
        VN2CN3_bit => VN_data_out(3129),
        VN2CN4_bit => VN_data_out(3130),
        VN2CN5_bit => VN_data_out(3131),
        VN2CN0_sign => VN_sign_out(3126),
        VN2CN1_sign => VN_sign_out(3127),
        VN2CN2_sign => VN_sign_out(3128),
        VN2CN3_sign => VN_sign_out(3129),
        VN2CN4_sign => VN_sign_out(3130),
        VN2CN5_sign => VN_sign_out(3131),
        codeword => codeword(521),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN522 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3137 downto 3132),
        Din0 => VN522_in0,
        Din1 => VN522_in1,
        Din2 => VN522_in2,
        Din3 => VN522_in3,
        Din4 => VN522_in4,
        Din5 => VN522_in5,
        VN2CN0_bit => VN_data_out(3132),
        VN2CN1_bit => VN_data_out(3133),
        VN2CN2_bit => VN_data_out(3134),
        VN2CN3_bit => VN_data_out(3135),
        VN2CN4_bit => VN_data_out(3136),
        VN2CN5_bit => VN_data_out(3137),
        VN2CN0_sign => VN_sign_out(3132),
        VN2CN1_sign => VN_sign_out(3133),
        VN2CN2_sign => VN_sign_out(3134),
        VN2CN3_sign => VN_sign_out(3135),
        VN2CN4_sign => VN_sign_out(3136),
        VN2CN5_sign => VN_sign_out(3137),
        codeword => codeword(522),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN523 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3143 downto 3138),
        Din0 => VN523_in0,
        Din1 => VN523_in1,
        Din2 => VN523_in2,
        Din3 => VN523_in3,
        Din4 => VN523_in4,
        Din5 => VN523_in5,
        VN2CN0_bit => VN_data_out(3138),
        VN2CN1_bit => VN_data_out(3139),
        VN2CN2_bit => VN_data_out(3140),
        VN2CN3_bit => VN_data_out(3141),
        VN2CN4_bit => VN_data_out(3142),
        VN2CN5_bit => VN_data_out(3143),
        VN2CN0_sign => VN_sign_out(3138),
        VN2CN1_sign => VN_sign_out(3139),
        VN2CN2_sign => VN_sign_out(3140),
        VN2CN3_sign => VN_sign_out(3141),
        VN2CN4_sign => VN_sign_out(3142),
        VN2CN5_sign => VN_sign_out(3143),
        codeword => codeword(523),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN524 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3149 downto 3144),
        Din0 => VN524_in0,
        Din1 => VN524_in1,
        Din2 => VN524_in2,
        Din3 => VN524_in3,
        Din4 => VN524_in4,
        Din5 => VN524_in5,
        VN2CN0_bit => VN_data_out(3144),
        VN2CN1_bit => VN_data_out(3145),
        VN2CN2_bit => VN_data_out(3146),
        VN2CN3_bit => VN_data_out(3147),
        VN2CN4_bit => VN_data_out(3148),
        VN2CN5_bit => VN_data_out(3149),
        VN2CN0_sign => VN_sign_out(3144),
        VN2CN1_sign => VN_sign_out(3145),
        VN2CN2_sign => VN_sign_out(3146),
        VN2CN3_sign => VN_sign_out(3147),
        VN2CN4_sign => VN_sign_out(3148),
        VN2CN5_sign => VN_sign_out(3149),
        codeword => codeword(524),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN525 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3155 downto 3150),
        Din0 => VN525_in0,
        Din1 => VN525_in1,
        Din2 => VN525_in2,
        Din3 => VN525_in3,
        Din4 => VN525_in4,
        Din5 => VN525_in5,
        VN2CN0_bit => VN_data_out(3150),
        VN2CN1_bit => VN_data_out(3151),
        VN2CN2_bit => VN_data_out(3152),
        VN2CN3_bit => VN_data_out(3153),
        VN2CN4_bit => VN_data_out(3154),
        VN2CN5_bit => VN_data_out(3155),
        VN2CN0_sign => VN_sign_out(3150),
        VN2CN1_sign => VN_sign_out(3151),
        VN2CN2_sign => VN_sign_out(3152),
        VN2CN3_sign => VN_sign_out(3153),
        VN2CN4_sign => VN_sign_out(3154),
        VN2CN5_sign => VN_sign_out(3155),
        codeword => codeword(525),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN526 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3161 downto 3156),
        Din0 => VN526_in0,
        Din1 => VN526_in1,
        Din2 => VN526_in2,
        Din3 => VN526_in3,
        Din4 => VN526_in4,
        Din5 => VN526_in5,
        VN2CN0_bit => VN_data_out(3156),
        VN2CN1_bit => VN_data_out(3157),
        VN2CN2_bit => VN_data_out(3158),
        VN2CN3_bit => VN_data_out(3159),
        VN2CN4_bit => VN_data_out(3160),
        VN2CN5_bit => VN_data_out(3161),
        VN2CN0_sign => VN_sign_out(3156),
        VN2CN1_sign => VN_sign_out(3157),
        VN2CN2_sign => VN_sign_out(3158),
        VN2CN3_sign => VN_sign_out(3159),
        VN2CN4_sign => VN_sign_out(3160),
        VN2CN5_sign => VN_sign_out(3161),
        codeword => codeword(526),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN527 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3167 downto 3162),
        Din0 => VN527_in0,
        Din1 => VN527_in1,
        Din2 => VN527_in2,
        Din3 => VN527_in3,
        Din4 => VN527_in4,
        Din5 => VN527_in5,
        VN2CN0_bit => VN_data_out(3162),
        VN2CN1_bit => VN_data_out(3163),
        VN2CN2_bit => VN_data_out(3164),
        VN2CN3_bit => VN_data_out(3165),
        VN2CN4_bit => VN_data_out(3166),
        VN2CN5_bit => VN_data_out(3167),
        VN2CN0_sign => VN_sign_out(3162),
        VN2CN1_sign => VN_sign_out(3163),
        VN2CN2_sign => VN_sign_out(3164),
        VN2CN3_sign => VN_sign_out(3165),
        VN2CN4_sign => VN_sign_out(3166),
        VN2CN5_sign => VN_sign_out(3167),
        codeword => codeword(527),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN528 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3173 downto 3168),
        Din0 => VN528_in0,
        Din1 => VN528_in1,
        Din2 => VN528_in2,
        Din3 => VN528_in3,
        Din4 => VN528_in4,
        Din5 => VN528_in5,
        VN2CN0_bit => VN_data_out(3168),
        VN2CN1_bit => VN_data_out(3169),
        VN2CN2_bit => VN_data_out(3170),
        VN2CN3_bit => VN_data_out(3171),
        VN2CN4_bit => VN_data_out(3172),
        VN2CN5_bit => VN_data_out(3173),
        VN2CN0_sign => VN_sign_out(3168),
        VN2CN1_sign => VN_sign_out(3169),
        VN2CN2_sign => VN_sign_out(3170),
        VN2CN3_sign => VN_sign_out(3171),
        VN2CN4_sign => VN_sign_out(3172),
        VN2CN5_sign => VN_sign_out(3173),
        codeword => codeword(528),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN529 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3179 downto 3174),
        Din0 => VN529_in0,
        Din1 => VN529_in1,
        Din2 => VN529_in2,
        Din3 => VN529_in3,
        Din4 => VN529_in4,
        Din5 => VN529_in5,
        VN2CN0_bit => VN_data_out(3174),
        VN2CN1_bit => VN_data_out(3175),
        VN2CN2_bit => VN_data_out(3176),
        VN2CN3_bit => VN_data_out(3177),
        VN2CN4_bit => VN_data_out(3178),
        VN2CN5_bit => VN_data_out(3179),
        VN2CN0_sign => VN_sign_out(3174),
        VN2CN1_sign => VN_sign_out(3175),
        VN2CN2_sign => VN_sign_out(3176),
        VN2CN3_sign => VN_sign_out(3177),
        VN2CN4_sign => VN_sign_out(3178),
        VN2CN5_sign => VN_sign_out(3179),
        codeword => codeword(529),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN530 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3185 downto 3180),
        Din0 => VN530_in0,
        Din1 => VN530_in1,
        Din2 => VN530_in2,
        Din3 => VN530_in3,
        Din4 => VN530_in4,
        Din5 => VN530_in5,
        VN2CN0_bit => VN_data_out(3180),
        VN2CN1_bit => VN_data_out(3181),
        VN2CN2_bit => VN_data_out(3182),
        VN2CN3_bit => VN_data_out(3183),
        VN2CN4_bit => VN_data_out(3184),
        VN2CN5_bit => VN_data_out(3185),
        VN2CN0_sign => VN_sign_out(3180),
        VN2CN1_sign => VN_sign_out(3181),
        VN2CN2_sign => VN_sign_out(3182),
        VN2CN3_sign => VN_sign_out(3183),
        VN2CN4_sign => VN_sign_out(3184),
        VN2CN5_sign => VN_sign_out(3185),
        codeword => codeword(530),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN531 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3191 downto 3186),
        Din0 => VN531_in0,
        Din1 => VN531_in1,
        Din2 => VN531_in2,
        Din3 => VN531_in3,
        Din4 => VN531_in4,
        Din5 => VN531_in5,
        VN2CN0_bit => VN_data_out(3186),
        VN2CN1_bit => VN_data_out(3187),
        VN2CN2_bit => VN_data_out(3188),
        VN2CN3_bit => VN_data_out(3189),
        VN2CN4_bit => VN_data_out(3190),
        VN2CN5_bit => VN_data_out(3191),
        VN2CN0_sign => VN_sign_out(3186),
        VN2CN1_sign => VN_sign_out(3187),
        VN2CN2_sign => VN_sign_out(3188),
        VN2CN3_sign => VN_sign_out(3189),
        VN2CN4_sign => VN_sign_out(3190),
        VN2CN5_sign => VN_sign_out(3191),
        codeword => codeword(531),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN532 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3197 downto 3192),
        Din0 => VN532_in0,
        Din1 => VN532_in1,
        Din2 => VN532_in2,
        Din3 => VN532_in3,
        Din4 => VN532_in4,
        Din5 => VN532_in5,
        VN2CN0_bit => VN_data_out(3192),
        VN2CN1_bit => VN_data_out(3193),
        VN2CN2_bit => VN_data_out(3194),
        VN2CN3_bit => VN_data_out(3195),
        VN2CN4_bit => VN_data_out(3196),
        VN2CN5_bit => VN_data_out(3197),
        VN2CN0_sign => VN_sign_out(3192),
        VN2CN1_sign => VN_sign_out(3193),
        VN2CN2_sign => VN_sign_out(3194),
        VN2CN3_sign => VN_sign_out(3195),
        VN2CN4_sign => VN_sign_out(3196),
        VN2CN5_sign => VN_sign_out(3197),
        codeword => codeword(532),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN533 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3203 downto 3198),
        Din0 => VN533_in0,
        Din1 => VN533_in1,
        Din2 => VN533_in2,
        Din3 => VN533_in3,
        Din4 => VN533_in4,
        Din5 => VN533_in5,
        VN2CN0_bit => VN_data_out(3198),
        VN2CN1_bit => VN_data_out(3199),
        VN2CN2_bit => VN_data_out(3200),
        VN2CN3_bit => VN_data_out(3201),
        VN2CN4_bit => VN_data_out(3202),
        VN2CN5_bit => VN_data_out(3203),
        VN2CN0_sign => VN_sign_out(3198),
        VN2CN1_sign => VN_sign_out(3199),
        VN2CN2_sign => VN_sign_out(3200),
        VN2CN3_sign => VN_sign_out(3201),
        VN2CN4_sign => VN_sign_out(3202),
        VN2CN5_sign => VN_sign_out(3203),
        codeword => codeword(533),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN534 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3209 downto 3204),
        Din0 => VN534_in0,
        Din1 => VN534_in1,
        Din2 => VN534_in2,
        Din3 => VN534_in3,
        Din4 => VN534_in4,
        Din5 => VN534_in5,
        VN2CN0_bit => VN_data_out(3204),
        VN2CN1_bit => VN_data_out(3205),
        VN2CN2_bit => VN_data_out(3206),
        VN2CN3_bit => VN_data_out(3207),
        VN2CN4_bit => VN_data_out(3208),
        VN2CN5_bit => VN_data_out(3209),
        VN2CN0_sign => VN_sign_out(3204),
        VN2CN1_sign => VN_sign_out(3205),
        VN2CN2_sign => VN_sign_out(3206),
        VN2CN3_sign => VN_sign_out(3207),
        VN2CN4_sign => VN_sign_out(3208),
        VN2CN5_sign => VN_sign_out(3209),
        codeword => codeword(534),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN535 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3215 downto 3210),
        Din0 => VN535_in0,
        Din1 => VN535_in1,
        Din2 => VN535_in2,
        Din3 => VN535_in3,
        Din4 => VN535_in4,
        Din5 => VN535_in5,
        VN2CN0_bit => VN_data_out(3210),
        VN2CN1_bit => VN_data_out(3211),
        VN2CN2_bit => VN_data_out(3212),
        VN2CN3_bit => VN_data_out(3213),
        VN2CN4_bit => VN_data_out(3214),
        VN2CN5_bit => VN_data_out(3215),
        VN2CN0_sign => VN_sign_out(3210),
        VN2CN1_sign => VN_sign_out(3211),
        VN2CN2_sign => VN_sign_out(3212),
        VN2CN3_sign => VN_sign_out(3213),
        VN2CN4_sign => VN_sign_out(3214),
        VN2CN5_sign => VN_sign_out(3215),
        codeword => codeword(535),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN536 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3221 downto 3216),
        Din0 => VN536_in0,
        Din1 => VN536_in1,
        Din2 => VN536_in2,
        Din3 => VN536_in3,
        Din4 => VN536_in4,
        Din5 => VN536_in5,
        VN2CN0_bit => VN_data_out(3216),
        VN2CN1_bit => VN_data_out(3217),
        VN2CN2_bit => VN_data_out(3218),
        VN2CN3_bit => VN_data_out(3219),
        VN2CN4_bit => VN_data_out(3220),
        VN2CN5_bit => VN_data_out(3221),
        VN2CN0_sign => VN_sign_out(3216),
        VN2CN1_sign => VN_sign_out(3217),
        VN2CN2_sign => VN_sign_out(3218),
        VN2CN3_sign => VN_sign_out(3219),
        VN2CN4_sign => VN_sign_out(3220),
        VN2CN5_sign => VN_sign_out(3221),
        codeword => codeword(536),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN537 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3227 downto 3222),
        Din0 => VN537_in0,
        Din1 => VN537_in1,
        Din2 => VN537_in2,
        Din3 => VN537_in3,
        Din4 => VN537_in4,
        Din5 => VN537_in5,
        VN2CN0_bit => VN_data_out(3222),
        VN2CN1_bit => VN_data_out(3223),
        VN2CN2_bit => VN_data_out(3224),
        VN2CN3_bit => VN_data_out(3225),
        VN2CN4_bit => VN_data_out(3226),
        VN2CN5_bit => VN_data_out(3227),
        VN2CN0_sign => VN_sign_out(3222),
        VN2CN1_sign => VN_sign_out(3223),
        VN2CN2_sign => VN_sign_out(3224),
        VN2CN3_sign => VN_sign_out(3225),
        VN2CN4_sign => VN_sign_out(3226),
        VN2CN5_sign => VN_sign_out(3227),
        codeword => codeword(537),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN538 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3233 downto 3228),
        Din0 => VN538_in0,
        Din1 => VN538_in1,
        Din2 => VN538_in2,
        Din3 => VN538_in3,
        Din4 => VN538_in4,
        Din5 => VN538_in5,
        VN2CN0_bit => VN_data_out(3228),
        VN2CN1_bit => VN_data_out(3229),
        VN2CN2_bit => VN_data_out(3230),
        VN2CN3_bit => VN_data_out(3231),
        VN2CN4_bit => VN_data_out(3232),
        VN2CN5_bit => VN_data_out(3233),
        VN2CN0_sign => VN_sign_out(3228),
        VN2CN1_sign => VN_sign_out(3229),
        VN2CN2_sign => VN_sign_out(3230),
        VN2CN3_sign => VN_sign_out(3231),
        VN2CN4_sign => VN_sign_out(3232),
        VN2CN5_sign => VN_sign_out(3233),
        codeword => codeword(538),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN539 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3239 downto 3234),
        Din0 => VN539_in0,
        Din1 => VN539_in1,
        Din2 => VN539_in2,
        Din3 => VN539_in3,
        Din4 => VN539_in4,
        Din5 => VN539_in5,
        VN2CN0_bit => VN_data_out(3234),
        VN2CN1_bit => VN_data_out(3235),
        VN2CN2_bit => VN_data_out(3236),
        VN2CN3_bit => VN_data_out(3237),
        VN2CN4_bit => VN_data_out(3238),
        VN2CN5_bit => VN_data_out(3239),
        VN2CN0_sign => VN_sign_out(3234),
        VN2CN1_sign => VN_sign_out(3235),
        VN2CN2_sign => VN_sign_out(3236),
        VN2CN3_sign => VN_sign_out(3237),
        VN2CN4_sign => VN_sign_out(3238),
        VN2CN5_sign => VN_sign_out(3239),
        codeword => codeword(539),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN540 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3245 downto 3240),
        Din0 => VN540_in0,
        Din1 => VN540_in1,
        Din2 => VN540_in2,
        Din3 => VN540_in3,
        Din4 => VN540_in4,
        Din5 => VN540_in5,
        VN2CN0_bit => VN_data_out(3240),
        VN2CN1_bit => VN_data_out(3241),
        VN2CN2_bit => VN_data_out(3242),
        VN2CN3_bit => VN_data_out(3243),
        VN2CN4_bit => VN_data_out(3244),
        VN2CN5_bit => VN_data_out(3245),
        VN2CN0_sign => VN_sign_out(3240),
        VN2CN1_sign => VN_sign_out(3241),
        VN2CN2_sign => VN_sign_out(3242),
        VN2CN3_sign => VN_sign_out(3243),
        VN2CN4_sign => VN_sign_out(3244),
        VN2CN5_sign => VN_sign_out(3245),
        codeword => codeword(540),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN541 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3251 downto 3246),
        Din0 => VN541_in0,
        Din1 => VN541_in1,
        Din2 => VN541_in2,
        Din3 => VN541_in3,
        Din4 => VN541_in4,
        Din5 => VN541_in5,
        VN2CN0_bit => VN_data_out(3246),
        VN2CN1_bit => VN_data_out(3247),
        VN2CN2_bit => VN_data_out(3248),
        VN2CN3_bit => VN_data_out(3249),
        VN2CN4_bit => VN_data_out(3250),
        VN2CN5_bit => VN_data_out(3251),
        VN2CN0_sign => VN_sign_out(3246),
        VN2CN1_sign => VN_sign_out(3247),
        VN2CN2_sign => VN_sign_out(3248),
        VN2CN3_sign => VN_sign_out(3249),
        VN2CN4_sign => VN_sign_out(3250),
        VN2CN5_sign => VN_sign_out(3251),
        codeword => codeword(541),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN542 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3257 downto 3252),
        Din0 => VN542_in0,
        Din1 => VN542_in1,
        Din2 => VN542_in2,
        Din3 => VN542_in3,
        Din4 => VN542_in4,
        Din5 => VN542_in5,
        VN2CN0_bit => VN_data_out(3252),
        VN2CN1_bit => VN_data_out(3253),
        VN2CN2_bit => VN_data_out(3254),
        VN2CN3_bit => VN_data_out(3255),
        VN2CN4_bit => VN_data_out(3256),
        VN2CN5_bit => VN_data_out(3257),
        VN2CN0_sign => VN_sign_out(3252),
        VN2CN1_sign => VN_sign_out(3253),
        VN2CN2_sign => VN_sign_out(3254),
        VN2CN3_sign => VN_sign_out(3255),
        VN2CN4_sign => VN_sign_out(3256),
        VN2CN5_sign => VN_sign_out(3257),
        codeword => codeword(542),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN543 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3263 downto 3258),
        Din0 => VN543_in0,
        Din1 => VN543_in1,
        Din2 => VN543_in2,
        Din3 => VN543_in3,
        Din4 => VN543_in4,
        Din5 => VN543_in5,
        VN2CN0_bit => VN_data_out(3258),
        VN2CN1_bit => VN_data_out(3259),
        VN2CN2_bit => VN_data_out(3260),
        VN2CN3_bit => VN_data_out(3261),
        VN2CN4_bit => VN_data_out(3262),
        VN2CN5_bit => VN_data_out(3263),
        VN2CN0_sign => VN_sign_out(3258),
        VN2CN1_sign => VN_sign_out(3259),
        VN2CN2_sign => VN_sign_out(3260),
        VN2CN3_sign => VN_sign_out(3261),
        VN2CN4_sign => VN_sign_out(3262),
        VN2CN5_sign => VN_sign_out(3263),
        codeword => codeword(543),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN544 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3269 downto 3264),
        Din0 => VN544_in0,
        Din1 => VN544_in1,
        Din2 => VN544_in2,
        Din3 => VN544_in3,
        Din4 => VN544_in4,
        Din5 => VN544_in5,
        VN2CN0_bit => VN_data_out(3264),
        VN2CN1_bit => VN_data_out(3265),
        VN2CN2_bit => VN_data_out(3266),
        VN2CN3_bit => VN_data_out(3267),
        VN2CN4_bit => VN_data_out(3268),
        VN2CN5_bit => VN_data_out(3269),
        VN2CN0_sign => VN_sign_out(3264),
        VN2CN1_sign => VN_sign_out(3265),
        VN2CN2_sign => VN_sign_out(3266),
        VN2CN3_sign => VN_sign_out(3267),
        VN2CN4_sign => VN_sign_out(3268),
        VN2CN5_sign => VN_sign_out(3269),
        codeword => codeword(544),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN545 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3275 downto 3270),
        Din0 => VN545_in0,
        Din1 => VN545_in1,
        Din2 => VN545_in2,
        Din3 => VN545_in3,
        Din4 => VN545_in4,
        Din5 => VN545_in5,
        VN2CN0_bit => VN_data_out(3270),
        VN2CN1_bit => VN_data_out(3271),
        VN2CN2_bit => VN_data_out(3272),
        VN2CN3_bit => VN_data_out(3273),
        VN2CN4_bit => VN_data_out(3274),
        VN2CN5_bit => VN_data_out(3275),
        VN2CN0_sign => VN_sign_out(3270),
        VN2CN1_sign => VN_sign_out(3271),
        VN2CN2_sign => VN_sign_out(3272),
        VN2CN3_sign => VN_sign_out(3273),
        VN2CN4_sign => VN_sign_out(3274),
        VN2CN5_sign => VN_sign_out(3275),
        codeword => codeword(545),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN546 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3281 downto 3276),
        Din0 => VN546_in0,
        Din1 => VN546_in1,
        Din2 => VN546_in2,
        Din3 => VN546_in3,
        Din4 => VN546_in4,
        Din5 => VN546_in5,
        VN2CN0_bit => VN_data_out(3276),
        VN2CN1_bit => VN_data_out(3277),
        VN2CN2_bit => VN_data_out(3278),
        VN2CN3_bit => VN_data_out(3279),
        VN2CN4_bit => VN_data_out(3280),
        VN2CN5_bit => VN_data_out(3281),
        VN2CN0_sign => VN_sign_out(3276),
        VN2CN1_sign => VN_sign_out(3277),
        VN2CN2_sign => VN_sign_out(3278),
        VN2CN3_sign => VN_sign_out(3279),
        VN2CN4_sign => VN_sign_out(3280),
        VN2CN5_sign => VN_sign_out(3281),
        codeword => codeword(546),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN547 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3287 downto 3282),
        Din0 => VN547_in0,
        Din1 => VN547_in1,
        Din2 => VN547_in2,
        Din3 => VN547_in3,
        Din4 => VN547_in4,
        Din5 => VN547_in5,
        VN2CN0_bit => VN_data_out(3282),
        VN2CN1_bit => VN_data_out(3283),
        VN2CN2_bit => VN_data_out(3284),
        VN2CN3_bit => VN_data_out(3285),
        VN2CN4_bit => VN_data_out(3286),
        VN2CN5_bit => VN_data_out(3287),
        VN2CN0_sign => VN_sign_out(3282),
        VN2CN1_sign => VN_sign_out(3283),
        VN2CN2_sign => VN_sign_out(3284),
        VN2CN3_sign => VN_sign_out(3285),
        VN2CN4_sign => VN_sign_out(3286),
        VN2CN5_sign => VN_sign_out(3287),
        codeword => codeword(547),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN548 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3293 downto 3288),
        Din0 => VN548_in0,
        Din1 => VN548_in1,
        Din2 => VN548_in2,
        Din3 => VN548_in3,
        Din4 => VN548_in4,
        Din5 => VN548_in5,
        VN2CN0_bit => VN_data_out(3288),
        VN2CN1_bit => VN_data_out(3289),
        VN2CN2_bit => VN_data_out(3290),
        VN2CN3_bit => VN_data_out(3291),
        VN2CN4_bit => VN_data_out(3292),
        VN2CN5_bit => VN_data_out(3293),
        VN2CN0_sign => VN_sign_out(3288),
        VN2CN1_sign => VN_sign_out(3289),
        VN2CN2_sign => VN_sign_out(3290),
        VN2CN3_sign => VN_sign_out(3291),
        VN2CN4_sign => VN_sign_out(3292),
        VN2CN5_sign => VN_sign_out(3293),
        codeword => codeword(548),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN549 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3299 downto 3294),
        Din0 => VN549_in0,
        Din1 => VN549_in1,
        Din2 => VN549_in2,
        Din3 => VN549_in3,
        Din4 => VN549_in4,
        Din5 => VN549_in5,
        VN2CN0_bit => VN_data_out(3294),
        VN2CN1_bit => VN_data_out(3295),
        VN2CN2_bit => VN_data_out(3296),
        VN2CN3_bit => VN_data_out(3297),
        VN2CN4_bit => VN_data_out(3298),
        VN2CN5_bit => VN_data_out(3299),
        VN2CN0_sign => VN_sign_out(3294),
        VN2CN1_sign => VN_sign_out(3295),
        VN2CN2_sign => VN_sign_out(3296),
        VN2CN3_sign => VN_sign_out(3297),
        VN2CN4_sign => VN_sign_out(3298),
        VN2CN5_sign => VN_sign_out(3299),
        codeword => codeword(549),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN550 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3305 downto 3300),
        Din0 => VN550_in0,
        Din1 => VN550_in1,
        Din2 => VN550_in2,
        Din3 => VN550_in3,
        Din4 => VN550_in4,
        Din5 => VN550_in5,
        VN2CN0_bit => VN_data_out(3300),
        VN2CN1_bit => VN_data_out(3301),
        VN2CN2_bit => VN_data_out(3302),
        VN2CN3_bit => VN_data_out(3303),
        VN2CN4_bit => VN_data_out(3304),
        VN2CN5_bit => VN_data_out(3305),
        VN2CN0_sign => VN_sign_out(3300),
        VN2CN1_sign => VN_sign_out(3301),
        VN2CN2_sign => VN_sign_out(3302),
        VN2CN3_sign => VN_sign_out(3303),
        VN2CN4_sign => VN_sign_out(3304),
        VN2CN5_sign => VN_sign_out(3305),
        codeword => codeword(550),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN551 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3311 downto 3306),
        Din0 => VN551_in0,
        Din1 => VN551_in1,
        Din2 => VN551_in2,
        Din3 => VN551_in3,
        Din4 => VN551_in4,
        Din5 => VN551_in5,
        VN2CN0_bit => VN_data_out(3306),
        VN2CN1_bit => VN_data_out(3307),
        VN2CN2_bit => VN_data_out(3308),
        VN2CN3_bit => VN_data_out(3309),
        VN2CN4_bit => VN_data_out(3310),
        VN2CN5_bit => VN_data_out(3311),
        VN2CN0_sign => VN_sign_out(3306),
        VN2CN1_sign => VN_sign_out(3307),
        VN2CN2_sign => VN_sign_out(3308),
        VN2CN3_sign => VN_sign_out(3309),
        VN2CN4_sign => VN_sign_out(3310),
        VN2CN5_sign => VN_sign_out(3311),
        codeword => codeword(551),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN552 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3317 downto 3312),
        Din0 => VN552_in0,
        Din1 => VN552_in1,
        Din2 => VN552_in2,
        Din3 => VN552_in3,
        Din4 => VN552_in4,
        Din5 => VN552_in5,
        VN2CN0_bit => VN_data_out(3312),
        VN2CN1_bit => VN_data_out(3313),
        VN2CN2_bit => VN_data_out(3314),
        VN2CN3_bit => VN_data_out(3315),
        VN2CN4_bit => VN_data_out(3316),
        VN2CN5_bit => VN_data_out(3317),
        VN2CN0_sign => VN_sign_out(3312),
        VN2CN1_sign => VN_sign_out(3313),
        VN2CN2_sign => VN_sign_out(3314),
        VN2CN3_sign => VN_sign_out(3315),
        VN2CN4_sign => VN_sign_out(3316),
        VN2CN5_sign => VN_sign_out(3317),
        codeword => codeword(552),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN553 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3323 downto 3318),
        Din0 => VN553_in0,
        Din1 => VN553_in1,
        Din2 => VN553_in2,
        Din3 => VN553_in3,
        Din4 => VN553_in4,
        Din5 => VN553_in5,
        VN2CN0_bit => VN_data_out(3318),
        VN2CN1_bit => VN_data_out(3319),
        VN2CN2_bit => VN_data_out(3320),
        VN2CN3_bit => VN_data_out(3321),
        VN2CN4_bit => VN_data_out(3322),
        VN2CN5_bit => VN_data_out(3323),
        VN2CN0_sign => VN_sign_out(3318),
        VN2CN1_sign => VN_sign_out(3319),
        VN2CN2_sign => VN_sign_out(3320),
        VN2CN3_sign => VN_sign_out(3321),
        VN2CN4_sign => VN_sign_out(3322),
        VN2CN5_sign => VN_sign_out(3323),
        codeword => codeword(553),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN554 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3329 downto 3324),
        Din0 => VN554_in0,
        Din1 => VN554_in1,
        Din2 => VN554_in2,
        Din3 => VN554_in3,
        Din4 => VN554_in4,
        Din5 => VN554_in5,
        VN2CN0_bit => VN_data_out(3324),
        VN2CN1_bit => VN_data_out(3325),
        VN2CN2_bit => VN_data_out(3326),
        VN2CN3_bit => VN_data_out(3327),
        VN2CN4_bit => VN_data_out(3328),
        VN2CN5_bit => VN_data_out(3329),
        VN2CN0_sign => VN_sign_out(3324),
        VN2CN1_sign => VN_sign_out(3325),
        VN2CN2_sign => VN_sign_out(3326),
        VN2CN3_sign => VN_sign_out(3327),
        VN2CN4_sign => VN_sign_out(3328),
        VN2CN5_sign => VN_sign_out(3329),
        codeword => codeword(554),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN555 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3335 downto 3330),
        Din0 => VN555_in0,
        Din1 => VN555_in1,
        Din2 => VN555_in2,
        Din3 => VN555_in3,
        Din4 => VN555_in4,
        Din5 => VN555_in5,
        VN2CN0_bit => VN_data_out(3330),
        VN2CN1_bit => VN_data_out(3331),
        VN2CN2_bit => VN_data_out(3332),
        VN2CN3_bit => VN_data_out(3333),
        VN2CN4_bit => VN_data_out(3334),
        VN2CN5_bit => VN_data_out(3335),
        VN2CN0_sign => VN_sign_out(3330),
        VN2CN1_sign => VN_sign_out(3331),
        VN2CN2_sign => VN_sign_out(3332),
        VN2CN3_sign => VN_sign_out(3333),
        VN2CN4_sign => VN_sign_out(3334),
        VN2CN5_sign => VN_sign_out(3335),
        codeword => codeword(555),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN556 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3341 downto 3336),
        Din0 => VN556_in0,
        Din1 => VN556_in1,
        Din2 => VN556_in2,
        Din3 => VN556_in3,
        Din4 => VN556_in4,
        Din5 => VN556_in5,
        VN2CN0_bit => VN_data_out(3336),
        VN2CN1_bit => VN_data_out(3337),
        VN2CN2_bit => VN_data_out(3338),
        VN2CN3_bit => VN_data_out(3339),
        VN2CN4_bit => VN_data_out(3340),
        VN2CN5_bit => VN_data_out(3341),
        VN2CN0_sign => VN_sign_out(3336),
        VN2CN1_sign => VN_sign_out(3337),
        VN2CN2_sign => VN_sign_out(3338),
        VN2CN3_sign => VN_sign_out(3339),
        VN2CN4_sign => VN_sign_out(3340),
        VN2CN5_sign => VN_sign_out(3341),
        codeword => codeword(556),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN557 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3347 downto 3342),
        Din0 => VN557_in0,
        Din1 => VN557_in1,
        Din2 => VN557_in2,
        Din3 => VN557_in3,
        Din4 => VN557_in4,
        Din5 => VN557_in5,
        VN2CN0_bit => VN_data_out(3342),
        VN2CN1_bit => VN_data_out(3343),
        VN2CN2_bit => VN_data_out(3344),
        VN2CN3_bit => VN_data_out(3345),
        VN2CN4_bit => VN_data_out(3346),
        VN2CN5_bit => VN_data_out(3347),
        VN2CN0_sign => VN_sign_out(3342),
        VN2CN1_sign => VN_sign_out(3343),
        VN2CN2_sign => VN_sign_out(3344),
        VN2CN3_sign => VN_sign_out(3345),
        VN2CN4_sign => VN_sign_out(3346),
        VN2CN5_sign => VN_sign_out(3347),
        codeword => codeword(557),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN558 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3353 downto 3348),
        Din0 => VN558_in0,
        Din1 => VN558_in1,
        Din2 => VN558_in2,
        Din3 => VN558_in3,
        Din4 => VN558_in4,
        Din5 => VN558_in5,
        VN2CN0_bit => VN_data_out(3348),
        VN2CN1_bit => VN_data_out(3349),
        VN2CN2_bit => VN_data_out(3350),
        VN2CN3_bit => VN_data_out(3351),
        VN2CN4_bit => VN_data_out(3352),
        VN2CN5_bit => VN_data_out(3353),
        VN2CN0_sign => VN_sign_out(3348),
        VN2CN1_sign => VN_sign_out(3349),
        VN2CN2_sign => VN_sign_out(3350),
        VN2CN3_sign => VN_sign_out(3351),
        VN2CN4_sign => VN_sign_out(3352),
        VN2CN5_sign => VN_sign_out(3353),
        codeword => codeword(558),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN559 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3359 downto 3354),
        Din0 => VN559_in0,
        Din1 => VN559_in1,
        Din2 => VN559_in2,
        Din3 => VN559_in3,
        Din4 => VN559_in4,
        Din5 => VN559_in5,
        VN2CN0_bit => VN_data_out(3354),
        VN2CN1_bit => VN_data_out(3355),
        VN2CN2_bit => VN_data_out(3356),
        VN2CN3_bit => VN_data_out(3357),
        VN2CN4_bit => VN_data_out(3358),
        VN2CN5_bit => VN_data_out(3359),
        VN2CN0_sign => VN_sign_out(3354),
        VN2CN1_sign => VN_sign_out(3355),
        VN2CN2_sign => VN_sign_out(3356),
        VN2CN3_sign => VN_sign_out(3357),
        VN2CN4_sign => VN_sign_out(3358),
        VN2CN5_sign => VN_sign_out(3359),
        codeword => codeword(559),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN560 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3365 downto 3360),
        Din0 => VN560_in0,
        Din1 => VN560_in1,
        Din2 => VN560_in2,
        Din3 => VN560_in3,
        Din4 => VN560_in4,
        Din5 => VN560_in5,
        VN2CN0_bit => VN_data_out(3360),
        VN2CN1_bit => VN_data_out(3361),
        VN2CN2_bit => VN_data_out(3362),
        VN2CN3_bit => VN_data_out(3363),
        VN2CN4_bit => VN_data_out(3364),
        VN2CN5_bit => VN_data_out(3365),
        VN2CN0_sign => VN_sign_out(3360),
        VN2CN1_sign => VN_sign_out(3361),
        VN2CN2_sign => VN_sign_out(3362),
        VN2CN3_sign => VN_sign_out(3363),
        VN2CN4_sign => VN_sign_out(3364),
        VN2CN5_sign => VN_sign_out(3365),
        codeword => codeword(560),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN561 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3371 downto 3366),
        Din0 => VN561_in0,
        Din1 => VN561_in1,
        Din2 => VN561_in2,
        Din3 => VN561_in3,
        Din4 => VN561_in4,
        Din5 => VN561_in5,
        VN2CN0_bit => VN_data_out(3366),
        VN2CN1_bit => VN_data_out(3367),
        VN2CN2_bit => VN_data_out(3368),
        VN2CN3_bit => VN_data_out(3369),
        VN2CN4_bit => VN_data_out(3370),
        VN2CN5_bit => VN_data_out(3371),
        VN2CN0_sign => VN_sign_out(3366),
        VN2CN1_sign => VN_sign_out(3367),
        VN2CN2_sign => VN_sign_out(3368),
        VN2CN3_sign => VN_sign_out(3369),
        VN2CN4_sign => VN_sign_out(3370),
        VN2CN5_sign => VN_sign_out(3371),
        codeword => codeword(561),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN562 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3377 downto 3372),
        Din0 => VN562_in0,
        Din1 => VN562_in1,
        Din2 => VN562_in2,
        Din3 => VN562_in3,
        Din4 => VN562_in4,
        Din5 => VN562_in5,
        VN2CN0_bit => VN_data_out(3372),
        VN2CN1_bit => VN_data_out(3373),
        VN2CN2_bit => VN_data_out(3374),
        VN2CN3_bit => VN_data_out(3375),
        VN2CN4_bit => VN_data_out(3376),
        VN2CN5_bit => VN_data_out(3377),
        VN2CN0_sign => VN_sign_out(3372),
        VN2CN1_sign => VN_sign_out(3373),
        VN2CN2_sign => VN_sign_out(3374),
        VN2CN3_sign => VN_sign_out(3375),
        VN2CN4_sign => VN_sign_out(3376),
        VN2CN5_sign => VN_sign_out(3377),
        codeword => codeword(562),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN563 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3383 downto 3378),
        Din0 => VN563_in0,
        Din1 => VN563_in1,
        Din2 => VN563_in2,
        Din3 => VN563_in3,
        Din4 => VN563_in4,
        Din5 => VN563_in5,
        VN2CN0_bit => VN_data_out(3378),
        VN2CN1_bit => VN_data_out(3379),
        VN2CN2_bit => VN_data_out(3380),
        VN2CN3_bit => VN_data_out(3381),
        VN2CN4_bit => VN_data_out(3382),
        VN2CN5_bit => VN_data_out(3383),
        VN2CN0_sign => VN_sign_out(3378),
        VN2CN1_sign => VN_sign_out(3379),
        VN2CN2_sign => VN_sign_out(3380),
        VN2CN3_sign => VN_sign_out(3381),
        VN2CN4_sign => VN_sign_out(3382),
        VN2CN5_sign => VN_sign_out(3383),
        codeword => codeword(563),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN564 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3389 downto 3384),
        Din0 => VN564_in0,
        Din1 => VN564_in1,
        Din2 => VN564_in2,
        Din3 => VN564_in3,
        Din4 => VN564_in4,
        Din5 => VN564_in5,
        VN2CN0_bit => VN_data_out(3384),
        VN2CN1_bit => VN_data_out(3385),
        VN2CN2_bit => VN_data_out(3386),
        VN2CN3_bit => VN_data_out(3387),
        VN2CN4_bit => VN_data_out(3388),
        VN2CN5_bit => VN_data_out(3389),
        VN2CN0_sign => VN_sign_out(3384),
        VN2CN1_sign => VN_sign_out(3385),
        VN2CN2_sign => VN_sign_out(3386),
        VN2CN3_sign => VN_sign_out(3387),
        VN2CN4_sign => VN_sign_out(3388),
        VN2CN5_sign => VN_sign_out(3389),
        codeword => codeword(564),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN565 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3395 downto 3390),
        Din0 => VN565_in0,
        Din1 => VN565_in1,
        Din2 => VN565_in2,
        Din3 => VN565_in3,
        Din4 => VN565_in4,
        Din5 => VN565_in5,
        VN2CN0_bit => VN_data_out(3390),
        VN2CN1_bit => VN_data_out(3391),
        VN2CN2_bit => VN_data_out(3392),
        VN2CN3_bit => VN_data_out(3393),
        VN2CN4_bit => VN_data_out(3394),
        VN2CN5_bit => VN_data_out(3395),
        VN2CN0_sign => VN_sign_out(3390),
        VN2CN1_sign => VN_sign_out(3391),
        VN2CN2_sign => VN_sign_out(3392),
        VN2CN3_sign => VN_sign_out(3393),
        VN2CN4_sign => VN_sign_out(3394),
        VN2CN5_sign => VN_sign_out(3395),
        codeword => codeword(565),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN566 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3401 downto 3396),
        Din0 => VN566_in0,
        Din1 => VN566_in1,
        Din2 => VN566_in2,
        Din3 => VN566_in3,
        Din4 => VN566_in4,
        Din5 => VN566_in5,
        VN2CN0_bit => VN_data_out(3396),
        VN2CN1_bit => VN_data_out(3397),
        VN2CN2_bit => VN_data_out(3398),
        VN2CN3_bit => VN_data_out(3399),
        VN2CN4_bit => VN_data_out(3400),
        VN2CN5_bit => VN_data_out(3401),
        VN2CN0_sign => VN_sign_out(3396),
        VN2CN1_sign => VN_sign_out(3397),
        VN2CN2_sign => VN_sign_out(3398),
        VN2CN3_sign => VN_sign_out(3399),
        VN2CN4_sign => VN_sign_out(3400),
        VN2CN5_sign => VN_sign_out(3401),
        codeword => codeword(566),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN567 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3407 downto 3402),
        Din0 => VN567_in0,
        Din1 => VN567_in1,
        Din2 => VN567_in2,
        Din3 => VN567_in3,
        Din4 => VN567_in4,
        Din5 => VN567_in5,
        VN2CN0_bit => VN_data_out(3402),
        VN2CN1_bit => VN_data_out(3403),
        VN2CN2_bit => VN_data_out(3404),
        VN2CN3_bit => VN_data_out(3405),
        VN2CN4_bit => VN_data_out(3406),
        VN2CN5_bit => VN_data_out(3407),
        VN2CN0_sign => VN_sign_out(3402),
        VN2CN1_sign => VN_sign_out(3403),
        VN2CN2_sign => VN_sign_out(3404),
        VN2CN3_sign => VN_sign_out(3405),
        VN2CN4_sign => VN_sign_out(3406),
        VN2CN5_sign => VN_sign_out(3407),
        codeword => codeword(567),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN568 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3413 downto 3408),
        Din0 => VN568_in0,
        Din1 => VN568_in1,
        Din2 => VN568_in2,
        Din3 => VN568_in3,
        Din4 => VN568_in4,
        Din5 => VN568_in5,
        VN2CN0_bit => VN_data_out(3408),
        VN2CN1_bit => VN_data_out(3409),
        VN2CN2_bit => VN_data_out(3410),
        VN2CN3_bit => VN_data_out(3411),
        VN2CN4_bit => VN_data_out(3412),
        VN2CN5_bit => VN_data_out(3413),
        VN2CN0_sign => VN_sign_out(3408),
        VN2CN1_sign => VN_sign_out(3409),
        VN2CN2_sign => VN_sign_out(3410),
        VN2CN3_sign => VN_sign_out(3411),
        VN2CN4_sign => VN_sign_out(3412),
        VN2CN5_sign => VN_sign_out(3413),
        codeword => codeword(568),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN569 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3419 downto 3414),
        Din0 => VN569_in0,
        Din1 => VN569_in1,
        Din2 => VN569_in2,
        Din3 => VN569_in3,
        Din4 => VN569_in4,
        Din5 => VN569_in5,
        VN2CN0_bit => VN_data_out(3414),
        VN2CN1_bit => VN_data_out(3415),
        VN2CN2_bit => VN_data_out(3416),
        VN2CN3_bit => VN_data_out(3417),
        VN2CN4_bit => VN_data_out(3418),
        VN2CN5_bit => VN_data_out(3419),
        VN2CN0_sign => VN_sign_out(3414),
        VN2CN1_sign => VN_sign_out(3415),
        VN2CN2_sign => VN_sign_out(3416),
        VN2CN3_sign => VN_sign_out(3417),
        VN2CN4_sign => VN_sign_out(3418),
        VN2CN5_sign => VN_sign_out(3419),
        codeword => codeword(569),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN570 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3425 downto 3420),
        Din0 => VN570_in0,
        Din1 => VN570_in1,
        Din2 => VN570_in2,
        Din3 => VN570_in3,
        Din4 => VN570_in4,
        Din5 => VN570_in5,
        VN2CN0_bit => VN_data_out(3420),
        VN2CN1_bit => VN_data_out(3421),
        VN2CN2_bit => VN_data_out(3422),
        VN2CN3_bit => VN_data_out(3423),
        VN2CN4_bit => VN_data_out(3424),
        VN2CN5_bit => VN_data_out(3425),
        VN2CN0_sign => VN_sign_out(3420),
        VN2CN1_sign => VN_sign_out(3421),
        VN2CN2_sign => VN_sign_out(3422),
        VN2CN3_sign => VN_sign_out(3423),
        VN2CN4_sign => VN_sign_out(3424),
        VN2CN5_sign => VN_sign_out(3425),
        codeword => codeword(570),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN571 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3431 downto 3426),
        Din0 => VN571_in0,
        Din1 => VN571_in1,
        Din2 => VN571_in2,
        Din3 => VN571_in3,
        Din4 => VN571_in4,
        Din5 => VN571_in5,
        VN2CN0_bit => VN_data_out(3426),
        VN2CN1_bit => VN_data_out(3427),
        VN2CN2_bit => VN_data_out(3428),
        VN2CN3_bit => VN_data_out(3429),
        VN2CN4_bit => VN_data_out(3430),
        VN2CN5_bit => VN_data_out(3431),
        VN2CN0_sign => VN_sign_out(3426),
        VN2CN1_sign => VN_sign_out(3427),
        VN2CN2_sign => VN_sign_out(3428),
        VN2CN3_sign => VN_sign_out(3429),
        VN2CN4_sign => VN_sign_out(3430),
        VN2CN5_sign => VN_sign_out(3431),
        codeword => codeword(571),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN572 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3437 downto 3432),
        Din0 => VN572_in0,
        Din1 => VN572_in1,
        Din2 => VN572_in2,
        Din3 => VN572_in3,
        Din4 => VN572_in4,
        Din5 => VN572_in5,
        VN2CN0_bit => VN_data_out(3432),
        VN2CN1_bit => VN_data_out(3433),
        VN2CN2_bit => VN_data_out(3434),
        VN2CN3_bit => VN_data_out(3435),
        VN2CN4_bit => VN_data_out(3436),
        VN2CN5_bit => VN_data_out(3437),
        VN2CN0_sign => VN_sign_out(3432),
        VN2CN1_sign => VN_sign_out(3433),
        VN2CN2_sign => VN_sign_out(3434),
        VN2CN3_sign => VN_sign_out(3435),
        VN2CN4_sign => VN_sign_out(3436),
        VN2CN5_sign => VN_sign_out(3437),
        codeword => codeword(572),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN573 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3443 downto 3438),
        Din0 => VN573_in0,
        Din1 => VN573_in1,
        Din2 => VN573_in2,
        Din3 => VN573_in3,
        Din4 => VN573_in4,
        Din5 => VN573_in5,
        VN2CN0_bit => VN_data_out(3438),
        VN2CN1_bit => VN_data_out(3439),
        VN2CN2_bit => VN_data_out(3440),
        VN2CN3_bit => VN_data_out(3441),
        VN2CN4_bit => VN_data_out(3442),
        VN2CN5_bit => VN_data_out(3443),
        VN2CN0_sign => VN_sign_out(3438),
        VN2CN1_sign => VN_sign_out(3439),
        VN2CN2_sign => VN_sign_out(3440),
        VN2CN3_sign => VN_sign_out(3441),
        VN2CN4_sign => VN_sign_out(3442),
        VN2CN5_sign => VN_sign_out(3443),
        codeword => codeword(573),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN574 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3449 downto 3444),
        Din0 => VN574_in0,
        Din1 => VN574_in1,
        Din2 => VN574_in2,
        Din3 => VN574_in3,
        Din4 => VN574_in4,
        Din5 => VN574_in5,
        VN2CN0_bit => VN_data_out(3444),
        VN2CN1_bit => VN_data_out(3445),
        VN2CN2_bit => VN_data_out(3446),
        VN2CN3_bit => VN_data_out(3447),
        VN2CN4_bit => VN_data_out(3448),
        VN2CN5_bit => VN_data_out(3449),
        VN2CN0_sign => VN_sign_out(3444),
        VN2CN1_sign => VN_sign_out(3445),
        VN2CN2_sign => VN_sign_out(3446),
        VN2CN3_sign => VN_sign_out(3447),
        VN2CN4_sign => VN_sign_out(3448),
        VN2CN5_sign => VN_sign_out(3449),
        codeword => codeword(574),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN575 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3455 downto 3450),
        Din0 => VN575_in0,
        Din1 => VN575_in1,
        Din2 => VN575_in2,
        Din3 => VN575_in3,
        Din4 => VN575_in4,
        Din5 => VN575_in5,
        VN2CN0_bit => VN_data_out(3450),
        VN2CN1_bit => VN_data_out(3451),
        VN2CN2_bit => VN_data_out(3452),
        VN2CN3_bit => VN_data_out(3453),
        VN2CN4_bit => VN_data_out(3454),
        VN2CN5_bit => VN_data_out(3455),
        VN2CN0_sign => VN_sign_out(3450),
        VN2CN1_sign => VN_sign_out(3451),
        VN2CN2_sign => VN_sign_out(3452),
        VN2CN3_sign => VN_sign_out(3453),
        VN2CN4_sign => VN_sign_out(3454),
        VN2CN5_sign => VN_sign_out(3455),
        codeword => codeword(575),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN576 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3461 downto 3456),
        Din0 => VN576_in0,
        Din1 => VN576_in1,
        Din2 => VN576_in2,
        Din3 => VN576_in3,
        Din4 => VN576_in4,
        Din5 => VN576_in5,
        VN2CN0_bit => VN_data_out(3456),
        VN2CN1_bit => VN_data_out(3457),
        VN2CN2_bit => VN_data_out(3458),
        VN2CN3_bit => VN_data_out(3459),
        VN2CN4_bit => VN_data_out(3460),
        VN2CN5_bit => VN_data_out(3461),
        VN2CN0_sign => VN_sign_out(3456),
        VN2CN1_sign => VN_sign_out(3457),
        VN2CN2_sign => VN_sign_out(3458),
        VN2CN3_sign => VN_sign_out(3459),
        VN2CN4_sign => VN_sign_out(3460),
        VN2CN5_sign => VN_sign_out(3461),
        codeword => codeword(576),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN577 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3467 downto 3462),
        Din0 => VN577_in0,
        Din1 => VN577_in1,
        Din2 => VN577_in2,
        Din3 => VN577_in3,
        Din4 => VN577_in4,
        Din5 => VN577_in5,
        VN2CN0_bit => VN_data_out(3462),
        VN2CN1_bit => VN_data_out(3463),
        VN2CN2_bit => VN_data_out(3464),
        VN2CN3_bit => VN_data_out(3465),
        VN2CN4_bit => VN_data_out(3466),
        VN2CN5_bit => VN_data_out(3467),
        VN2CN0_sign => VN_sign_out(3462),
        VN2CN1_sign => VN_sign_out(3463),
        VN2CN2_sign => VN_sign_out(3464),
        VN2CN3_sign => VN_sign_out(3465),
        VN2CN4_sign => VN_sign_out(3466),
        VN2CN5_sign => VN_sign_out(3467),
        codeword => codeword(577),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN578 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3473 downto 3468),
        Din0 => VN578_in0,
        Din1 => VN578_in1,
        Din2 => VN578_in2,
        Din3 => VN578_in3,
        Din4 => VN578_in4,
        Din5 => VN578_in5,
        VN2CN0_bit => VN_data_out(3468),
        VN2CN1_bit => VN_data_out(3469),
        VN2CN2_bit => VN_data_out(3470),
        VN2CN3_bit => VN_data_out(3471),
        VN2CN4_bit => VN_data_out(3472),
        VN2CN5_bit => VN_data_out(3473),
        VN2CN0_sign => VN_sign_out(3468),
        VN2CN1_sign => VN_sign_out(3469),
        VN2CN2_sign => VN_sign_out(3470),
        VN2CN3_sign => VN_sign_out(3471),
        VN2CN4_sign => VN_sign_out(3472),
        VN2CN5_sign => VN_sign_out(3473),
        codeword => codeword(578),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN579 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3479 downto 3474),
        Din0 => VN579_in0,
        Din1 => VN579_in1,
        Din2 => VN579_in2,
        Din3 => VN579_in3,
        Din4 => VN579_in4,
        Din5 => VN579_in5,
        VN2CN0_bit => VN_data_out(3474),
        VN2CN1_bit => VN_data_out(3475),
        VN2CN2_bit => VN_data_out(3476),
        VN2CN3_bit => VN_data_out(3477),
        VN2CN4_bit => VN_data_out(3478),
        VN2CN5_bit => VN_data_out(3479),
        VN2CN0_sign => VN_sign_out(3474),
        VN2CN1_sign => VN_sign_out(3475),
        VN2CN2_sign => VN_sign_out(3476),
        VN2CN3_sign => VN_sign_out(3477),
        VN2CN4_sign => VN_sign_out(3478),
        VN2CN5_sign => VN_sign_out(3479),
        codeword => codeword(579),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN580 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3485 downto 3480),
        Din0 => VN580_in0,
        Din1 => VN580_in1,
        Din2 => VN580_in2,
        Din3 => VN580_in3,
        Din4 => VN580_in4,
        Din5 => VN580_in5,
        VN2CN0_bit => VN_data_out(3480),
        VN2CN1_bit => VN_data_out(3481),
        VN2CN2_bit => VN_data_out(3482),
        VN2CN3_bit => VN_data_out(3483),
        VN2CN4_bit => VN_data_out(3484),
        VN2CN5_bit => VN_data_out(3485),
        VN2CN0_sign => VN_sign_out(3480),
        VN2CN1_sign => VN_sign_out(3481),
        VN2CN2_sign => VN_sign_out(3482),
        VN2CN3_sign => VN_sign_out(3483),
        VN2CN4_sign => VN_sign_out(3484),
        VN2CN5_sign => VN_sign_out(3485),
        codeword => codeword(580),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN581 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3491 downto 3486),
        Din0 => VN581_in0,
        Din1 => VN581_in1,
        Din2 => VN581_in2,
        Din3 => VN581_in3,
        Din4 => VN581_in4,
        Din5 => VN581_in5,
        VN2CN0_bit => VN_data_out(3486),
        VN2CN1_bit => VN_data_out(3487),
        VN2CN2_bit => VN_data_out(3488),
        VN2CN3_bit => VN_data_out(3489),
        VN2CN4_bit => VN_data_out(3490),
        VN2CN5_bit => VN_data_out(3491),
        VN2CN0_sign => VN_sign_out(3486),
        VN2CN1_sign => VN_sign_out(3487),
        VN2CN2_sign => VN_sign_out(3488),
        VN2CN3_sign => VN_sign_out(3489),
        VN2CN4_sign => VN_sign_out(3490),
        VN2CN5_sign => VN_sign_out(3491),
        codeword => codeword(581),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN582 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3497 downto 3492),
        Din0 => VN582_in0,
        Din1 => VN582_in1,
        Din2 => VN582_in2,
        Din3 => VN582_in3,
        Din4 => VN582_in4,
        Din5 => VN582_in5,
        VN2CN0_bit => VN_data_out(3492),
        VN2CN1_bit => VN_data_out(3493),
        VN2CN2_bit => VN_data_out(3494),
        VN2CN3_bit => VN_data_out(3495),
        VN2CN4_bit => VN_data_out(3496),
        VN2CN5_bit => VN_data_out(3497),
        VN2CN0_sign => VN_sign_out(3492),
        VN2CN1_sign => VN_sign_out(3493),
        VN2CN2_sign => VN_sign_out(3494),
        VN2CN3_sign => VN_sign_out(3495),
        VN2CN4_sign => VN_sign_out(3496),
        VN2CN5_sign => VN_sign_out(3497),
        codeword => codeword(582),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN583 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3503 downto 3498),
        Din0 => VN583_in0,
        Din1 => VN583_in1,
        Din2 => VN583_in2,
        Din3 => VN583_in3,
        Din4 => VN583_in4,
        Din5 => VN583_in5,
        VN2CN0_bit => VN_data_out(3498),
        VN2CN1_bit => VN_data_out(3499),
        VN2CN2_bit => VN_data_out(3500),
        VN2CN3_bit => VN_data_out(3501),
        VN2CN4_bit => VN_data_out(3502),
        VN2CN5_bit => VN_data_out(3503),
        VN2CN0_sign => VN_sign_out(3498),
        VN2CN1_sign => VN_sign_out(3499),
        VN2CN2_sign => VN_sign_out(3500),
        VN2CN3_sign => VN_sign_out(3501),
        VN2CN4_sign => VN_sign_out(3502),
        VN2CN5_sign => VN_sign_out(3503),
        codeword => codeword(583),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN584 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3509 downto 3504),
        Din0 => VN584_in0,
        Din1 => VN584_in1,
        Din2 => VN584_in2,
        Din3 => VN584_in3,
        Din4 => VN584_in4,
        Din5 => VN584_in5,
        VN2CN0_bit => VN_data_out(3504),
        VN2CN1_bit => VN_data_out(3505),
        VN2CN2_bit => VN_data_out(3506),
        VN2CN3_bit => VN_data_out(3507),
        VN2CN4_bit => VN_data_out(3508),
        VN2CN5_bit => VN_data_out(3509),
        VN2CN0_sign => VN_sign_out(3504),
        VN2CN1_sign => VN_sign_out(3505),
        VN2CN2_sign => VN_sign_out(3506),
        VN2CN3_sign => VN_sign_out(3507),
        VN2CN4_sign => VN_sign_out(3508),
        VN2CN5_sign => VN_sign_out(3509),
        codeword => codeword(584),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN585 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3515 downto 3510),
        Din0 => VN585_in0,
        Din1 => VN585_in1,
        Din2 => VN585_in2,
        Din3 => VN585_in3,
        Din4 => VN585_in4,
        Din5 => VN585_in5,
        VN2CN0_bit => VN_data_out(3510),
        VN2CN1_bit => VN_data_out(3511),
        VN2CN2_bit => VN_data_out(3512),
        VN2CN3_bit => VN_data_out(3513),
        VN2CN4_bit => VN_data_out(3514),
        VN2CN5_bit => VN_data_out(3515),
        VN2CN0_sign => VN_sign_out(3510),
        VN2CN1_sign => VN_sign_out(3511),
        VN2CN2_sign => VN_sign_out(3512),
        VN2CN3_sign => VN_sign_out(3513),
        VN2CN4_sign => VN_sign_out(3514),
        VN2CN5_sign => VN_sign_out(3515),
        codeword => codeword(585),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN586 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3521 downto 3516),
        Din0 => VN586_in0,
        Din1 => VN586_in1,
        Din2 => VN586_in2,
        Din3 => VN586_in3,
        Din4 => VN586_in4,
        Din5 => VN586_in5,
        VN2CN0_bit => VN_data_out(3516),
        VN2CN1_bit => VN_data_out(3517),
        VN2CN2_bit => VN_data_out(3518),
        VN2CN3_bit => VN_data_out(3519),
        VN2CN4_bit => VN_data_out(3520),
        VN2CN5_bit => VN_data_out(3521),
        VN2CN0_sign => VN_sign_out(3516),
        VN2CN1_sign => VN_sign_out(3517),
        VN2CN2_sign => VN_sign_out(3518),
        VN2CN3_sign => VN_sign_out(3519),
        VN2CN4_sign => VN_sign_out(3520),
        VN2CN5_sign => VN_sign_out(3521),
        codeword => codeword(586),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN587 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3527 downto 3522),
        Din0 => VN587_in0,
        Din1 => VN587_in1,
        Din2 => VN587_in2,
        Din3 => VN587_in3,
        Din4 => VN587_in4,
        Din5 => VN587_in5,
        VN2CN0_bit => VN_data_out(3522),
        VN2CN1_bit => VN_data_out(3523),
        VN2CN2_bit => VN_data_out(3524),
        VN2CN3_bit => VN_data_out(3525),
        VN2CN4_bit => VN_data_out(3526),
        VN2CN5_bit => VN_data_out(3527),
        VN2CN0_sign => VN_sign_out(3522),
        VN2CN1_sign => VN_sign_out(3523),
        VN2CN2_sign => VN_sign_out(3524),
        VN2CN3_sign => VN_sign_out(3525),
        VN2CN4_sign => VN_sign_out(3526),
        VN2CN5_sign => VN_sign_out(3527),
        codeword => codeword(587),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN588 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3533 downto 3528),
        Din0 => VN588_in0,
        Din1 => VN588_in1,
        Din2 => VN588_in2,
        Din3 => VN588_in3,
        Din4 => VN588_in4,
        Din5 => VN588_in5,
        VN2CN0_bit => VN_data_out(3528),
        VN2CN1_bit => VN_data_out(3529),
        VN2CN2_bit => VN_data_out(3530),
        VN2CN3_bit => VN_data_out(3531),
        VN2CN4_bit => VN_data_out(3532),
        VN2CN5_bit => VN_data_out(3533),
        VN2CN0_sign => VN_sign_out(3528),
        VN2CN1_sign => VN_sign_out(3529),
        VN2CN2_sign => VN_sign_out(3530),
        VN2CN3_sign => VN_sign_out(3531),
        VN2CN4_sign => VN_sign_out(3532),
        VN2CN5_sign => VN_sign_out(3533),
        codeword => codeword(588),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN589 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3539 downto 3534),
        Din0 => VN589_in0,
        Din1 => VN589_in1,
        Din2 => VN589_in2,
        Din3 => VN589_in3,
        Din4 => VN589_in4,
        Din5 => VN589_in5,
        VN2CN0_bit => VN_data_out(3534),
        VN2CN1_bit => VN_data_out(3535),
        VN2CN2_bit => VN_data_out(3536),
        VN2CN3_bit => VN_data_out(3537),
        VN2CN4_bit => VN_data_out(3538),
        VN2CN5_bit => VN_data_out(3539),
        VN2CN0_sign => VN_sign_out(3534),
        VN2CN1_sign => VN_sign_out(3535),
        VN2CN2_sign => VN_sign_out(3536),
        VN2CN3_sign => VN_sign_out(3537),
        VN2CN4_sign => VN_sign_out(3538),
        VN2CN5_sign => VN_sign_out(3539),
        codeword => codeword(589),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN590 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3545 downto 3540),
        Din0 => VN590_in0,
        Din1 => VN590_in1,
        Din2 => VN590_in2,
        Din3 => VN590_in3,
        Din4 => VN590_in4,
        Din5 => VN590_in5,
        VN2CN0_bit => VN_data_out(3540),
        VN2CN1_bit => VN_data_out(3541),
        VN2CN2_bit => VN_data_out(3542),
        VN2CN3_bit => VN_data_out(3543),
        VN2CN4_bit => VN_data_out(3544),
        VN2CN5_bit => VN_data_out(3545),
        VN2CN0_sign => VN_sign_out(3540),
        VN2CN1_sign => VN_sign_out(3541),
        VN2CN2_sign => VN_sign_out(3542),
        VN2CN3_sign => VN_sign_out(3543),
        VN2CN4_sign => VN_sign_out(3544),
        VN2CN5_sign => VN_sign_out(3545),
        codeword => codeword(590),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN591 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3551 downto 3546),
        Din0 => VN591_in0,
        Din1 => VN591_in1,
        Din2 => VN591_in2,
        Din3 => VN591_in3,
        Din4 => VN591_in4,
        Din5 => VN591_in5,
        VN2CN0_bit => VN_data_out(3546),
        VN2CN1_bit => VN_data_out(3547),
        VN2CN2_bit => VN_data_out(3548),
        VN2CN3_bit => VN_data_out(3549),
        VN2CN4_bit => VN_data_out(3550),
        VN2CN5_bit => VN_data_out(3551),
        VN2CN0_sign => VN_sign_out(3546),
        VN2CN1_sign => VN_sign_out(3547),
        VN2CN2_sign => VN_sign_out(3548),
        VN2CN3_sign => VN_sign_out(3549),
        VN2CN4_sign => VN_sign_out(3550),
        VN2CN5_sign => VN_sign_out(3551),
        codeword => codeword(591),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN592 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3557 downto 3552),
        Din0 => VN592_in0,
        Din1 => VN592_in1,
        Din2 => VN592_in2,
        Din3 => VN592_in3,
        Din4 => VN592_in4,
        Din5 => VN592_in5,
        VN2CN0_bit => VN_data_out(3552),
        VN2CN1_bit => VN_data_out(3553),
        VN2CN2_bit => VN_data_out(3554),
        VN2CN3_bit => VN_data_out(3555),
        VN2CN4_bit => VN_data_out(3556),
        VN2CN5_bit => VN_data_out(3557),
        VN2CN0_sign => VN_sign_out(3552),
        VN2CN1_sign => VN_sign_out(3553),
        VN2CN2_sign => VN_sign_out(3554),
        VN2CN3_sign => VN_sign_out(3555),
        VN2CN4_sign => VN_sign_out(3556),
        VN2CN5_sign => VN_sign_out(3557),
        codeword => codeword(592),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN593 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3563 downto 3558),
        Din0 => VN593_in0,
        Din1 => VN593_in1,
        Din2 => VN593_in2,
        Din3 => VN593_in3,
        Din4 => VN593_in4,
        Din5 => VN593_in5,
        VN2CN0_bit => VN_data_out(3558),
        VN2CN1_bit => VN_data_out(3559),
        VN2CN2_bit => VN_data_out(3560),
        VN2CN3_bit => VN_data_out(3561),
        VN2CN4_bit => VN_data_out(3562),
        VN2CN5_bit => VN_data_out(3563),
        VN2CN0_sign => VN_sign_out(3558),
        VN2CN1_sign => VN_sign_out(3559),
        VN2CN2_sign => VN_sign_out(3560),
        VN2CN3_sign => VN_sign_out(3561),
        VN2CN4_sign => VN_sign_out(3562),
        VN2CN5_sign => VN_sign_out(3563),
        codeword => codeword(593),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN594 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3569 downto 3564),
        Din0 => VN594_in0,
        Din1 => VN594_in1,
        Din2 => VN594_in2,
        Din3 => VN594_in3,
        Din4 => VN594_in4,
        Din5 => VN594_in5,
        VN2CN0_bit => VN_data_out(3564),
        VN2CN1_bit => VN_data_out(3565),
        VN2CN2_bit => VN_data_out(3566),
        VN2CN3_bit => VN_data_out(3567),
        VN2CN4_bit => VN_data_out(3568),
        VN2CN5_bit => VN_data_out(3569),
        VN2CN0_sign => VN_sign_out(3564),
        VN2CN1_sign => VN_sign_out(3565),
        VN2CN2_sign => VN_sign_out(3566),
        VN2CN3_sign => VN_sign_out(3567),
        VN2CN4_sign => VN_sign_out(3568),
        VN2CN5_sign => VN_sign_out(3569),
        codeword => codeword(594),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN595 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3575 downto 3570),
        Din0 => VN595_in0,
        Din1 => VN595_in1,
        Din2 => VN595_in2,
        Din3 => VN595_in3,
        Din4 => VN595_in4,
        Din5 => VN595_in5,
        VN2CN0_bit => VN_data_out(3570),
        VN2CN1_bit => VN_data_out(3571),
        VN2CN2_bit => VN_data_out(3572),
        VN2CN3_bit => VN_data_out(3573),
        VN2CN4_bit => VN_data_out(3574),
        VN2CN5_bit => VN_data_out(3575),
        VN2CN0_sign => VN_sign_out(3570),
        VN2CN1_sign => VN_sign_out(3571),
        VN2CN2_sign => VN_sign_out(3572),
        VN2CN3_sign => VN_sign_out(3573),
        VN2CN4_sign => VN_sign_out(3574),
        VN2CN5_sign => VN_sign_out(3575),
        codeword => codeword(595),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN596 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3581 downto 3576),
        Din0 => VN596_in0,
        Din1 => VN596_in1,
        Din2 => VN596_in2,
        Din3 => VN596_in3,
        Din4 => VN596_in4,
        Din5 => VN596_in5,
        VN2CN0_bit => VN_data_out(3576),
        VN2CN1_bit => VN_data_out(3577),
        VN2CN2_bit => VN_data_out(3578),
        VN2CN3_bit => VN_data_out(3579),
        VN2CN4_bit => VN_data_out(3580),
        VN2CN5_bit => VN_data_out(3581),
        VN2CN0_sign => VN_sign_out(3576),
        VN2CN1_sign => VN_sign_out(3577),
        VN2CN2_sign => VN_sign_out(3578),
        VN2CN3_sign => VN_sign_out(3579),
        VN2CN4_sign => VN_sign_out(3580),
        VN2CN5_sign => VN_sign_out(3581),
        codeword => codeword(596),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN597 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3587 downto 3582),
        Din0 => VN597_in0,
        Din1 => VN597_in1,
        Din2 => VN597_in2,
        Din3 => VN597_in3,
        Din4 => VN597_in4,
        Din5 => VN597_in5,
        VN2CN0_bit => VN_data_out(3582),
        VN2CN1_bit => VN_data_out(3583),
        VN2CN2_bit => VN_data_out(3584),
        VN2CN3_bit => VN_data_out(3585),
        VN2CN4_bit => VN_data_out(3586),
        VN2CN5_bit => VN_data_out(3587),
        VN2CN0_sign => VN_sign_out(3582),
        VN2CN1_sign => VN_sign_out(3583),
        VN2CN2_sign => VN_sign_out(3584),
        VN2CN3_sign => VN_sign_out(3585),
        VN2CN4_sign => VN_sign_out(3586),
        VN2CN5_sign => VN_sign_out(3587),
        codeword => codeword(597),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN598 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3593 downto 3588),
        Din0 => VN598_in0,
        Din1 => VN598_in1,
        Din2 => VN598_in2,
        Din3 => VN598_in3,
        Din4 => VN598_in4,
        Din5 => VN598_in5,
        VN2CN0_bit => VN_data_out(3588),
        VN2CN1_bit => VN_data_out(3589),
        VN2CN2_bit => VN_data_out(3590),
        VN2CN3_bit => VN_data_out(3591),
        VN2CN4_bit => VN_data_out(3592),
        VN2CN5_bit => VN_data_out(3593),
        VN2CN0_sign => VN_sign_out(3588),
        VN2CN1_sign => VN_sign_out(3589),
        VN2CN2_sign => VN_sign_out(3590),
        VN2CN3_sign => VN_sign_out(3591),
        VN2CN4_sign => VN_sign_out(3592),
        VN2CN5_sign => VN_sign_out(3593),
        codeword => codeword(598),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN599 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3599 downto 3594),
        Din0 => VN599_in0,
        Din1 => VN599_in1,
        Din2 => VN599_in2,
        Din3 => VN599_in3,
        Din4 => VN599_in4,
        Din5 => VN599_in5,
        VN2CN0_bit => VN_data_out(3594),
        VN2CN1_bit => VN_data_out(3595),
        VN2CN2_bit => VN_data_out(3596),
        VN2CN3_bit => VN_data_out(3597),
        VN2CN4_bit => VN_data_out(3598),
        VN2CN5_bit => VN_data_out(3599),
        VN2CN0_sign => VN_sign_out(3594),
        VN2CN1_sign => VN_sign_out(3595),
        VN2CN2_sign => VN_sign_out(3596),
        VN2CN3_sign => VN_sign_out(3597),
        VN2CN4_sign => VN_sign_out(3598),
        VN2CN5_sign => VN_sign_out(3599),
        codeword => codeword(599),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN600 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3605 downto 3600),
        Din0 => VN600_in0,
        Din1 => VN600_in1,
        Din2 => VN600_in2,
        Din3 => VN600_in3,
        Din4 => VN600_in4,
        Din5 => VN600_in5,
        VN2CN0_bit => VN_data_out(3600),
        VN2CN1_bit => VN_data_out(3601),
        VN2CN2_bit => VN_data_out(3602),
        VN2CN3_bit => VN_data_out(3603),
        VN2CN4_bit => VN_data_out(3604),
        VN2CN5_bit => VN_data_out(3605),
        VN2CN0_sign => VN_sign_out(3600),
        VN2CN1_sign => VN_sign_out(3601),
        VN2CN2_sign => VN_sign_out(3602),
        VN2CN3_sign => VN_sign_out(3603),
        VN2CN4_sign => VN_sign_out(3604),
        VN2CN5_sign => VN_sign_out(3605),
        codeword => codeword(600),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN601 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3611 downto 3606),
        Din0 => VN601_in0,
        Din1 => VN601_in1,
        Din2 => VN601_in2,
        Din3 => VN601_in3,
        Din4 => VN601_in4,
        Din5 => VN601_in5,
        VN2CN0_bit => VN_data_out(3606),
        VN2CN1_bit => VN_data_out(3607),
        VN2CN2_bit => VN_data_out(3608),
        VN2CN3_bit => VN_data_out(3609),
        VN2CN4_bit => VN_data_out(3610),
        VN2CN5_bit => VN_data_out(3611),
        VN2CN0_sign => VN_sign_out(3606),
        VN2CN1_sign => VN_sign_out(3607),
        VN2CN2_sign => VN_sign_out(3608),
        VN2CN3_sign => VN_sign_out(3609),
        VN2CN4_sign => VN_sign_out(3610),
        VN2CN5_sign => VN_sign_out(3611),
        codeword => codeword(601),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN602 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3617 downto 3612),
        Din0 => VN602_in0,
        Din1 => VN602_in1,
        Din2 => VN602_in2,
        Din3 => VN602_in3,
        Din4 => VN602_in4,
        Din5 => VN602_in5,
        VN2CN0_bit => VN_data_out(3612),
        VN2CN1_bit => VN_data_out(3613),
        VN2CN2_bit => VN_data_out(3614),
        VN2CN3_bit => VN_data_out(3615),
        VN2CN4_bit => VN_data_out(3616),
        VN2CN5_bit => VN_data_out(3617),
        VN2CN0_sign => VN_sign_out(3612),
        VN2CN1_sign => VN_sign_out(3613),
        VN2CN2_sign => VN_sign_out(3614),
        VN2CN3_sign => VN_sign_out(3615),
        VN2CN4_sign => VN_sign_out(3616),
        VN2CN5_sign => VN_sign_out(3617),
        codeword => codeword(602),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN603 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3623 downto 3618),
        Din0 => VN603_in0,
        Din1 => VN603_in1,
        Din2 => VN603_in2,
        Din3 => VN603_in3,
        Din4 => VN603_in4,
        Din5 => VN603_in5,
        VN2CN0_bit => VN_data_out(3618),
        VN2CN1_bit => VN_data_out(3619),
        VN2CN2_bit => VN_data_out(3620),
        VN2CN3_bit => VN_data_out(3621),
        VN2CN4_bit => VN_data_out(3622),
        VN2CN5_bit => VN_data_out(3623),
        VN2CN0_sign => VN_sign_out(3618),
        VN2CN1_sign => VN_sign_out(3619),
        VN2CN2_sign => VN_sign_out(3620),
        VN2CN3_sign => VN_sign_out(3621),
        VN2CN4_sign => VN_sign_out(3622),
        VN2CN5_sign => VN_sign_out(3623),
        codeword => codeword(603),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN604 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3629 downto 3624),
        Din0 => VN604_in0,
        Din1 => VN604_in1,
        Din2 => VN604_in2,
        Din3 => VN604_in3,
        Din4 => VN604_in4,
        Din5 => VN604_in5,
        VN2CN0_bit => VN_data_out(3624),
        VN2CN1_bit => VN_data_out(3625),
        VN2CN2_bit => VN_data_out(3626),
        VN2CN3_bit => VN_data_out(3627),
        VN2CN4_bit => VN_data_out(3628),
        VN2CN5_bit => VN_data_out(3629),
        VN2CN0_sign => VN_sign_out(3624),
        VN2CN1_sign => VN_sign_out(3625),
        VN2CN2_sign => VN_sign_out(3626),
        VN2CN3_sign => VN_sign_out(3627),
        VN2CN4_sign => VN_sign_out(3628),
        VN2CN5_sign => VN_sign_out(3629),
        codeword => codeword(604),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN605 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3635 downto 3630),
        Din0 => VN605_in0,
        Din1 => VN605_in1,
        Din2 => VN605_in2,
        Din3 => VN605_in3,
        Din4 => VN605_in4,
        Din5 => VN605_in5,
        VN2CN0_bit => VN_data_out(3630),
        VN2CN1_bit => VN_data_out(3631),
        VN2CN2_bit => VN_data_out(3632),
        VN2CN3_bit => VN_data_out(3633),
        VN2CN4_bit => VN_data_out(3634),
        VN2CN5_bit => VN_data_out(3635),
        VN2CN0_sign => VN_sign_out(3630),
        VN2CN1_sign => VN_sign_out(3631),
        VN2CN2_sign => VN_sign_out(3632),
        VN2CN3_sign => VN_sign_out(3633),
        VN2CN4_sign => VN_sign_out(3634),
        VN2CN5_sign => VN_sign_out(3635),
        codeword => codeword(605),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN606 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3641 downto 3636),
        Din0 => VN606_in0,
        Din1 => VN606_in1,
        Din2 => VN606_in2,
        Din3 => VN606_in3,
        Din4 => VN606_in4,
        Din5 => VN606_in5,
        VN2CN0_bit => VN_data_out(3636),
        VN2CN1_bit => VN_data_out(3637),
        VN2CN2_bit => VN_data_out(3638),
        VN2CN3_bit => VN_data_out(3639),
        VN2CN4_bit => VN_data_out(3640),
        VN2CN5_bit => VN_data_out(3641),
        VN2CN0_sign => VN_sign_out(3636),
        VN2CN1_sign => VN_sign_out(3637),
        VN2CN2_sign => VN_sign_out(3638),
        VN2CN3_sign => VN_sign_out(3639),
        VN2CN4_sign => VN_sign_out(3640),
        VN2CN5_sign => VN_sign_out(3641),
        codeword => codeword(606),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN607 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3647 downto 3642),
        Din0 => VN607_in0,
        Din1 => VN607_in1,
        Din2 => VN607_in2,
        Din3 => VN607_in3,
        Din4 => VN607_in4,
        Din5 => VN607_in5,
        VN2CN0_bit => VN_data_out(3642),
        VN2CN1_bit => VN_data_out(3643),
        VN2CN2_bit => VN_data_out(3644),
        VN2CN3_bit => VN_data_out(3645),
        VN2CN4_bit => VN_data_out(3646),
        VN2CN5_bit => VN_data_out(3647),
        VN2CN0_sign => VN_sign_out(3642),
        VN2CN1_sign => VN_sign_out(3643),
        VN2CN2_sign => VN_sign_out(3644),
        VN2CN3_sign => VN_sign_out(3645),
        VN2CN4_sign => VN_sign_out(3646),
        VN2CN5_sign => VN_sign_out(3647),
        codeword => codeword(607),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN608 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3653 downto 3648),
        Din0 => VN608_in0,
        Din1 => VN608_in1,
        Din2 => VN608_in2,
        Din3 => VN608_in3,
        Din4 => VN608_in4,
        Din5 => VN608_in5,
        VN2CN0_bit => VN_data_out(3648),
        VN2CN1_bit => VN_data_out(3649),
        VN2CN2_bit => VN_data_out(3650),
        VN2CN3_bit => VN_data_out(3651),
        VN2CN4_bit => VN_data_out(3652),
        VN2CN5_bit => VN_data_out(3653),
        VN2CN0_sign => VN_sign_out(3648),
        VN2CN1_sign => VN_sign_out(3649),
        VN2CN2_sign => VN_sign_out(3650),
        VN2CN3_sign => VN_sign_out(3651),
        VN2CN4_sign => VN_sign_out(3652),
        VN2CN5_sign => VN_sign_out(3653),
        codeword => codeword(608),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN609 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3659 downto 3654),
        Din0 => VN609_in0,
        Din1 => VN609_in1,
        Din2 => VN609_in2,
        Din3 => VN609_in3,
        Din4 => VN609_in4,
        Din5 => VN609_in5,
        VN2CN0_bit => VN_data_out(3654),
        VN2CN1_bit => VN_data_out(3655),
        VN2CN2_bit => VN_data_out(3656),
        VN2CN3_bit => VN_data_out(3657),
        VN2CN4_bit => VN_data_out(3658),
        VN2CN5_bit => VN_data_out(3659),
        VN2CN0_sign => VN_sign_out(3654),
        VN2CN1_sign => VN_sign_out(3655),
        VN2CN2_sign => VN_sign_out(3656),
        VN2CN3_sign => VN_sign_out(3657),
        VN2CN4_sign => VN_sign_out(3658),
        VN2CN5_sign => VN_sign_out(3659),
        codeword => codeword(609),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN610 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3665 downto 3660),
        Din0 => VN610_in0,
        Din1 => VN610_in1,
        Din2 => VN610_in2,
        Din3 => VN610_in3,
        Din4 => VN610_in4,
        Din5 => VN610_in5,
        VN2CN0_bit => VN_data_out(3660),
        VN2CN1_bit => VN_data_out(3661),
        VN2CN2_bit => VN_data_out(3662),
        VN2CN3_bit => VN_data_out(3663),
        VN2CN4_bit => VN_data_out(3664),
        VN2CN5_bit => VN_data_out(3665),
        VN2CN0_sign => VN_sign_out(3660),
        VN2CN1_sign => VN_sign_out(3661),
        VN2CN2_sign => VN_sign_out(3662),
        VN2CN3_sign => VN_sign_out(3663),
        VN2CN4_sign => VN_sign_out(3664),
        VN2CN5_sign => VN_sign_out(3665),
        codeword => codeword(610),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN611 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3671 downto 3666),
        Din0 => VN611_in0,
        Din1 => VN611_in1,
        Din2 => VN611_in2,
        Din3 => VN611_in3,
        Din4 => VN611_in4,
        Din5 => VN611_in5,
        VN2CN0_bit => VN_data_out(3666),
        VN2CN1_bit => VN_data_out(3667),
        VN2CN2_bit => VN_data_out(3668),
        VN2CN3_bit => VN_data_out(3669),
        VN2CN4_bit => VN_data_out(3670),
        VN2CN5_bit => VN_data_out(3671),
        VN2CN0_sign => VN_sign_out(3666),
        VN2CN1_sign => VN_sign_out(3667),
        VN2CN2_sign => VN_sign_out(3668),
        VN2CN3_sign => VN_sign_out(3669),
        VN2CN4_sign => VN_sign_out(3670),
        VN2CN5_sign => VN_sign_out(3671),
        codeword => codeword(611),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN612 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3677 downto 3672),
        Din0 => VN612_in0,
        Din1 => VN612_in1,
        Din2 => VN612_in2,
        Din3 => VN612_in3,
        Din4 => VN612_in4,
        Din5 => VN612_in5,
        VN2CN0_bit => VN_data_out(3672),
        VN2CN1_bit => VN_data_out(3673),
        VN2CN2_bit => VN_data_out(3674),
        VN2CN3_bit => VN_data_out(3675),
        VN2CN4_bit => VN_data_out(3676),
        VN2CN5_bit => VN_data_out(3677),
        VN2CN0_sign => VN_sign_out(3672),
        VN2CN1_sign => VN_sign_out(3673),
        VN2CN2_sign => VN_sign_out(3674),
        VN2CN3_sign => VN_sign_out(3675),
        VN2CN4_sign => VN_sign_out(3676),
        VN2CN5_sign => VN_sign_out(3677),
        codeword => codeword(612),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN613 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3683 downto 3678),
        Din0 => VN613_in0,
        Din1 => VN613_in1,
        Din2 => VN613_in2,
        Din3 => VN613_in3,
        Din4 => VN613_in4,
        Din5 => VN613_in5,
        VN2CN0_bit => VN_data_out(3678),
        VN2CN1_bit => VN_data_out(3679),
        VN2CN2_bit => VN_data_out(3680),
        VN2CN3_bit => VN_data_out(3681),
        VN2CN4_bit => VN_data_out(3682),
        VN2CN5_bit => VN_data_out(3683),
        VN2CN0_sign => VN_sign_out(3678),
        VN2CN1_sign => VN_sign_out(3679),
        VN2CN2_sign => VN_sign_out(3680),
        VN2CN3_sign => VN_sign_out(3681),
        VN2CN4_sign => VN_sign_out(3682),
        VN2CN5_sign => VN_sign_out(3683),
        codeword => codeword(613),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN614 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3689 downto 3684),
        Din0 => VN614_in0,
        Din1 => VN614_in1,
        Din2 => VN614_in2,
        Din3 => VN614_in3,
        Din4 => VN614_in4,
        Din5 => VN614_in5,
        VN2CN0_bit => VN_data_out(3684),
        VN2CN1_bit => VN_data_out(3685),
        VN2CN2_bit => VN_data_out(3686),
        VN2CN3_bit => VN_data_out(3687),
        VN2CN4_bit => VN_data_out(3688),
        VN2CN5_bit => VN_data_out(3689),
        VN2CN0_sign => VN_sign_out(3684),
        VN2CN1_sign => VN_sign_out(3685),
        VN2CN2_sign => VN_sign_out(3686),
        VN2CN3_sign => VN_sign_out(3687),
        VN2CN4_sign => VN_sign_out(3688),
        VN2CN5_sign => VN_sign_out(3689),
        codeword => codeword(614),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN615 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3695 downto 3690),
        Din0 => VN615_in0,
        Din1 => VN615_in1,
        Din2 => VN615_in2,
        Din3 => VN615_in3,
        Din4 => VN615_in4,
        Din5 => VN615_in5,
        VN2CN0_bit => VN_data_out(3690),
        VN2CN1_bit => VN_data_out(3691),
        VN2CN2_bit => VN_data_out(3692),
        VN2CN3_bit => VN_data_out(3693),
        VN2CN4_bit => VN_data_out(3694),
        VN2CN5_bit => VN_data_out(3695),
        VN2CN0_sign => VN_sign_out(3690),
        VN2CN1_sign => VN_sign_out(3691),
        VN2CN2_sign => VN_sign_out(3692),
        VN2CN3_sign => VN_sign_out(3693),
        VN2CN4_sign => VN_sign_out(3694),
        VN2CN5_sign => VN_sign_out(3695),
        codeword => codeword(615),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN616 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3701 downto 3696),
        Din0 => VN616_in0,
        Din1 => VN616_in1,
        Din2 => VN616_in2,
        Din3 => VN616_in3,
        Din4 => VN616_in4,
        Din5 => VN616_in5,
        VN2CN0_bit => VN_data_out(3696),
        VN2CN1_bit => VN_data_out(3697),
        VN2CN2_bit => VN_data_out(3698),
        VN2CN3_bit => VN_data_out(3699),
        VN2CN4_bit => VN_data_out(3700),
        VN2CN5_bit => VN_data_out(3701),
        VN2CN0_sign => VN_sign_out(3696),
        VN2CN1_sign => VN_sign_out(3697),
        VN2CN2_sign => VN_sign_out(3698),
        VN2CN3_sign => VN_sign_out(3699),
        VN2CN4_sign => VN_sign_out(3700),
        VN2CN5_sign => VN_sign_out(3701),
        codeword => codeword(616),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN617 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3707 downto 3702),
        Din0 => VN617_in0,
        Din1 => VN617_in1,
        Din2 => VN617_in2,
        Din3 => VN617_in3,
        Din4 => VN617_in4,
        Din5 => VN617_in5,
        VN2CN0_bit => VN_data_out(3702),
        VN2CN1_bit => VN_data_out(3703),
        VN2CN2_bit => VN_data_out(3704),
        VN2CN3_bit => VN_data_out(3705),
        VN2CN4_bit => VN_data_out(3706),
        VN2CN5_bit => VN_data_out(3707),
        VN2CN0_sign => VN_sign_out(3702),
        VN2CN1_sign => VN_sign_out(3703),
        VN2CN2_sign => VN_sign_out(3704),
        VN2CN3_sign => VN_sign_out(3705),
        VN2CN4_sign => VN_sign_out(3706),
        VN2CN5_sign => VN_sign_out(3707),
        codeword => codeword(617),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN618 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3713 downto 3708),
        Din0 => VN618_in0,
        Din1 => VN618_in1,
        Din2 => VN618_in2,
        Din3 => VN618_in3,
        Din4 => VN618_in4,
        Din5 => VN618_in5,
        VN2CN0_bit => VN_data_out(3708),
        VN2CN1_bit => VN_data_out(3709),
        VN2CN2_bit => VN_data_out(3710),
        VN2CN3_bit => VN_data_out(3711),
        VN2CN4_bit => VN_data_out(3712),
        VN2CN5_bit => VN_data_out(3713),
        VN2CN0_sign => VN_sign_out(3708),
        VN2CN1_sign => VN_sign_out(3709),
        VN2CN2_sign => VN_sign_out(3710),
        VN2CN3_sign => VN_sign_out(3711),
        VN2CN4_sign => VN_sign_out(3712),
        VN2CN5_sign => VN_sign_out(3713),
        codeword => codeword(618),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN619 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3719 downto 3714),
        Din0 => VN619_in0,
        Din1 => VN619_in1,
        Din2 => VN619_in2,
        Din3 => VN619_in3,
        Din4 => VN619_in4,
        Din5 => VN619_in5,
        VN2CN0_bit => VN_data_out(3714),
        VN2CN1_bit => VN_data_out(3715),
        VN2CN2_bit => VN_data_out(3716),
        VN2CN3_bit => VN_data_out(3717),
        VN2CN4_bit => VN_data_out(3718),
        VN2CN5_bit => VN_data_out(3719),
        VN2CN0_sign => VN_sign_out(3714),
        VN2CN1_sign => VN_sign_out(3715),
        VN2CN2_sign => VN_sign_out(3716),
        VN2CN3_sign => VN_sign_out(3717),
        VN2CN4_sign => VN_sign_out(3718),
        VN2CN5_sign => VN_sign_out(3719),
        codeword => codeword(619),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN620 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3725 downto 3720),
        Din0 => VN620_in0,
        Din1 => VN620_in1,
        Din2 => VN620_in2,
        Din3 => VN620_in3,
        Din4 => VN620_in4,
        Din5 => VN620_in5,
        VN2CN0_bit => VN_data_out(3720),
        VN2CN1_bit => VN_data_out(3721),
        VN2CN2_bit => VN_data_out(3722),
        VN2CN3_bit => VN_data_out(3723),
        VN2CN4_bit => VN_data_out(3724),
        VN2CN5_bit => VN_data_out(3725),
        VN2CN0_sign => VN_sign_out(3720),
        VN2CN1_sign => VN_sign_out(3721),
        VN2CN2_sign => VN_sign_out(3722),
        VN2CN3_sign => VN_sign_out(3723),
        VN2CN4_sign => VN_sign_out(3724),
        VN2CN5_sign => VN_sign_out(3725),
        codeword => codeword(620),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN621 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3731 downto 3726),
        Din0 => VN621_in0,
        Din1 => VN621_in1,
        Din2 => VN621_in2,
        Din3 => VN621_in3,
        Din4 => VN621_in4,
        Din5 => VN621_in5,
        VN2CN0_bit => VN_data_out(3726),
        VN2CN1_bit => VN_data_out(3727),
        VN2CN2_bit => VN_data_out(3728),
        VN2CN3_bit => VN_data_out(3729),
        VN2CN4_bit => VN_data_out(3730),
        VN2CN5_bit => VN_data_out(3731),
        VN2CN0_sign => VN_sign_out(3726),
        VN2CN1_sign => VN_sign_out(3727),
        VN2CN2_sign => VN_sign_out(3728),
        VN2CN3_sign => VN_sign_out(3729),
        VN2CN4_sign => VN_sign_out(3730),
        VN2CN5_sign => VN_sign_out(3731),
        codeword => codeword(621),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN622 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3737 downto 3732),
        Din0 => VN622_in0,
        Din1 => VN622_in1,
        Din2 => VN622_in2,
        Din3 => VN622_in3,
        Din4 => VN622_in4,
        Din5 => VN622_in5,
        VN2CN0_bit => VN_data_out(3732),
        VN2CN1_bit => VN_data_out(3733),
        VN2CN2_bit => VN_data_out(3734),
        VN2CN3_bit => VN_data_out(3735),
        VN2CN4_bit => VN_data_out(3736),
        VN2CN5_bit => VN_data_out(3737),
        VN2CN0_sign => VN_sign_out(3732),
        VN2CN1_sign => VN_sign_out(3733),
        VN2CN2_sign => VN_sign_out(3734),
        VN2CN3_sign => VN_sign_out(3735),
        VN2CN4_sign => VN_sign_out(3736),
        VN2CN5_sign => VN_sign_out(3737),
        codeword => codeword(622),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN623 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3743 downto 3738),
        Din0 => VN623_in0,
        Din1 => VN623_in1,
        Din2 => VN623_in2,
        Din3 => VN623_in3,
        Din4 => VN623_in4,
        Din5 => VN623_in5,
        VN2CN0_bit => VN_data_out(3738),
        VN2CN1_bit => VN_data_out(3739),
        VN2CN2_bit => VN_data_out(3740),
        VN2CN3_bit => VN_data_out(3741),
        VN2CN4_bit => VN_data_out(3742),
        VN2CN5_bit => VN_data_out(3743),
        VN2CN0_sign => VN_sign_out(3738),
        VN2CN1_sign => VN_sign_out(3739),
        VN2CN2_sign => VN_sign_out(3740),
        VN2CN3_sign => VN_sign_out(3741),
        VN2CN4_sign => VN_sign_out(3742),
        VN2CN5_sign => VN_sign_out(3743),
        codeword => codeword(623),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN624 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3749 downto 3744),
        Din0 => VN624_in0,
        Din1 => VN624_in1,
        Din2 => VN624_in2,
        Din3 => VN624_in3,
        Din4 => VN624_in4,
        Din5 => VN624_in5,
        VN2CN0_bit => VN_data_out(3744),
        VN2CN1_bit => VN_data_out(3745),
        VN2CN2_bit => VN_data_out(3746),
        VN2CN3_bit => VN_data_out(3747),
        VN2CN4_bit => VN_data_out(3748),
        VN2CN5_bit => VN_data_out(3749),
        VN2CN0_sign => VN_sign_out(3744),
        VN2CN1_sign => VN_sign_out(3745),
        VN2CN2_sign => VN_sign_out(3746),
        VN2CN3_sign => VN_sign_out(3747),
        VN2CN4_sign => VN_sign_out(3748),
        VN2CN5_sign => VN_sign_out(3749),
        codeword => codeword(624),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN625 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3755 downto 3750),
        Din0 => VN625_in0,
        Din1 => VN625_in1,
        Din2 => VN625_in2,
        Din3 => VN625_in3,
        Din4 => VN625_in4,
        Din5 => VN625_in5,
        VN2CN0_bit => VN_data_out(3750),
        VN2CN1_bit => VN_data_out(3751),
        VN2CN2_bit => VN_data_out(3752),
        VN2CN3_bit => VN_data_out(3753),
        VN2CN4_bit => VN_data_out(3754),
        VN2CN5_bit => VN_data_out(3755),
        VN2CN0_sign => VN_sign_out(3750),
        VN2CN1_sign => VN_sign_out(3751),
        VN2CN2_sign => VN_sign_out(3752),
        VN2CN3_sign => VN_sign_out(3753),
        VN2CN4_sign => VN_sign_out(3754),
        VN2CN5_sign => VN_sign_out(3755),
        codeword => codeword(625),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN626 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3761 downto 3756),
        Din0 => VN626_in0,
        Din1 => VN626_in1,
        Din2 => VN626_in2,
        Din3 => VN626_in3,
        Din4 => VN626_in4,
        Din5 => VN626_in5,
        VN2CN0_bit => VN_data_out(3756),
        VN2CN1_bit => VN_data_out(3757),
        VN2CN2_bit => VN_data_out(3758),
        VN2CN3_bit => VN_data_out(3759),
        VN2CN4_bit => VN_data_out(3760),
        VN2CN5_bit => VN_data_out(3761),
        VN2CN0_sign => VN_sign_out(3756),
        VN2CN1_sign => VN_sign_out(3757),
        VN2CN2_sign => VN_sign_out(3758),
        VN2CN3_sign => VN_sign_out(3759),
        VN2CN4_sign => VN_sign_out(3760),
        VN2CN5_sign => VN_sign_out(3761),
        codeword => codeword(626),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN627 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3767 downto 3762),
        Din0 => VN627_in0,
        Din1 => VN627_in1,
        Din2 => VN627_in2,
        Din3 => VN627_in3,
        Din4 => VN627_in4,
        Din5 => VN627_in5,
        VN2CN0_bit => VN_data_out(3762),
        VN2CN1_bit => VN_data_out(3763),
        VN2CN2_bit => VN_data_out(3764),
        VN2CN3_bit => VN_data_out(3765),
        VN2CN4_bit => VN_data_out(3766),
        VN2CN5_bit => VN_data_out(3767),
        VN2CN0_sign => VN_sign_out(3762),
        VN2CN1_sign => VN_sign_out(3763),
        VN2CN2_sign => VN_sign_out(3764),
        VN2CN3_sign => VN_sign_out(3765),
        VN2CN4_sign => VN_sign_out(3766),
        VN2CN5_sign => VN_sign_out(3767),
        codeword => codeword(627),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN628 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3773 downto 3768),
        Din0 => VN628_in0,
        Din1 => VN628_in1,
        Din2 => VN628_in2,
        Din3 => VN628_in3,
        Din4 => VN628_in4,
        Din5 => VN628_in5,
        VN2CN0_bit => VN_data_out(3768),
        VN2CN1_bit => VN_data_out(3769),
        VN2CN2_bit => VN_data_out(3770),
        VN2CN3_bit => VN_data_out(3771),
        VN2CN4_bit => VN_data_out(3772),
        VN2CN5_bit => VN_data_out(3773),
        VN2CN0_sign => VN_sign_out(3768),
        VN2CN1_sign => VN_sign_out(3769),
        VN2CN2_sign => VN_sign_out(3770),
        VN2CN3_sign => VN_sign_out(3771),
        VN2CN4_sign => VN_sign_out(3772),
        VN2CN5_sign => VN_sign_out(3773),
        codeword => codeword(628),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN629 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3779 downto 3774),
        Din0 => VN629_in0,
        Din1 => VN629_in1,
        Din2 => VN629_in2,
        Din3 => VN629_in3,
        Din4 => VN629_in4,
        Din5 => VN629_in5,
        VN2CN0_bit => VN_data_out(3774),
        VN2CN1_bit => VN_data_out(3775),
        VN2CN2_bit => VN_data_out(3776),
        VN2CN3_bit => VN_data_out(3777),
        VN2CN4_bit => VN_data_out(3778),
        VN2CN5_bit => VN_data_out(3779),
        VN2CN0_sign => VN_sign_out(3774),
        VN2CN1_sign => VN_sign_out(3775),
        VN2CN2_sign => VN_sign_out(3776),
        VN2CN3_sign => VN_sign_out(3777),
        VN2CN4_sign => VN_sign_out(3778),
        VN2CN5_sign => VN_sign_out(3779),
        codeword => codeword(629),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN630 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3785 downto 3780),
        Din0 => VN630_in0,
        Din1 => VN630_in1,
        Din2 => VN630_in2,
        Din3 => VN630_in3,
        Din4 => VN630_in4,
        Din5 => VN630_in5,
        VN2CN0_bit => VN_data_out(3780),
        VN2CN1_bit => VN_data_out(3781),
        VN2CN2_bit => VN_data_out(3782),
        VN2CN3_bit => VN_data_out(3783),
        VN2CN4_bit => VN_data_out(3784),
        VN2CN5_bit => VN_data_out(3785),
        VN2CN0_sign => VN_sign_out(3780),
        VN2CN1_sign => VN_sign_out(3781),
        VN2CN2_sign => VN_sign_out(3782),
        VN2CN3_sign => VN_sign_out(3783),
        VN2CN4_sign => VN_sign_out(3784),
        VN2CN5_sign => VN_sign_out(3785),
        codeword => codeword(630),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN631 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3791 downto 3786),
        Din0 => VN631_in0,
        Din1 => VN631_in1,
        Din2 => VN631_in2,
        Din3 => VN631_in3,
        Din4 => VN631_in4,
        Din5 => VN631_in5,
        VN2CN0_bit => VN_data_out(3786),
        VN2CN1_bit => VN_data_out(3787),
        VN2CN2_bit => VN_data_out(3788),
        VN2CN3_bit => VN_data_out(3789),
        VN2CN4_bit => VN_data_out(3790),
        VN2CN5_bit => VN_data_out(3791),
        VN2CN0_sign => VN_sign_out(3786),
        VN2CN1_sign => VN_sign_out(3787),
        VN2CN2_sign => VN_sign_out(3788),
        VN2CN3_sign => VN_sign_out(3789),
        VN2CN4_sign => VN_sign_out(3790),
        VN2CN5_sign => VN_sign_out(3791),
        codeword => codeword(631),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN632 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3797 downto 3792),
        Din0 => VN632_in0,
        Din1 => VN632_in1,
        Din2 => VN632_in2,
        Din3 => VN632_in3,
        Din4 => VN632_in4,
        Din5 => VN632_in5,
        VN2CN0_bit => VN_data_out(3792),
        VN2CN1_bit => VN_data_out(3793),
        VN2CN2_bit => VN_data_out(3794),
        VN2CN3_bit => VN_data_out(3795),
        VN2CN4_bit => VN_data_out(3796),
        VN2CN5_bit => VN_data_out(3797),
        VN2CN0_sign => VN_sign_out(3792),
        VN2CN1_sign => VN_sign_out(3793),
        VN2CN2_sign => VN_sign_out(3794),
        VN2CN3_sign => VN_sign_out(3795),
        VN2CN4_sign => VN_sign_out(3796),
        VN2CN5_sign => VN_sign_out(3797),
        codeword => codeword(632),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN633 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3803 downto 3798),
        Din0 => VN633_in0,
        Din1 => VN633_in1,
        Din2 => VN633_in2,
        Din3 => VN633_in3,
        Din4 => VN633_in4,
        Din5 => VN633_in5,
        VN2CN0_bit => VN_data_out(3798),
        VN2CN1_bit => VN_data_out(3799),
        VN2CN2_bit => VN_data_out(3800),
        VN2CN3_bit => VN_data_out(3801),
        VN2CN4_bit => VN_data_out(3802),
        VN2CN5_bit => VN_data_out(3803),
        VN2CN0_sign => VN_sign_out(3798),
        VN2CN1_sign => VN_sign_out(3799),
        VN2CN2_sign => VN_sign_out(3800),
        VN2CN3_sign => VN_sign_out(3801),
        VN2CN4_sign => VN_sign_out(3802),
        VN2CN5_sign => VN_sign_out(3803),
        codeword => codeword(633),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN634 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3809 downto 3804),
        Din0 => VN634_in0,
        Din1 => VN634_in1,
        Din2 => VN634_in2,
        Din3 => VN634_in3,
        Din4 => VN634_in4,
        Din5 => VN634_in5,
        VN2CN0_bit => VN_data_out(3804),
        VN2CN1_bit => VN_data_out(3805),
        VN2CN2_bit => VN_data_out(3806),
        VN2CN3_bit => VN_data_out(3807),
        VN2CN4_bit => VN_data_out(3808),
        VN2CN5_bit => VN_data_out(3809),
        VN2CN0_sign => VN_sign_out(3804),
        VN2CN1_sign => VN_sign_out(3805),
        VN2CN2_sign => VN_sign_out(3806),
        VN2CN3_sign => VN_sign_out(3807),
        VN2CN4_sign => VN_sign_out(3808),
        VN2CN5_sign => VN_sign_out(3809),
        codeword => codeword(634),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN635 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3815 downto 3810),
        Din0 => VN635_in0,
        Din1 => VN635_in1,
        Din2 => VN635_in2,
        Din3 => VN635_in3,
        Din4 => VN635_in4,
        Din5 => VN635_in5,
        VN2CN0_bit => VN_data_out(3810),
        VN2CN1_bit => VN_data_out(3811),
        VN2CN2_bit => VN_data_out(3812),
        VN2CN3_bit => VN_data_out(3813),
        VN2CN4_bit => VN_data_out(3814),
        VN2CN5_bit => VN_data_out(3815),
        VN2CN0_sign => VN_sign_out(3810),
        VN2CN1_sign => VN_sign_out(3811),
        VN2CN2_sign => VN_sign_out(3812),
        VN2CN3_sign => VN_sign_out(3813),
        VN2CN4_sign => VN_sign_out(3814),
        VN2CN5_sign => VN_sign_out(3815),
        codeword => codeword(635),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN636 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3821 downto 3816),
        Din0 => VN636_in0,
        Din1 => VN636_in1,
        Din2 => VN636_in2,
        Din3 => VN636_in3,
        Din4 => VN636_in4,
        Din5 => VN636_in5,
        VN2CN0_bit => VN_data_out(3816),
        VN2CN1_bit => VN_data_out(3817),
        VN2CN2_bit => VN_data_out(3818),
        VN2CN3_bit => VN_data_out(3819),
        VN2CN4_bit => VN_data_out(3820),
        VN2CN5_bit => VN_data_out(3821),
        VN2CN0_sign => VN_sign_out(3816),
        VN2CN1_sign => VN_sign_out(3817),
        VN2CN2_sign => VN_sign_out(3818),
        VN2CN3_sign => VN_sign_out(3819),
        VN2CN4_sign => VN_sign_out(3820),
        VN2CN5_sign => VN_sign_out(3821),
        codeword => codeword(636),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN637 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3827 downto 3822),
        Din0 => VN637_in0,
        Din1 => VN637_in1,
        Din2 => VN637_in2,
        Din3 => VN637_in3,
        Din4 => VN637_in4,
        Din5 => VN637_in5,
        VN2CN0_bit => VN_data_out(3822),
        VN2CN1_bit => VN_data_out(3823),
        VN2CN2_bit => VN_data_out(3824),
        VN2CN3_bit => VN_data_out(3825),
        VN2CN4_bit => VN_data_out(3826),
        VN2CN5_bit => VN_data_out(3827),
        VN2CN0_sign => VN_sign_out(3822),
        VN2CN1_sign => VN_sign_out(3823),
        VN2CN2_sign => VN_sign_out(3824),
        VN2CN3_sign => VN_sign_out(3825),
        VN2CN4_sign => VN_sign_out(3826),
        VN2CN5_sign => VN_sign_out(3827),
        codeword => codeword(637),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN638 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3833 downto 3828),
        Din0 => VN638_in0,
        Din1 => VN638_in1,
        Din2 => VN638_in2,
        Din3 => VN638_in3,
        Din4 => VN638_in4,
        Din5 => VN638_in5,
        VN2CN0_bit => VN_data_out(3828),
        VN2CN1_bit => VN_data_out(3829),
        VN2CN2_bit => VN_data_out(3830),
        VN2CN3_bit => VN_data_out(3831),
        VN2CN4_bit => VN_data_out(3832),
        VN2CN5_bit => VN_data_out(3833),
        VN2CN0_sign => VN_sign_out(3828),
        VN2CN1_sign => VN_sign_out(3829),
        VN2CN2_sign => VN_sign_out(3830),
        VN2CN3_sign => VN_sign_out(3831),
        VN2CN4_sign => VN_sign_out(3832),
        VN2CN5_sign => VN_sign_out(3833),
        codeword => codeword(638),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN639 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3839 downto 3834),
        Din0 => VN639_in0,
        Din1 => VN639_in1,
        Din2 => VN639_in2,
        Din3 => VN639_in3,
        Din4 => VN639_in4,
        Din5 => VN639_in5,
        VN2CN0_bit => VN_data_out(3834),
        VN2CN1_bit => VN_data_out(3835),
        VN2CN2_bit => VN_data_out(3836),
        VN2CN3_bit => VN_data_out(3837),
        VN2CN4_bit => VN_data_out(3838),
        VN2CN5_bit => VN_data_out(3839),
        VN2CN0_sign => VN_sign_out(3834),
        VN2CN1_sign => VN_sign_out(3835),
        VN2CN2_sign => VN_sign_out(3836),
        VN2CN3_sign => VN_sign_out(3837),
        VN2CN4_sign => VN_sign_out(3838),
        VN2CN5_sign => VN_sign_out(3839),
        codeword => codeword(639),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN640 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3845 downto 3840),
        Din0 => VN640_in0,
        Din1 => VN640_in1,
        Din2 => VN640_in2,
        Din3 => VN640_in3,
        Din4 => VN640_in4,
        Din5 => VN640_in5,
        VN2CN0_bit => VN_data_out(3840),
        VN2CN1_bit => VN_data_out(3841),
        VN2CN2_bit => VN_data_out(3842),
        VN2CN3_bit => VN_data_out(3843),
        VN2CN4_bit => VN_data_out(3844),
        VN2CN5_bit => VN_data_out(3845),
        VN2CN0_sign => VN_sign_out(3840),
        VN2CN1_sign => VN_sign_out(3841),
        VN2CN2_sign => VN_sign_out(3842),
        VN2CN3_sign => VN_sign_out(3843),
        VN2CN4_sign => VN_sign_out(3844),
        VN2CN5_sign => VN_sign_out(3845),
        codeword => codeword(640),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN641 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3851 downto 3846),
        Din0 => VN641_in0,
        Din1 => VN641_in1,
        Din2 => VN641_in2,
        Din3 => VN641_in3,
        Din4 => VN641_in4,
        Din5 => VN641_in5,
        VN2CN0_bit => VN_data_out(3846),
        VN2CN1_bit => VN_data_out(3847),
        VN2CN2_bit => VN_data_out(3848),
        VN2CN3_bit => VN_data_out(3849),
        VN2CN4_bit => VN_data_out(3850),
        VN2CN5_bit => VN_data_out(3851),
        VN2CN0_sign => VN_sign_out(3846),
        VN2CN1_sign => VN_sign_out(3847),
        VN2CN2_sign => VN_sign_out(3848),
        VN2CN3_sign => VN_sign_out(3849),
        VN2CN4_sign => VN_sign_out(3850),
        VN2CN5_sign => VN_sign_out(3851),
        codeword => codeword(641),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN642 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3857 downto 3852),
        Din0 => VN642_in0,
        Din1 => VN642_in1,
        Din2 => VN642_in2,
        Din3 => VN642_in3,
        Din4 => VN642_in4,
        Din5 => VN642_in5,
        VN2CN0_bit => VN_data_out(3852),
        VN2CN1_bit => VN_data_out(3853),
        VN2CN2_bit => VN_data_out(3854),
        VN2CN3_bit => VN_data_out(3855),
        VN2CN4_bit => VN_data_out(3856),
        VN2CN5_bit => VN_data_out(3857),
        VN2CN0_sign => VN_sign_out(3852),
        VN2CN1_sign => VN_sign_out(3853),
        VN2CN2_sign => VN_sign_out(3854),
        VN2CN3_sign => VN_sign_out(3855),
        VN2CN4_sign => VN_sign_out(3856),
        VN2CN5_sign => VN_sign_out(3857),
        codeword => codeword(642),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN643 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3863 downto 3858),
        Din0 => VN643_in0,
        Din1 => VN643_in1,
        Din2 => VN643_in2,
        Din3 => VN643_in3,
        Din4 => VN643_in4,
        Din5 => VN643_in5,
        VN2CN0_bit => VN_data_out(3858),
        VN2CN1_bit => VN_data_out(3859),
        VN2CN2_bit => VN_data_out(3860),
        VN2CN3_bit => VN_data_out(3861),
        VN2CN4_bit => VN_data_out(3862),
        VN2CN5_bit => VN_data_out(3863),
        VN2CN0_sign => VN_sign_out(3858),
        VN2CN1_sign => VN_sign_out(3859),
        VN2CN2_sign => VN_sign_out(3860),
        VN2CN3_sign => VN_sign_out(3861),
        VN2CN4_sign => VN_sign_out(3862),
        VN2CN5_sign => VN_sign_out(3863),
        codeword => codeword(643),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN644 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3869 downto 3864),
        Din0 => VN644_in0,
        Din1 => VN644_in1,
        Din2 => VN644_in2,
        Din3 => VN644_in3,
        Din4 => VN644_in4,
        Din5 => VN644_in5,
        VN2CN0_bit => VN_data_out(3864),
        VN2CN1_bit => VN_data_out(3865),
        VN2CN2_bit => VN_data_out(3866),
        VN2CN3_bit => VN_data_out(3867),
        VN2CN4_bit => VN_data_out(3868),
        VN2CN5_bit => VN_data_out(3869),
        VN2CN0_sign => VN_sign_out(3864),
        VN2CN1_sign => VN_sign_out(3865),
        VN2CN2_sign => VN_sign_out(3866),
        VN2CN3_sign => VN_sign_out(3867),
        VN2CN4_sign => VN_sign_out(3868),
        VN2CN5_sign => VN_sign_out(3869),
        codeword => codeword(644),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN645 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3875 downto 3870),
        Din0 => VN645_in0,
        Din1 => VN645_in1,
        Din2 => VN645_in2,
        Din3 => VN645_in3,
        Din4 => VN645_in4,
        Din5 => VN645_in5,
        VN2CN0_bit => VN_data_out(3870),
        VN2CN1_bit => VN_data_out(3871),
        VN2CN2_bit => VN_data_out(3872),
        VN2CN3_bit => VN_data_out(3873),
        VN2CN4_bit => VN_data_out(3874),
        VN2CN5_bit => VN_data_out(3875),
        VN2CN0_sign => VN_sign_out(3870),
        VN2CN1_sign => VN_sign_out(3871),
        VN2CN2_sign => VN_sign_out(3872),
        VN2CN3_sign => VN_sign_out(3873),
        VN2CN4_sign => VN_sign_out(3874),
        VN2CN5_sign => VN_sign_out(3875),
        codeword => codeword(645),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN646 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3881 downto 3876),
        Din0 => VN646_in0,
        Din1 => VN646_in1,
        Din2 => VN646_in2,
        Din3 => VN646_in3,
        Din4 => VN646_in4,
        Din5 => VN646_in5,
        VN2CN0_bit => VN_data_out(3876),
        VN2CN1_bit => VN_data_out(3877),
        VN2CN2_bit => VN_data_out(3878),
        VN2CN3_bit => VN_data_out(3879),
        VN2CN4_bit => VN_data_out(3880),
        VN2CN5_bit => VN_data_out(3881),
        VN2CN0_sign => VN_sign_out(3876),
        VN2CN1_sign => VN_sign_out(3877),
        VN2CN2_sign => VN_sign_out(3878),
        VN2CN3_sign => VN_sign_out(3879),
        VN2CN4_sign => VN_sign_out(3880),
        VN2CN5_sign => VN_sign_out(3881),
        codeword => codeword(646),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN647 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3887 downto 3882),
        Din0 => VN647_in0,
        Din1 => VN647_in1,
        Din2 => VN647_in2,
        Din3 => VN647_in3,
        Din4 => VN647_in4,
        Din5 => VN647_in5,
        VN2CN0_bit => VN_data_out(3882),
        VN2CN1_bit => VN_data_out(3883),
        VN2CN2_bit => VN_data_out(3884),
        VN2CN3_bit => VN_data_out(3885),
        VN2CN4_bit => VN_data_out(3886),
        VN2CN5_bit => VN_data_out(3887),
        VN2CN0_sign => VN_sign_out(3882),
        VN2CN1_sign => VN_sign_out(3883),
        VN2CN2_sign => VN_sign_out(3884),
        VN2CN3_sign => VN_sign_out(3885),
        VN2CN4_sign => VN_sign_out(3886),
        VN2CN5_sign => VN_sign_out(3887),
        codeword => codeword(647),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN648 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3893 downto 3888),
        Din0 => VN648_in0,
        Din1 => VN648_in1,
        Din2 => VN648_in2,
        Din3 => VN648_in3,
        Din4 => VN648_in4,
        Din5 => VN648_in5,
        VN2CN0_bit => VN_data_out(3888),
        VN2CN1_bit => VN_data_out(3889),
        VN2CN2_bit => VN_data_out(3890),
        VN2CN3_bit => VN_data_out(3891),
        VN2CN4_bit => VN_data_out(3892),
        VN2CN5_bit => VN_data_out(3893),
        VN2CN0_sign => VN_sign_out(3888),
        VN2CN1_sign => VN_sign_out(3889),
        VN2CN2_sign => VN_sign_out(3890),
        VN2CN3_sign => VN_sign_out(3891),
        VN2CN4_sign => VN_sign_out(3892),
        VN2CN5_sign => VN_sign_out(3893),
        codeword => codeword(648),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN649 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3899 downto 3894),
        Din0 => VN649_in0,
        Din1 => VN649_in1,
        Din2 => VN649_in2,
        Din3 => VN649_in3,
        Din4 => VN649_in4,
        Din5 => VN649_in5,
        VN2CN0_bit => VN_data_out(3894),
        VN2CN1_bit => VN_data_out(3895),
        VN2CN2_bit => VN_data_out(3896),
        VN2CN3_bit => VN_data_out(3897),
        VN2CN4_bit => VN_data_out(3898),
        VN2CN5_bit => VN_data_out(3899),
        VN2CN0_sign => VN_sign_out(3894),
        VN2CN1_sign => VN_sign_out(3895),
        VN2CN2_sign => VN_sign_out(3896),
        VN2CN3_sign => VN_sign_out(3897),
        VN2CN4_sign => VN_sign_out(3898),
        VN2CN5_sign => VN_sign_out(3899),
        codeword => codeword(649),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN650 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3905 downto 3900),
        Din0 => VN650_in0,
        Din1 => VN650_in1,
        Din2 => VN650_in2,
        Din3 => VN650_in3,
        Din4 => VN650_in4,
        Din5 => VN650_in5,
        VN2CN0_bit => VN_data_out(3900),
        VN2CN1_bit => VN_data_out(3901),
        VN2CN2_bit => VN_data_out(3902),
        VN2CN3_bit => VN_data_out(3903),
        VN2CN4_bit => VN_data_out(3904),
        VN2CN5_bit => VN_data_out(3905),
        VN2CN0_sign => VN_sign_out(3900),
        VN2CN1_sign => VN_sign_out(3901),
        VN2CN2_sign => VN_sign_out(3902),
        VN2CN3_sign => VN_sign_out(3903),
        VN2CN4_sign => VN_sign_out(3904),
        VN2CN5_sign => VN_sign_out(3905),
        codeword => codeword(650),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN651 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3911 downto 3906),
        Din0 => VN651_in0,
        Din1 => VN651_in1,
        Din2 => VN651_in2,
        Din3 => VN651_in3,
        Din4 => VN651_in4,
        Din5 => VN651_in5,
        VN2CN0_bit => VN_data_out(3906),
        VN2CN1_bit => VN_data_out(3907),
        VN2CN2_bit => VN_data_out(3908),
        VN2CN3_bit => VN_data_out(3909),
        VN2CN4_bit => VN_data_out(3910),
        VN2CN5_bit => VN_data_out(3911),
        VN2CN0_sign => VN_sign_out(3906),
        VN2CN1_sign => VN_sign_out(3907),
        VN2CN2_sign => VN_sign_out(3908),
        VN2CN3_sign => VN_sign_out(3909),
        VN2CN4_sign => VN_sign_out(3910),
        VN2CN5_sign => VN_sign_out(3911),
        codeword => codeword(651),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN652 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3917 downto 3912),
        Din0 => VN652_in0,
        Din1 => VN652_in1,
        Din2 => VN652_in2,
        Din3 => VN652_in3,
        Din4 => VN652_in4,
        Din5 => VN652_in5,
        VN2CN0_bit => VN_data_out(3912),
        VN2CN1_bit => VN_data_out(3913),
        VN2CN2_bit => VN_data_out(3914),
        VN2CN3_bit => VN_data_out(3915),
        VN2CN4_bit => VN_data_out(3916),
        VN2CN5_bit => VN_data_out(3917),
        VN2CN0_sign => VN_sign_out(3912),
        VN2CN1_sign => VN_sign_out(3913),
        VN2CN2_sign => VN_sign_out(3914),
        VN2CN3_sign => VN_sign_out(3915),
        VN2CN4_sign => VN_sign_out(3916),
        VN2CN5_sign => VN_sign_out(3917),
        codeword => codeword(652),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN653 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3923 downto 3918),
        Din0 => VN653_in0,
        Din1 => VN653_in1,
        Din2 => VN653_in2,
        Din3 => VN653_in3,
        Din4 => VN653_in4,
        Din5 => VN653_in5,
        VN2CN0_bit => VN_data_out(3918),
        VN2CN1_bit => VN_data_out(3919),
        VN2CN2_bit => VN_data_out(3920),
        VN2CN3_bit => VN_data_out(3921),
        VN2CN4_bit => VN_data_out(3922),
        VN2CN5_bit => VN_data_out(3923),
        VN2CN0_sign => VN_sign_out(3918),
        VN2CN1_sign => VN_sign_out(3919),
        VN2CN2_sign => VN_sign_out(3920),
        VN2CN3_sign => VN_sign_out(3921),
        VN2CN4_sign => VN_sign_out(3922),
        VN2CN5_sign => VN_sign_out(3923),
        codeword => codeword(653),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN654 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3929 downto 3924),
        Din0 => VN654_in0,
        Din1 => VN654_in1,
        Din2 => VN654_in2,
        Din3 => VN654_in3,
        Din4 => VN654_in4,
        Din5 => VN654_in5,
        VN2CN0_bit => VN_data_out(3924),
        VN2CN1_bit => VN_data_out(3925),
        VN2CN2_bit => VN_data_out(3926),
        VN2CN3_bit => VN_data_out(3927),
        VN2CN4_bit => VN_data_out(3928),
        VN2CN5_bit => VN_data_out(3929),
        VN2CN0_sign => VN_sign_out(3924),
        VN2CN1_sign => VN_sign_out(3925),
        VN2CN2_sign => VN_sign_out(3926),
        VN2CN3_sign => VN_sign_out(3927),
        VN2CN4_sign => VN_sign_out(3928),
        VN2CN5_sign => VN_sign_out(3929),
        codeword => codeword(654),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN655 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3935 downto 3930),
        Din0 => VN655_in0,
        Din1 => VN655_in1,
        Din2 => VN655_in2,
        Din3 => VN655_in3,
        Din4 => VN655_in4,
        Din5 => VN655_in5,
        VN2CN0_bit => VN_data_out(3930),
        VN2CN1_bit => VN_data_out(3931),
        VN2CN2_bit => VN_data_out(3932),
        VN2CN3_bit => VN_data_out(3933),
        VN2CN4_bit => VN_data_out(3934),
        VN2CN5_bit => VN_data_out(3935),
        VN2CN0_sign => VN_sign_out(3930),
        VN2CN1_sign => VN_sign_out(3931),
        VN2CN2_sign => VN_sign_out(3932),
        VN2CN3_sign => VN_sign_out(3933),
        VN2CN4_sign => VN_sign_out(3934),
        VN2CN5_sign => VN_sign_out(3935),
        codeword => codeword(655),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN656 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3941 downto 3936),
        Din0 => VN656_in0,
        Din1 => VN656_in1,
        Din2 => VN656_in2,
        Din3 => VN656_in3,
        Din4 => VN656_in4,
        Din5 => VN656_in5,
        VN2CN0_bit => VN_data_out(3936),
        VN2CN1_bit => VN_data_out(3937),
        VN2CN2_bit => VN_data_out(3938),
        VN2CN3_bit => VN_data_out(3939),
        VN2CN4_bit => VN_data_out(3940),
        VN2CN5_bit => VN_data_out(3941),
        VN2CN0_sign => VN_sign_out(3936),
        VN2CN1_sign => VN_sign_out(3937),
        VN2CN2_sign => VN_sign_out(3938),
        VN2CN3_sign => VN_sign_out(3939),
        VN2CN4_sign => VN_sign_out(3940),
        VN2CN5_sign => VN_sign_out(3941),
        codeword => codeword(656),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN657 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3947 downto 3942),
        Din0 => VN657_in0,
        Din1 => VN657_in1,
        Din2 => VN657_in2,
        Din3 => VN657_in3,
        Din4 => VN657_in4,
        Din5 => VN657_in5,
        VN2CN0_bit => VN_data_out(3942),
        VN2CN1_bit => VN_data_out(3943),
        VN2CN2_bit => VN_data_out(3944),
        VN2CN3_bit => VN_data_out(3945),
        VN2CN4_bit => VN_data_out(3946),
        VN2CN5_bit => VN_data_out(3947),
        VN2CN0_sign => VN_sign_out(3942),
        VN2CN1_sign => VN_sign_out(3943),
        VN2CN2_sign => VN_sign_out(3944),
        VN2CN3_sign => VN_sign_out(3945),
        VN2CN4_sign => VN_sign_out(3946),
        VN2CN5_sign => VN_sign_out(3947),
        codeword => codeword(657),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN658 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3953 downto 3948),
        Din0 => VN658_in0,
        Din1 => VN658_in1,
        Din2 => VN658_in2,
        Din3 => VN658_in3,
        Din4 => VN658_in4,
        Din5 => VN658_in5,
        VN2CN0_bit => VN_data_out(3948),
        VN2CN1_bit => VN_data_out(3949),
        VN2CN2_bit => VN_data_out(3950),
        VN2CN3_bit => VN_data_out(3951),
        VN2CN4_bit => VN_data_out(3952),
        VN2CN5_bit => VN_data_out(3953),
        VN2CN0_sign => VN_sign_out(3948),
        VN2CN1_sign => VN_sign_out(3949),
        VN2CN2_sign => VN_sign_out(3950),
        VN2CN3_sign => VN_sign_out(3951),
        VN2CN4_sign => VN_sign_out(3952),
        VN2CN5_sign => VN_sign_out(3953),
        codeword => codeword(658),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN659 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3959 downto 3954),
        Din0 => VN659_in0,
        Din1 => VN659_in1,
        Din2 => VN659_in2,
        Din3 => VN659_in3,
        Din4 => VN659_in4,
        Din5 => VN659_in5,
        VN2CN0_bit => VN_data_out(3954),
        VN2CN1_bit => VN_data_out(3955),
        VN2CN2_bit => VN_data_out(3956),
        VN2CN3_bit => VN_data_out(3957),
        VN2CN4_bit => VN_data_out(3958),
        VN2CN5_bit => VN_data_out(3959),
        VN2CN0_sign => VN_sign_out(3954),
        VN2CN1_sign => VN_sign_out(3955),
        VN2CN2_sign => VN_sign_out(3956),
        VN2CN3_sign => VN_sign_out(3957),
        VN2CN4_sign => VN_sign_out(3958),
        VN2CN5_sign => VN_sign_out(3959),
        codeword => codeword(659),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN660 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3965 downto 3960),
        Din0 => VN660_in0,
        Din1 => VN660_in1,
        Din2 => VN660_in2,
        Din3 => VN660_in3,
        Din4 => VN660_in4,
        Din5 => VN660_in5,
        VN2CN0_bit => VN_data_out(3960),
        VN2CN1_bit => VN_data_out(3961),
        VN2CN2_bit => VN_data_out(3962),
        VN2CN3_bit => VN_data_out(3963),
        VN2CN4_bit => VN_data_out(3964),
        VN2CN5_bit => VN_data_out(3965),
        VN2CN0_sign => VN_sign_out(3960),
        VN2CN1_sign => VN_sign_out(3961),
        VN2CN2_sign => VN_sign_out(3962),
        VN2CN3_sign => VN_sign_out(3963),
        VN2CN4_sign => VN_sign_out(3964),
        VN2CN5_sign => VN_sign_out(3965),
        codeword => codeword(660),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN661 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3971 downto 3966),
        Din0 => VN661_in0,
        Din1 => VN661_in1,
        Din2 => VN661_in2,
        Din3 => VN661_in3,
        Din4 => VN661_in4,
        Din5 => VN661_in5,
        VN2CN0_bit => VN_data_out(3966),
        VN2CN1_bit => VN_data_out(3967),
        VN2CN2_bit => VN_data_out(3968),
        VN2CN3_bit => VN_data_out(3969),
        VN2CN4_bit => VN_data_out(3970),
        VN2CN5_bit => VN_data_out(3971),
        VN2CN0_sign => VN_sign_out(3966),
        VN2CN1_sign => VN_sign_out(3967),
        VN2CN2_sign => VN_sign_out(3968),
        VN2CN3_sign => VN_sign_out(3969),
        VN2CN4_sign => VN_sign_out(3970),
        VN2CN5_sign => VN_sign_out(3971),
        codeword => codeword(661),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN662 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3977 downto 3972),
        Din0 => VN662_in0,
        Din1 => VN662_in1,
        Din2 => VN662_in2,
        Din3 => VN662_in3,
        Din4 => VN662_in4,
        Din5 => VN662_in5,
        VN2CN0_bit => VN_data_out(3972),
        VN2CN1_bit => VN_data_out(3973),
        VN2CN2_bit => VN_data_out(3974),
        VN2CN3_bit => VN_data_out(3975),
        VN2CN4_bit => VN_data_out(3976),
        VN2CN5_bit => VN_data_out(3977),
        VN2CN0_sign => VN_sign_out(3972),
        VN2CN1_sign => VN_sign_out(3973),
        VN2CN2_sign => VN_sign_out(3974),
        VN2CN3_sign => VN_sign_out(3975),
        VN2CN4_sign => VN_sign_out(3976),
        VN2CN5_sign => VN_sign_out(3977),
        codeword => codeword(662),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN663 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3983 downto 3978),
        Din0 => VN663_in0,
        Din1 => VN663_in1,
        Din2 => VN663_in2,
        Din3 => VN663_in3,
        Din4 => VN663_in4,
        Din5 => VN663_in5,
        VN2CN0_bit => VN_data_out(3978),
        VN2CN1_bit => VN_data_out(3979),
        VN2CN2_bit => VN_data_out(3980),
        VN2CN3_bit => VN_data_out(3981),
        VN2CN4_bit => VN_data_out(3982),
        VN2CN5_bit => VN_data_out(3983),
        VN2CN0_sign => VN_sign_out(3978),
        VN2CN1_sign => VN_sign_out(3979),
        VN2CN2_sign => VN_sign_out(3980),
        VN2CN3_sign => VN_sign_out(3981),
        VN2CN4_sign => VN_sign_out(3982),
        VN2CN5_sign => VN_sign_out(3983),
        codeword => codeword(663),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN664 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3989 downto 3984),
        Din0 => VN664_in0,
        Din1 => VN664_in1,
        Din2 => VN664_in2,
        Din3 => VN664_in3,
        Din4 => VN664_in4,
        Din5 => VN664_in5,
        VN2CN0_bit => VN_data_out(3984),
        VN2CN1_bit => VN_data_out(3985),
        VN2CN2_bit => VN_data_out(3986),
        VN2CN3_bit => VN_data_out(3987),
        VN2CN4_bit => VN_data_out(3988),
        VN2CN5_bit => VN_data_out(3989),
        VN2CN0_sign => VN_sign_out(3984),
        VN2CN1_sign => VN_sign_out(3985),
        VN2CN2_sign => VN_sign_out(3986),
        VN2CN3_sign => VN_sign_out(3987),
        VN2CN4_sign => VN_sign_out(3988),
        VN2CN5_sign => VN_sign_out(3989),
        codeword => codeword(664),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN665 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(3995 downto 3990),
        Din0 => VN665_in0,
        Din1 => VN665_in1,
        Din2 => VN665_in2,
        Din3 => VN665_in3,
        Din4 => VN665_in4,
        Din5 => VN665_in5,
        VN2CN0_bit => VN_data_out(3990),
        VN2CN1_bit => VN_data_out(3991),
        VN2CN2_bit => VN_data_out(3992),
        VN2CN3_bit => VN_data_out(3993),
        VN2CN4_bit => VN_data_out(3994),
        VN2CN5_bit => VN_data_out(3995),
        VN2CN0_sign => VN_sign_out(3990),
        VN2CN1_sign => VN_sign_out(3991),
        VN2CN2_sign => VN_sign_out(3992),
        VN2CN3_sign => VN_sign_out(3993),
        VN2CN4_sign => VN_sign_out(3994),
        VN2CN5_sign => VN_sign_out(3995),
        codeword => codeword(665),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN666 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4001 downto 3996),
        Din0 => VN666_in0,
        Din1 => VN666_in1,
        Din2 => VN666_in2,
        Din3 => VN666_in3,
        Din4 => VN666_in4,
        Din5 => VN666_in5,
        VN2CN0_bit => VN_data_out(3996),
        VN2CN1_bit => VN_data_out(3997),
        VN2CN2_bit => VN_data_out(3998),
        VN2CN3_bit => VN_data_out(3999),
        VN2CN4_bit => VN_data_out(4000),
        VN2CN5_bit => VN_data_out(4001),
        VN2CN0_sign => VN_sign_out(3996),
        VN2CN1_sign => VN_sign_out(3997),
        VN2CN2_sign => VN_sign_out(3998),
        VN2CN3_sign => VN_sign_out(3999),
        VN2CN4_sign => VN_sign_out(4000),
        VN2CN5_sign => VN_sign_out(4001),
        codeword => codeword(666),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN667 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4007 downto 4002),
        Din0 => VN667_in0,
        Din1 => VN667_in1,
        Din2 => VN667_in2,
        Din3 => VN667_in3,
        Din4 => VN667_in4,
        Din5 => VN667_in5,
        VN2CN0_bit => VN_data_out(4002),
        VN2CN1_bit => VN_data_out(4003),
        VN2CN2_bit => VN_data_out(4004),
        VN2CN3_bit => VN_data_out(4005),
        VN2CN4_bit => VN_data_out(4006),
        VN2CN5_bit => VN_data_out(4007),
        VN2CN0_sign => VN_sign_out(4002),
        VN2CN1_sign => VN_sign_out(4003),
        VN2CN2_sign => VN_sign_out(4004),
        VN2CN3_sign => VN_sign_out(4005),
        VN2CN4_sign => VN_sign_out(4006),
        VN2CN5_sign => VN_sign_out(4007),
        codeword => codeword(667),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN668 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4013 downto 4008),
        Din0 => VN668_in0,
        Din1 => VN668_in1,
        Din2 => VN668_in2,
        Din3 => VN668_in3,
        Din4 => VN668_in4,
        Din5 => VN668_in5,
        VN2CN0_bit => VN_data_out(4008),
        VN2CN1_bit => VN_data_out(4009),
        VN2CN2_bit => VN_data_out(4010),
        VN2CN3_bit => VN_data_out(4011),
        VN2CN4_bit => VN_data_out(4012),
        VN2CN5_bit => VN_data_out(4013),
        VN2CN0_sign => VN_sign_out(4008),
        VN2CN1_sign => VN_sign_out(4009),
        VN2CN2_sign => VN_sign_out(4010),
        VN2CN3_sign => VN_sign_out(4011),
        VN2CN4_sign => VN_sign_out(4012),
        VN2CN5_sign => VN_sign_out(4013),
        codeword => codeword(668),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN669 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4019 downto 4014),
        Din0 => VN669_in0,
        Din1 => VN669_in1,
        Din2 => VN669_in2,
        Din3 => VN669_in3,
        Din4 => VN669_in4,
        Din5 => VN669_in5,
        VN2CN0_bit => VN_data_out(4014),
        VN2CN1_bit => VN_data_out(4015),
        VN2CN2_bit => VN_data_out(4016),
        VN2CN3_bit => VN_data_out(4017),
        VN2CN4_bit => VN_data_out(4018),
        VN2CN5_bit => VN_data_out(4019),
        VN2CN0_sign => VN_sign_out(4014),
        VN2CN1_sign => VN_sign_out(4015),
        VN2CN2_sign => VN_sign_out(4016),
        VN2CN3_sign => VN_sign_out(4017),
        VN2CN4_sign => VN_sign_out(4018),
        VN2CN5_sign => VN_sign_out(4019),
        codeword => codeword(669),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN670 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4025 downto 4020),
        Din0 => VN670_in0,
        Din1 => VN670_in1,
        Din2 => VN670_in2,
        Din3 => VN670_in3,
        Din4 => VN670_in4,
        Din5 => VN670_in5,
        VN2CN0_bit => VN_data_out(4020),
        VN2CN1_bit => VN_data_out(4021),
        VN2CN2_bit => VN_data_out(4022),
        VN2CN3_bit => VN_data_out(4023),
        VN2CN4_bit => VN_data_out(4024),
        VN2CN5_bit => VN_data_out(4025),
        VN2CN0_sign => VN_sign_out(4020),
        VN2CN1_sign => VN_sign_out(4021),
        VN2CN2_sign => VN_sign_out(4022),
        VN2CN3_sign => VN_sign_out(4023),
        VN2CN4_sign => VN_sign_out(4024),
        VN2CN5_sign => VN_sign_out(4025),
        codeword => codeword(670),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN671 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4031 downto 4026),
        Din0 => VN671_in0,
        Din1 => VN671_in1,
        Din2 => VN671_in2,
        Din3 => VN671_in3,
        Din4 => VN671_in4,
        Din5 => VN671_in5,
        VN2CN0_bit => VN_data_out(4026),
        VN2CN1_bit => VN_data_out(4027),
        VN2CN2_bit => VN_data_out(4028),
        VN2CN3_bit => VN_data_out(4029),
        VN2CN4_bit => VN_data_out(4030),
        VN2CN5_bit => VN_data_out(4031),
        VN2CN0_sign => VN_sign_out(4026),
        VN2CN1_sign => VN_sign_out(4027),
        VN2CN2_sign => VN_sign_out(4028),
        VN2CN3_sign => VN_sign_out(4029),
        VN2CN4_sign => VN_sign_out(4030),
        VN2CN5_sign => VN_sign_out(4031),
        codeword => codeword(671),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN672 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4037 downto 4032),
        Din0 => VN672_in0,
        Din1 => VN672_in1,
        Din2 => VN672_in2,
        Din3 => VN672_in3,
        Din4 => VN672_in4,
        Din5 => VN672_in5,
        VN2CN0_bit => VN_data_out(4032),
        VN2CN1_bit => VN_data_out(4033),
        VN2CN2_bit => VN_data_out(4034),
        VN2CN3_bit => VN_data_out(4035),
        VN2CN4_bit => VN_data_out(4036),
        VN2CN5_bit => VN_data_out(4037),
        VN2CN0_sign => VN_sign_out(4032),
        VN2CN1_sign => VN_sign_out(4033),
        VN2CN2_sign => VN_sign_out(4034),
        VN2CN3_sign => VN_sign_out(4035),
        VN2CN4_sign => VN_sign_out(4036),
        VN2CN5_sign => VN_sign_out(4037),
        codeword => codeword(672),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN673 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4043 downto 4038),
        Din0 => VN673_in0,
        Din1 => VN673_in1,
        Din2 => VN673_in2,
        Din3 => VN673_in3,
        Din4 => VN673_in4,
        Din5 => VN673_in5,
        VN2CN0_bit => VN_data_out(4038),
        VN2CN1_bit => VN_data_out(4039),
        VN2CN2_bit => VN_data_out(4040),
        VN2CN3_bit => VN_data_out(4041),
        VN2CN4_bit => VN_data_out(4042),
        VN2CN5_bit => VN_data_out(4043),
        VN2CN0_sign => VN_sign_out(4038),
        VN2CN1_sign => VN_sign_out(4039),
        VN2CN2_sign => VN_sign_out(4040),
        VN2CN3_sign => VN_sign_out(4041),
        VN2CN4_sign => VN_sign_out(4042),
        VN2CN5_sign => VN_sign_out(4043),
        codeword => codeword(673),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN674 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4049 downto 4044),
        Din0 => VN674_in0,
        Din1 => VN674_in1,
        Din2 => VN674_in2,
        Din3 => VN674_in3,
        Din4 => VN674_in4,
        Din5 => VN674_in5,
        VN2CN0_bit => VN_data_out(4044),
        VN2CN1_bit => VN_data_out(4045),
        VN2CN2_bit => VN_data_out(4046),
        VN2CN3_bit => VN_data_out(4047),
        VN2CN4_bit => VN_data_out(4048),
        VN2CN5_bit => VN_data_out(4049),
        VN2CN0_sign => VN_sign_out(4044),
        VN2CN1_sign => VN_sign_out(4045),
        VN2CN2_sign => VN_sign_out(4046),
        VN2CN3_sign => VN_sign_out(4047),
        VN2CN4_sign => VN_sign_out(4048),
        VN2CN5_sign => VN_sign_out(4049),
        codeword => codeword(674),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN675 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4055 downto 4050),
        Din0 => VN675_in0,
        Din1 => VN675_in1,
        Din2 => VN675_in2,
        Din3 => VN675_in3,
        Din4 => VN675_in4,
        Din5 => VN675_in5,
        VN2CN0_bit => VN_data_out(4050),
        VN2CN1_bit => VN_data_out(4051),
        VN2CN2_bit => VN_data_out(4052),
        VN2CN3_bit => VN_data_out(4053),
        VN2CN4_bit => VN_data_out(4054),
        VN2CN5_bit => VN_data_out(4055),
        VN2CN0_sign => VN_sign_out(4050),
        VN2CN1_sign => VN_sign_out(4051),
        VN2CN2_sign => VN_sign_out(4052),
        VN2CN3_sign => VN_sign_out(4053),
        VN2CN4_sign => VN_sign_out(4054),
        VN2CN5_sign => VN_sign_out(4055),
        codeword => codeword(675),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN676 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4061 downto 4056),
        Din0 => VN676_in0,
        Din1 => VN676_in1,
        Din2 => VN676_in2,
        Din3 => VN676_in3,
        Din4 => VN676_in4,
        Din5 => VN676_in5,
        VN2CN0_bit => VN_data_out(4056),
        VN2CN1_bit => VN_data_out(4057),
        VN2CN2_bit => VN_data_out(4058),
        VN2CN3_bit => VN_data_out(4059),
        VN2CN4_bit => VN_data_out(4060),
        VN2CN5_bit => VN_data_out(4061),
        VN2CN0_sign => VN_sign_out(4056),
        VN2CN1_sign => VN_sign_out(4057),
        VN2CN2_sign => VN_sign_out(4058),
        VN2CN3_sign => VN_sign_out(4059),
        VN2CN4_sign => VN_sign_out(4060),
        VN2CN5_sign => VN_sign_out(4061),
        codeword => codeword(676),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN677 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4067 downto 4062),
        Din0 => VN677_in0,
        Din1 => VN677_in1,
        Din2 => VN677_in2,
        Din3 => VN677_in3,
        Din4 => VN677_in4,
        Din5 => VN677_in5,
        VN2CN0_bit => VN_data_out(4062),
        VN2CN1_bit => VN_data_out(4063),
        VN2CN2_bit => VN_data_out(4064),
        VN2CN3_bit => VN_data_out(4065),
        VN2CN4_bit => VN_data_out(4066),
        VN2CN5_bit => VN_data_out(4067),
        VN2CN0_sign => VN_sign_out(4062),
        VN2CN1_sign => VN_sign_out(4063),
        VN2CN2_sign => VN_sign_out(4064),
        VN2CN3_sign => VN_sign_out(4065),
        VN2CN4_sign => VN_sign_out(4066),
        VN2CN5_sign => VN_sign_out(4067),
        codeword => codeword(677),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN678 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4073 downto 4068),
        Din0 => VN678_in0,
        Din1 => VN678_in1,
        Din2 => VN678_in2,
        Din3 => VN678_in3,
        Din4 => VN678_in4,
        Din5 => VN678_in5,
        VN2CN0_bit => VN_data_out(4068),
        VN2CN1_bit => VN_data_out(4069),
        VN2CN2_bit => VN_data_out(4070),
        VN2CN3_bit => VN_data_out(4071),
        VN2CN4_bit => VN_data_out(4072),
        VN2CN5_bit => VN_data_out(4073),
        VN2CN0_sign => VN_sign_out(4068),
        VN2CN1_sign => VN_sign_out(4069),
        VN2CN2_sign => VN_sign_out(4070),
        VN2CN3_sign => VN_sign_out(4071),
        VN2CN4_sign => VN_sign_out(4072),
        VN2CN5_sign => VN_sign_out(4073),
        codeword => codeword(678),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN679 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4079 downto 4074),
        Din0 => VN679_in0,
        Din1 => VN679_in1,
        Din2 => VN679_in2,
        Din3 => VN679_in3,
        Din4 => VN679_in4,
        Din5 => VN679_in5,
        VN2CN0_bit => VN_data_out(4074),
        VN2CN1_bit => VN_data_out(4075),
        VN2CN2_bit => VN_data_out(4076),
        VN2CN3_bit => VN_data_out(4077),
        VN2CN4_bit => VN_data_out(4078),
        VN2CN5_bit => VN_data_out(4079),
        VN2CN0_sign => VN_sign_out(4074),
        VN2CN1_sign => VN_sign_out(4075),
        VN2CN2_sign => VN_sign_out(4076),
        VN2CN3_sign => VN_sign_out(4077),
        VN2CN4_sign => VN_sign_out(4078),
        VN2CN5_sign => VN_sign_out(4079),
        codeword => codeword(679),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN680 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4085 downto 4080),
        Din0 => VN680_in0,
        Din1 => VN680_in1,
        Din2 => VN680_in2,
        Din3 => VN680_in3,
        Din4 => VN680_in4,
        Din5 => VN680_in5,
        VN2CN0_bit => VN_data_out(4080),
        VN2CN1_bit => VN_data_out(4081),
        VN2CN2_bit => VN_data_out(4082),
        VN2CN3_bit => VN_data_out(4083),
        VN2CN4_bit => VN_data_out(4084),
        VN2CN5_bit => VN_data_out(4085),
        VN2CN0_sign => VN_sign_out(4080),
        VN2CN1_sign => VN_sign_out(4081),
        VN2CN2_sign => VN_sign_out(4082),
        VN2CN3_sign => VN_sign_out(4083),
        VN2CN4_sign => VN_sign_out(4084),
        VN2CN5_sign => VN_sign_out(4085),
        codeword => codeword(680),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN681 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4091 downto 4086),
        Din0 => VN681_in0,
        Din1 => VN681_in1,
        Din2 => VN681_in2,
        Din3 => VN681_in3,
        Din4 => VN681_in4,
        Din5 => VN681_in5,
        VN2CN0_bit => VN_data_out(4086),
        VN2CN1_bit => VN_data_out(4087),
        VN2CN2_bit => VN_data_out(4088),
        VN2CN3_bit => VN_data_out(4089),
        VN2CN4_bit => VN_data_out(4090),
        VN2CN5_bit => VN_data_out(4091),
        VN2CN0_sign => VN_sign_out(4086),
        VN2CN1_sign => VN_sign_out(4087),
        VN2CN2_sign => VN_sign_out(4088),
        VN2CN3_sign => VN_sign_out(4089),
        VN2CN4_sign => VN_sign_out(4090),
        VN2CN5_sign => VN_sign_out(4091),
        codeword => codeword(681),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN682 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4097 downto 4092),
        Din0 => VN682_in0,
        Din1 => VN682_in1,
        Din2 => VN682_in2,
        Din3 => VN682_in3,
        Din4 => VN682_in4,
        Din5 => VN682_in5,
        VN2CN0_bit => VN_data_out(4092),
        VN2CN1_bit => VN_data_out(4093),
        VN2CN2_bit => VN_data_out(4094),
        VN2CN3_bit => VN_data_out(4095),
        VN2CN4_bit => VN_data_out(4096),
        VN2CN5_bit => VN_data_out(4097),
        VN2CN0_sign => VN_sign_out(4092),
        VN2CN1_sign => VN_sign_out(4093),
        VN2CN2_sign => VN_sign_out(4094),
        VN2CN3_sign => VN_sign_out(4095),
        VN2CN4_sign => VN_sign_out(4096),
        VN2CN5_sign => VN_sign_out(4097),
        codeword => codeword(682),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN683 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4103 downto 4098),
        Din0 => VN683_in0,
        Din1 => VN683_in1,
        Din2 => VN683_in2,
        Din3 => VN683_in3,
        Din4 => VN683_in4,
        Din5 => VN683_in5,
        VN2CN0_bit => VN_data_out(4098),
        VN2CN1_bit => VN_data_out(4099),
        VN2CN2_bit => VN_data_out(4100),
        VN2CN3_bit => VN_data_out(4101),
        VN2CN4_bit => VN_data_out(4102),
        VN2CN5_bit => VN_data_out(4103),
        VN2CN0_sign => VN_sign_out(4098),
        VN2CN1_sign => VN_sign_out(4099),
        VN2CN2_sign => VN_sign_out(4100),
        VN2CN3_sign => VN_sign_out(4101),
        VN2CN4_sign => VN_sign_out(4102),
        VN2CN5_sign => VN_sign_out(4103),
        codeword => codeword(683),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN684 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4109 downto 4104),
        Din0 => VN684_in0,
        Din1 => VN684_in1,
        Din2 => VN684_in2,
        Din3 => VN684_in3,
        Din4 => VN684_in4,
        Din5 => VN684_in5,
        VN2CN0_bit => VN_data_out(4104),
        VN2CN1_bit => VN_data_out(4105),
        VN2CN2_bit => VN_data_out(4106),
        VN2CN3_bit => VN_data_out(4107),
        VN2CN4_bit => VN_data_out(4108),
        VN2CN5_bit => VN_data_out(4109),
        VN2CN0_sign => VN_sign_out(4104),
        VN2CN1_sign => VN_sign_out(4105),
        VN2CN2_sign => VN_sign_out(4106),
        VN2CN3_sign => VN_sign_out(4107),
        VN2CN4_sign => VN_sign_out(4108),
        VN2CN5_sign => VN_sign_out(4109),
        codeword => codeword(684),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN685 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4115 downto 4110),
        Din0 => VN685_in0,
        Din1 => VN685_in1,
        Din2 => VN685_in2,
        Din3 => VN685_in3,
        Din4 => VN685_in4,
        Din5 => VN685_in5,
        VN2CN0_bit => VN_data_out(4110),
        VN2CN1_bit => VN_data_out(4111),
        VN2CN2_bit => VN_data_out(4112),
        VN2CN3_bit => VN_data_out(4113),
        VN2CN4_bit => VN_data_out(4114),
        VN2CN5_bit => VN_data_out(4115),
        VN2CN0_sign => VN_sign_out(4110),
        VN2CN1_sign => VN_sign_out(4111),
        VN2CN2_sign => VN_sign_out(4112),
        VN2CN3_sign => VN_sign_out(4113),
        VN2CN4_sign => VN_sign_out(4114),
        VN2CN5_sign => VN_sign_out(4115),
        codeword => codeword(685),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN686 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4121 downto 4116),
        Din0 => VN686_in0,
        Din1 => VN686_in1,
        Din2 => VN686_in2,
        Din3 => VN686_in3,
        Din4 => VN686_in4,
        Din5 => VN686_in5,
        VN2CN0_bit => VN_data_out(4116),
        VN2CN1_bit => VN_data_out(4117),
        VN2CN2_bit => VN_data_out(4118),
        VN2CN3_bit => VN_data_out(4119),
        VN2CN4_bit => VN_data_out(4120),
        VN2CN5_bit => VN_data_out(4121),
        VN2CN0_sign => VN_sign_out(4116),
        VN2CN1_sign => VN_sign_out(4117),
        VN2CN2_sign => VN_sign_out(4118),
        VN2CN3_sign => VN_sign_out(4119),
        VN2CN4_sign => VN_sign_out(4120),
        VN2CN5_sign => VN_sign_out(4121),
        codeword => codeword(686),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN687 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4127 downto 4122),
        Din0 => VN687_in0,
        Din1 => VN687_in1,
        Din2 => VN687_in2,
        Din3 => VN687_in3,
        Din4 => VN687_in4,
        Din5 => VN687_in5,
        VN2CN0_bit => VN_data_out(4122),
        VN2CN1_bit => VN_data_out(4123),
        VN2CN2_bit => VN_data_out(4124),
        VN2CN3_bit => VN_data_out(4125),
        VN2CN4_bit => VN_data_out(4126),
        VN2CN5_bit => VN_data_out(4127),
        VN2CN0_sign => VN_sign_out(4122),
        VN2CN1_sign => VN_sign_out(4123),
        VN2CN2_sign => VN_sign_out(4124),
        VN2CN3_sign => VN_sign_out(4125),
        VN2CN4_sign => VN_sign_out(4126),
        VN2CN5_sign => VN_sign_out(4127),
        codeword => codeword(687),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN688 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4133 downto 4128),
        Din0 => VN688_in0,
        Din1 => VN688_in1,
        Din2 => VN688_in2,
        Din3 => VN688_in3,
        Din4 => VN688_in4,
        Din5 => VN688_in5,
        VN2CN0_bit => VN_data_out(4128),
        VN2CN1_bit => VN_data_out(4129),
        VN2CN2_bit => VN_data_out(4130),
        VN2CN3_bit => VN_data_out(4131),
        VN2CN4_bit => VN_data_out(4132),
        VN2CN5_bit => VN_data_out(4133),
        VN2CN0_sign => VN_sign_out(4128),
        VN2CN1_sign => VN_sign_out(4129),
        VN2CN2_sign => VN_sign_out(4130),
        VN2CN3_sign => VN_sign_out(4131),
        VN2CN4_sign => VN_sign_out(4132),
        VN2CN5_sign => VN_sign_out(4133),
        codeword => codeword(688),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN689 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4139 downto 4134),
        Din0 => VN689_in0,
        Din1 => VN689_in1,
        Din2 => VN689_in2,
        Din3 => VN689_in3,
        Din4 => VN689_in4,
        Din5 => VN689_in5,
        VN2CN0_bit => VN_data_out(4134),
        VN2CN1_bit => VN_data_out(4135),
        VN2CN2_bit => VN_data_out(4136),
        VN2CN3_bit => VN_data_out(4137),
        VN2CN4_bit => VN_data_out(4138),
        VN2CN5_bit => VN_data_out(4139),
        VN2CN0_sign => VN_sign_out(4134),
        VN2CN1_sign => VN_sign_out(4135),
        VN2CN2_sign => VN_sign_out(4136),
        VN2CN3_sign => VN_sign_out(4137),
        VN2CN4_sign => VN_sign_out(4138),
        VN2CN5_sign => VN_sign_out(4139),
        codeword => codeword(689),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN690 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4145 downto 4140),
        Din0 => VN690_in0,
        Din1 => VN690_in1,
        Din2 => VN690_in2,
        Din3 => VN690_in3,
        Din4 => VN690_in4,
        Din5 => VN690_in5,
        VN2CN0_bit => VN_data_out(4140),
        VN2CN1_bit => VN_data_out(4141),
        VN2CN2_bit => VN_data_out(4142),
        VN2CN3_bit => VN_data_out(4143),
        VN2CN4_bit => VN_data_out(4144),
        VN2CN5_bit => VN_data_out(4145),
        VN2CN0_sign => VN_sign_out(4140),
        VN2CN1_sign => VN_sign_out(4141),
        VN2CN2_sign => VN_sign_out(4142),
        VN2CN3_sign => VN_sign_out(4143),
        VN2CN4_sign => VN_sign_out(4144),
        VN2CN5_sign => VN_sign_out(4145),
        codeword => codeword(690),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN691 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4151 downto 4146),
        Din0 => VN691_in0,
        Din1 => VN691_in1,
        Din2 => VN691_in2,
        Din3 => VN691_in3,
        Din4 => VN691_in4,
        Din5 => VN691_in5,
        VN2CN0_bit => VN_data_out(4146),
        VN2CN1_bit => VN_data_out(4147),
        VN2CN2_bit => VN_data_out(4148),
        VN2CN3_bit => VN_data_out(4149),
        VN2CN4_bit => VN_data_out(4150),
        VN2CN5_bit => VN_data_out(4151),
        VN2CN0_sign => VN_sign_out(4146),
        VN2CN1_sign => VN_sign_out(4147),
        VN2CN2_sign => VN_sign_out(4148),
        VN2CN3_sign => VN_sign_out(4149),
        VN2CN4_sign => VN_sign_out(4150),
        VN2CN5_sign => VN_sign_out(4151),
        codeword => codeword(691),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN692 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4157 downto 4152),
        Din0 => VN692_in0,
        Din1 => VN692_in1,
        Din2 => VN692_in2,
        Din3 => VN692_in3,
        Din4 => VN692_in4,
        Din5 => VN692_in5,
        VN2CN0_bit => VN_data_out(4152),
        VN2CN1_bit => VN_data_out(4153),
        VN2CN2_bit => VN_data_out(4154),
        VN2CN3_bit => VN_data_out(4155),
        VN2CN4_bit => VN_data_out(4156),
        VN2CN5_bit => VN_data_out(4157),
        VN2CN0_sign => VN_sign_out(4152),
        VN2CN1_sign => VN_sign_out(4153),
        VN2CN2_sign => VN_sign_out(4154),
        VN2CN3_sign => VN_sign_out(4155),
        VN2CN4_sign => VN_sign_out(4156),
        VN2CN5_sign => VN_sign_out(4157),
        codeword => codeword(692),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN693 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4163 downto 4158),
        Din0 => VN693_in0,
        Din1 => VN693_in1,
        Din2 => VN693_in2,
        Din3 => VN693_in3,
        Din4 => VN693_in4,
        Din5 => VN693_in5,
        VN2CN0_bit => VN_data_out(4158),
        VN2CN1_bit => VN_data_out(4159),
        VN2CN2_bit => VN_data_out(4160),
        VN2CN3_bit => VN_data_out(4161),
        VN2CN4_bit => VN_data_out(4162),
        VN2CN5_bit => VN_data_out(4163),
        VN2CN0_sign => VN_sign_out(4158),
        VN2CN1_sign => VN_sign_out(4159),
        VN2CN2_sign => VN_sign_out(4160),
        VN2CN3_sign => VN_sign_out(4161),
        VN2CN4_sign => VN_sign_out(4162),
        VN2CN5_sign => VN_sign_out(4163),
        codeword => codeword(693),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN694 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4169 downto 4164),
        Din0 => VN694_in0,
        Din1 => VN694_in1,
        Din2 => VN694_in2,
        Din3 => VN694_in3,
        Din4 => VN694_in4,
        Din5 => VN694_in5,
        VN2CN0_bit => VN_data_out(4164),
        VN2CN1_bit => VN_data_out(4165),
        VN2CN2_bit => VN_data_out(4166),
        VN2CN3_bit => VN_data_out(4167),
        VN2CN4_bit => VN_data_out(4168),
        VN2CN5_bit => VN_data_out(4169),
        VN2CN0_sign => VN_sign_out(4164),
        VN2CN1_sign => VN_sign_out(4165),
        VN2CN2_sign => VN_sign_out(4166),
        VN2CN3_sign => VN_sign_out(4167),
        VN2CN4_sign => VN_sign_out(4168),
        VN2CN5_sign => VN_sign_out(4169),
        codeword => codeword(694),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN695 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4175 downto 4170),
        Din0 => VN695_in0,
        Din1 => VN695_in1,
        Din2 => VN695_in2,
        Din3 => VN695_in3,
        Din4 => VN695_in4,
        Din5 => VN695_in5,
        VN2CN0_bit => VN_data_out(4170),
        VN2CN1_bit => VN_data_out(4171),
        VN2CN2_bit => VN_data_out(4172),
        VN2CN3_bit => VN_data_out(4173),
        VN2CN4_bit => VN_data_out(4174),
        VN2CN5_bit => VN_data_out(4175),
        VN2CN0_sign => VN_sign_out(4170),
        VN2CN1_sign => VN_sign_out(4171),
        VN2CN2_sign => VN_sign_out(4172),
        VN2CN3_sign => VN_sign_out(4173),
        VN2CN4_sign => VN_sign_out(4174),
        VN2CN5_sign => VN_sign_out(4175),
        codeword => codeword(695),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN696 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4181 downto 4176),
        Din0 => VN696_in0,
        Din1 => VN696_in1,
        Din2 => VN696_in2,
        Din3 => VN696_in3,
        Din4 => VN696_in4,
        Din5 => VN696_in5,
        VN2CN0_bit => VN_data_out(4176),
        VN2CN1_bit => VN_data_out(4177),
        VN2CN2_bit => VN_data_out(4178),
        VN2CN3_bit => VN_data_out(4179),
        VN2CN4_bit => VN_data_out(4180),
        VN2CN5_bit => VN_data_out(4181),
        VN2CN0_sign => VN_sign_out(4176),
        VN2CN1_sign => VN_sign_out(4177),
        VN2CN2_sign => VN_sign_out(4178),
        VN2CN3_sign => VN_sign_out(4179),
        VN2CN4_sign => VN_sign_out(4180),
        VN2CN5_sign => VN_sign_out(4181),
        codeword => codeword(696),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN697 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4187 downto 4182),
        Din0 => VN697_in0,
        Din1 => VN697_in1,
        Din2 => VN697_in2,
        Din3 => VN697_in3,
        Din4 => VN697_in4,
        Din5 => VN697_in5,
        VN2CN0_bit => VN_data_out(4182),
        VN2CN1_bit => VN_data_out(4183),
        VN2CN2_bit => VN_data_out(4184),
        VN2CN3_bit => VN_data_out(4185),
        VN2CN4_bit => VN_data_out(4186),
        VN2CN5_bit => VN_data_out(4187),
        VN2CN0_sign => VN_sign_out(4182),
        VN2CN1_sign => VN_sign_out(4183),
        VN2CN2_sign => VN_sign_out(4184),
        VN2CN3_sign => VN_sign_out(4185),
        VN2CN4_sign => VN_sign_out(4186),
        VN2CN5_sign => VN_sign_out(4187),
        codeword => codeword(697),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN698 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4193 downto 4188),
        Din0 => VN698_in0,
        Din1 => VN698_in1,
        Din2 => VN698_in2,
        Din3 => VN698_in3,
        Din4 => VN698_in4,
        Din5 => VN698_in5,
        VN2CN0_bit => VN_data_out(4188),
        VN2CN1_bit => VN_data_out(4189),
        VN2CN2_bit => VN_data_out(4190),
        VN2CN3_bit => VN_data_out(4191),
        VN2CN4_bit => VN_data_out(4192),
        VN2CN5_bit => VN_data_out(4193),
        VN2CN0_sign => VN_sign_out(4188),
        VN2CN1_sign => VN_sign_out(4189),
        VN2CN2_sign => VN_sign_out(4190),
        VN2CN3_sign => VN_sign_out(4191),
        VN2CN4_sign => VN_sign_out(4192),
        VN2CN5_sign => VN_sign_out(4193),
        codeword => codeword(698),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN699 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4199 downto 4194),
        Din0 => VN699_in0,
        Din1 => VN699_in1,
        Din2 => VN699_in2,
        Din3 => VN699_in3,
        Din4 => VN699_in4,
        Din5 => VN699_in5,
        VN2CN0_bit => VN_data_out(4194),
        VN2CN1_bit => VN_data_out(4195),
        VN2CN2_bit => VN_data_out(4196),
        VN2CN3_bit => VN_data_out(4197),
        VN2CN4_bit => VN_data_out(4198),
        VN2CN5_bit => VN_data_out(4199),
        VN2CN0_sign => VN_sign_out(4194),
        VN2CN1_sign => VN_sign_out(4195),
        VN2CN2_sign => VN_sign_out(4196),
        VN2CN3_sign => VN_sign_out(4197),
        VN2CN4_sign => VN_sign_out(4198),
        VN2CN5_sign => VN_sign_out(4199),
        codeword => codeword(699),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN700 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4205 downto 4200),
        Din0 => VN700_in0,
        Din1 => VN700_in1,
        Din2 => VN700_in2,
        Din3 => VN700_in3,
        Din4 => VN700_in4,
        Din5 => VN700_in5,
        VN2CN0_bit => VN_data_out(4200),
        VN2CN1_bit => VN_data_out(4201),
        VN2CN2_bit => VN_data_out(4202),
        VN2CN3_bit => VN_data_out(4203),
        VN2CN4_bit => VN_data_out(4204),
        VN2CN5_bit => VN_data_out(4205),
        VN2CN0_sign => VN_sign_out(4200),
        VN2CN1_sign => VN_sign_out(4201),
        VN2CN2_sign => VN_sign_out(4202),
        VN2CN3_sign => VN_sign_out(4203),
        VN2CN4_sign => VN_sign_out(4204),
        VN2CN5_sign => VN_sign_out(4205),
        codeword => codeword(700),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN701 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4211 downto 4206),
        Din0 => VN701_in0,
        Din1 => VN701_in1,
        Din2 => VN701_in2,
        Din3 => VN701_in3,
        Din4 => VN701_in4,
        Din5 => VN701_in5,
        VN2CN0_bit => VN_data_out(4206),
        VN2CN1_bit => VN_data_out(4207),
        VN2CN2_bit => VN_data_out(4208),
        VN2CN3_bit => VN_data_out(4209),
        VN2CN4_bit => VN_data_out(4210),
        VN2CN5_bit => VN_data_out(4211),
        VN2CN0_sign => VN_sign_out(4206),
        VN2CN1_sign => VN_sign_out(4207),
        VN2CN2_sign => VN_sign_out(4208),
        VN2CN3_sign => VN_sign_out(4209),
        VN2CN4_sign => VN_sign_out(4210),
        VN2CN5_sign => VN_sign_out(4211),
        codeword => codeword(701),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN702 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4217 downto 4212),
        Din0 => VN702_in0,
        Din1 => VN702_in1,
        Din2 => VN702_in2,
        Din3 => VN702_in3,
        Din4 => VN702_in4,
        Din5 => VN702_in5,
        VN2CN0_bit => VN_data_out(4212),
        VN2CN1_bit => VN_data_out(4213),
        VN2CN2_bit => VN_data_out(4214),
        VN2CN3_bit => VN_data_out(4215),
        VN2CN4_bit => VN_data_out(4216),
        VN2CN5_bit => VN_data_out(4217),
        VN2CN0_sign => VN_sign_out(4212),
        VN2CN1_sign => VN_sign_out(4213),
        VN2CN2_sign => VN_sign_out(4214),
        VN2CN3_sign => VN_sign_out(4215),
        VN2CN4_sign => VN_sign_out(4216),
        VN2CN5_sign => VN_sign_out(4217),
        codeword => codeword(702),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN703 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4223 downto 4218),
        Din0 => VN703_in0,
        Din1 => VN703_in1,
        Din2 => VN703_in2,
        Din3 => VN703_in3,
        Din4 => VN703_in4,
        Din5 => VN703_in5,
        VN2CN0_bit => VN_data_out(4218),
        VN2CN1_bit => VN_data_out(4219),
        VN2CN2_bit => VN_data_out(4220),
        VN2CN3_bit => VN_data_out(4221),
        VN2CN4_bit => VN_data_out(4222),
        VN2CN5_bit => VN_data_out(4223),
        VN2CN0_sign => VN_sign_out(4218),
        VN2CN1_sign => VN_sign_out(4219),
        VN2CN2_sign => VN_sign_out(4220),
        VN2CN3_sign => VN_sign_out(4221),
        VN2CN4_sign => VN_sign_out(4222),
        VN2CN5_sign => VN_sign_out(4223),
        codeword => codeword(703),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN704 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4229 downto 4224),
        Din0 => VN704_in0,
        Din1 => VN704_in1,
        Din2 => VN704_in2,
        Din3 => VN704_in3,
        Din4 => VN704_in4,
        Din5 => VN704_in5,
        VN2CN0_bit => VN_data_out(4224),
        VN2CN1_bit => VN_data_out(4225),
        VN2CN2_bit => VN_data_out(4226),
        VN2CN3_bit => VN_data_out(4227),
        VN2CN4_bit => VN_data_out(4228),
        VN2CN5_bit => VN_data_out(4229),
        VN2CN0_sign => VN_sign_out(4224),
        VN2CN1_sign => VN_sign_out(4225),
        VN2CN2_sign => VN_sign_out(4226),
        VN2CN3_sign => VN_sign_out(4227),
        VN2CN4_sign => VN_sign_out(4228),
        VN2CN5_sign => VN_sign_out(4229),
        codeword => codeword(704),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN705 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4235 downto 4230),
        Din0 => VN705_in0,
        Din1 => VN705_in1,
        Din2 => VN705_in2,
        Din3 => VN705_in3,
        Din4 => VN705_in4,
        Din5 => VN705_in5,
        VN2CN0_bit => VN_data_out(4230),
        VN2CN1_bit => VN_data_out(4231),
        VN2CN2_bit => VN_data_out(4232),
        VN2CN3_bit => VN_data_out(4233),
        VN2CN4_bit => VN_data_out(4234),
        VN2CN5_bit => VN_data_out(4235),
        VN2CN0_sign => VN_sign_out(4230),
        VN2CN1_sign => VN_sign_out(4231),
        VN2CN2_sign => VN_sign_out(4232),
        VN2CN3_sign => VN_sign_out(4233),
        VN2CN4_sign => VN_sign_out(4234),
        VN2CN5_sign => VN_sign_out(4235),
        codeword => codeword(705),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN706 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4241 downto 4236),
        Din0 => VN706_in0,
        Din1 => VN706_in1,
        Din2 => VN706_in2,
        Din3 => VN706_in3,
        Din4 => VN706_in4,
        Din5 => VN706_in5,
        VN2CN0_bit => VN_data_out(4236),
        VN2CN1_bit => VN_data_out(4237),
        VN2CN2_bit => VN_data_out(4238),
        VN2CN3_bit => VN_data_out(4239),
        VN2CN4_bit => VN_data_out(4240),
        VN2CN5_bit => VN_data_out(4241),
        VN2CN0_sign => VN_sign_out(4236),
        VN2CN1_sign => VN_sign_out(4237),
        VN2CN2_sign => VN_sign_out(4238),
        VN2CN3_sign => VN_sign_out(4239),
        VN2CN4_sign => VN_sign_out(4240),
        VN2CN5_sign => VN_sign_out(4241),
        codeword => codeword(706),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN707 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4247 downto 4242),
        Din0 => VN707_in0,
        Din1 => VN707_in1,
        Din2 => VN707_in2,
        Din3 => VN707_in3,
        Din4 => VN707_in4,
        Din5 => VN707_in5,
        VN2CN0_bit => VN_data_out(4242),
        VN2CN1_bit => VN_data_out(4243),
        VN2CN2_bit => VN_data_out(4244),
        VN2CN3_bit => VN_data_out(4245),
        VN2CN4_bit => VN_data_out(4246),
        VN2CN5_bit => VN_data_out(4247),
        VN2CN0_sign => VN_sign_out(4242),
        VN2CN1_sign => VN_sign_out(4243),
        VN2CN2_sign => VN_sign_out(4244),
        VN2CN3_sign => VN_sign_out(4245),
        VN2CN4_sign => VN_sign_out(4246),
        VN2CN5_sign => VN_sign_out(4247),
        codeword => codeword(707),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN708 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4253 downto 4248),
        Din0 => VN708_in0,
        Din1 => VN708_in1,
        Din2 => VN708_in2,
        Din3 => VN708_in3,
        Din4 => VN708_in4,
        Din5 => VN708_in5,
        VN2CN0_bit => VN_data_out(4248),
        VN2CN1_bit => VN_data_out(4249),
        VN2CN2_bit => VN_data_out(4250),
        VN2CN3_bit => VN_data_out(4251),
        VN2CN4_bit => VN_data_out(4252),
        VN2CN5_bit => VN_data_out(4253),
        VN2CN0_sign => VN_sign_out(4248),
        VN2CN1_sign => VN_sign_out(4249),
        VN2CN2_sign => VN_sign_out(4250),
        VN2CN3_sign => VN_sign_out(4251),
        VN2CN4_sign => VN_sign_out(4252),
        VN2CN5_sign => VN_sign_out(4253),
        codeword => codeword(708),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN709 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4259 downto 4254),
        Din0 => VN709_in0,
        Din1 => VN709_in1,
        Din2 => VN709_in2,
        Din3 => VN709_in3,
        Din4 => VN709_in4,
        Din5 => VN709_in5,
        VN2CN0_bit => VN_data_out(4254),
        VN2CN1_bit => VN_data_out(4255),
        VN2CN2_bit => VN_data_out(4256),
        VN2CN3_bit => VN_data_out(4257),
        VN2CN4_bit => VN_data_out(4258),
        VN2CN5_bit => VN_data_out(4259),
        VN2CN0_sign => VN_sign_out(4254),
        VN2CN1_sign => VN_sign_out(4255),
        VN2CN2_sign => VN_sign_out(4256),
        VN2CN3_sign => VN_sign_out(4257),
        VN2CN4_sign => VN_sign_out(4258),
        VN2CN5_sign => VN_sign_out(4259),
        codeword => codeword(709),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN710 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4265 downto 4260),
        Din0 => VN710_in0,
        Din1 => VN710_in1,
        Din2 => VN710_in2,
        Din3 => VN710_in3,
        Din4 => VN710_in4,
        Din5 => VN710_in5,
        VN2CN0_bit => VN_data_out(4260),
        VN2CN1_bit => VN_data_out(4261),
        VN2CN2_bit => VN_data_out(4262),
        VN2CN3_bit => VN_data_out(4263),
        VN2CN4_bit => VN_data_out(4264),
        VN2CN5_bit => VN_data_out(4265),
        VN2CN0_sign => VN_sign_out(4260),
        VN2CN1_sign => VN_sign_out(4261),
        VN2CN2_sign => VN_sign_out(4262),
        VN2CN3_sign => VN_sign_out(4263),
        VN2CN4_sign => VN_sign_out(4264),
        VN2CN5_sign => VN_sign_out(4265),
        codeword => codeword(710),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN711 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4271 downto 4266),
        Din0 => VN711_in0,
        Din1 => VN711_in1,
        Din2 => VN711_in2,
        Din3 => VN711_in3,
        Din4 => VN711_in4,
        Din5 => VN711_in5,
        VN2CN0_bit => VN_data_out(4266),
        VN2CN1_bit => VN_data_out(4267),
        VN2CN2_bit => VN_data_out(4268),
        VN2CN3_bit => VN_data_out(4269),
        VN2CN4_bit => VN_data_out(4270),
        VN2CN5_bit => VN_data_out(4271),
        VN2CN0_sign => VN_sign_out(4266),
        VN2CN1_sign => VN_sign_out(4267),
        VN2CN2_sign => VN_sign_out(4268),
        VN2CN3_sign => VN_sign_out(4269),
        VN2CN4_sign => VN_sign_out(4270),
        VN2CN5_sign => VN_sign_out(4271),
        codeword => codeword(711),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN712 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4277 downto 4272),
        Din0 => VN712_in0,
        Din1 => VN712_in1,
        Din2 => VN712_in2,
        Din3 => VN712_in3,
        Din4 => VN712_in4,
        Din5 => VN712_in5,
        VN2CN0_bit => VN_data_out(4272),
        VN2CN1_bit => VN_data_out(4273),
        VN2CN2_bit => VN_data_out(4274),
        VN2CN3_bit => VN_data_out(4275),
        VN2CN4_bit => VN_data_out(4276),
        VN2CN5_bit => VN_data_out(4277),
        VN2CN0_sign => VN_sign_out(4272),
        VN2CN1_sign => VN_sign_out(4273),
        VN2CN2_sign => VN_sign_out(4274),
        VN2CN3_sign => VN_sign_out(4275),
        VN2CN4_sign => VN_sign_out(4276),
        VN2CN5_sign => VN_sign_out(4277),
        codeword => codeword(712),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN713 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4283 downto 4278),
        Din0 => VN713_in0,
        Din1 => VN713_in1,
        Din2 => VN713_in2,
        Din3 => VN713_in3,
        Din4 => VN713_in4,
        Din5 => VN713_in5,
        VN2CN0_bit => VN_data_out(4278),
        VN2CN1_bit => VN_data_out(4279),
        VN2CN2_bit => VN_data_out(4280),
        VN2CN3_bit => VN_data_out(4281),
        VN2CN4_bit => VN_data_out(4282),
        VN2CN5_bit => VN_data_out(4283),
        VN2CN0_sign => VN_sign_out(4278),
        VN2CN1_sign => VN_sign_out(4279),
        VN2CN2_sign => VN_sign_out(4280),
        VN2CN3_sign => VN_sign_out(4281),
        VN2CN4_sign => VN_sign_out(4282),
        VN2CN5_sign => VN_sign_out(4283),
        codeword => codeword(713),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN714 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4289 downto 4284),
        Din0 => VN714_in0,
        Din1 => VN714_in1,
        Din2 => VN714_in2,
        Din3 => VN714_in3,
        Din4 => VN714_in4,
        Din5 => VN714_in5,
        VN2CN0_bit => VN_data_out(4284),
        VN2CN1_bit => VN_data_out(4285),
        VN2CN2_bit => VN_data_out(4286),
        VN2CN3_bit => VN_data_out(4287),
        VN2CN4_bit => VN_data_out(4288),
        VN2CN5_bit => VN_data_out(4289),
        VN2CN0_sign => VN_sign_out(4284),
        VN2CN1_sign => VN_sign_out(4285),
        VN2CN2_sign => VN_sign_out(4286),
        VN2CN3_sign => VN_sign_out(4287),
        VN2CN4_sign => VN_sign_out(4288),
        VN2CN5_sign => VN_sign_out(4289),
        codeword => codeword(714),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN715 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4295 downto 4290),
        Din0 => VN715_in0,
        Din1 => VN715_in1,
        Din2 => VN715_in2,
        Din3 => VN715_in3,
        Din4 => VN715_in4,
        Din5 => VN715_in5,
        VN2CN0_bit => VN_data_out(4290),
        VN2CN1_bit => VN_data_out(4291),
        VN2CN2_bit => VN_data_out(4292),
        VN2CN3_bit => VN_data_out(4293),
        VN2CN4_bit => VN_data_out(4294),
        VN2CN5_bit => VN_data_out(4295),
        VN2CN0_sign => VN_sign_out(4290),
        VN2CN1_sign => VN_sign_out(4291),
        VN2CN2_sign => VN_sign_out(4292),
        VN2CN3_sign => VN_sign_out(4293),
        VN2CN4_sign => VN_sign_out(4294),
        VN2CN5_sign => VN_sign_out(4295),
        codeword => codeword(715),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN716 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4301 downto 4296),
        Din0 => VN716_in0,
        Din1 => VN716_in1,
        Din2 => VN716_in2,
        Din3 => VN716_in3,
        Din4 => VN716_in4,
        Din5 => VN716_in5,
        VN2CN0_bit => VN_data_out(4296),
        VN2CN1_bit => VN_data_out(4297),
        VN2CN2_bit => VN_data_out(4298),
        VN2CN3_bit => VN_data_out(4299),
        VN2CN4_bit => VN_data_out(4300),
        VN2CN5_bit => VN_data_out(4301),
        VN2CN0_sign => VN_sign_out(4296),
        VN2CN1_sign => VN_sign_out(4297),
        VN2CN2_sign => VN_sign_out(4298),
        VN2CN3_sign => VN_sign_out(4299),
        VN2CN4_sign => VN_sign_out(4300),
        VN2CN5_sign => VN_sign_out(4301),
        codeword => codeword(716),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN717 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4307 downto 4302),
        Din0 => VN717_in0,
        Din1 => VN717_in1,
        Din2 => VN717_in2,
        Din3 => VN717_in3,
        Din4 => VN717_in4,
        Din5 => VN717_in5,
        VN2CN0_bit => VN_data_out(4302),
        VN2CN1_bit => VN_data_out(4303),
        VN2CN2_bit => VN_data_out(4304),
        VN2CN3_bit => VN_data_out(4305),
        VN2CN4_bit => VN_data_out(4306),
        VN2CN5_bit => VN_data_out(4307),
        VN2CN0_sign => VN_sign_out(4302),
        VN2CN1_sign => VN_sign_out(4303),
        VN2CN2_sign => VN_sign_out(4304),
        VN2CN3_sign => VN_sign_out(4305),
        VN2CN4_sign => VN_sign_out(4306),
        VN2CN5_sign => VN_sign_out(4307),
        codeword => codeword(717),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN718 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4313 downto 4308),
        Din0 => VN718_in0,
        Din1 => VN718_in1,
        Din2 => VN718_in2,
        Din3 => VN718_in3,
        Din4 => VN718_in4,
        Din5 => VN718_in5,
        VN2CN0_bit => VN_data_out(4308),
        VN2CN1_bit => VN_data_out(4309),
        VN2CN2_bit => VN_data_out(4310),
        VN2CN3_bit => VN_data_out(4311),
        VN2CN4_bit => VN_data_out(4312),
        VN2CN5_bit => VN_data_out(4313),
        VN2CN0_sign => VN_sign_out(4308),
        VN2CN1_sign => VN_sign_out(4309),
        VN2CN2_sign => VN_sign_out(4310),
        VN2CN3_sign => VN_sign_out(4311),
        VN2CN4_sign => VN_sign_out(4312),
        VN2CN5_sign => VN_sign_out(4313),
        codeword => codeword(718),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN719 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4319 downto 4314),
        Din0 => VN719_in0,
        Din1 => VN719_in1,
        Din2 => VN719_in2,
        Din3 => VN719_in3,
        Din4 => VN719_in4,
        Din5 => VN719_in5,
        VN2CN0_bit => VN_data_out(4314),
        VN2CN1_bit => VN_data_out(4315),
        VN2CN2_bit => VN_data_out(4316),
        VN2CN3_bit => VN_data_out(4317),
        VN2CN4_bit => VN_data_out(4318),
        VN2CN5_bit => VN_data_out(4319),
        VN2CN0_sign => VN_sign_out(4314),
        VN2CN1_sign => VN_sign_out(4315),
        VN2CN2_sign => VN_sign_out(4316),
        VN2CN3_sign => VN_sign_out(4317),
        VN2CN4_sign => VN_sign_out(4318),
        VN2CN5_sign => VN_sign_out(4319),
        codeword => codeword(719),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN720 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4325 downto 4320),
        Din0 => VN720_in0,
        Din1 => VN720_in1,
        Din2 => VN720_in2,
        Din3 => VN720_in3,
        Din4 => VN720_in4,
        Din5 => VN720_in5,
        VN2CN0_bit => VN_data_out(4320),
        VN2CN1_bit => VN_data_out(4321),
        VN2CN2_bit => VN_data_out(4322),
        VN2CN3_bit => VN_data_out(4323),
        VN2CN4_bit => VN_data_out(4324),
        VN2CN5_bit => VN_data_out(4325),
        VN2CN0_sign => VN_sign_out(4320),
        VN2CN1_sign => VN_sign_out(4321),
        VN2CN2_sign => VN_sign_out(4322),
        VN2CN3_sign => VN_sign_out(4323),
        VN2CN4_sign => VN_sign_out(4324),
        VN2CN5_sign => VN_sign_out(4325),
        codeword => codeword(720),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN721 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4331 downto 4326),
        Din0 => VN721_in0,
        Din1 => VN721_in1,
        Din2 => VN721_in2,
        Din3 => VN721_in3,
        Din4 => VN721_in4,
        Din5 => VN721_in5,
        VN2CN0_bit => VN_data_out(4326),
        VN2CN1_bit => VN_data_out(4327),
        VN2CN2_bit => VN_data_out(4328),
        VN2CN3_bit => VN_data_out(4329),
        VN2CN4_bit => VN_data_out(4330),
        VN2CN5_bit => VN_data_out(4331),
        VN2CN0_sign => VN_sign_out(4326),
        VN2CN1_sign => VN_sign_out(4327),
        VN2CN2_sign => VN_sign_out(4328),
        VN2CN3_sign => VN_sign_out(4329),
        VN2CN4_sign => VN_sign_out(4330),
        VN2CN5_sign => VN_sign_out(4331),
        codeword => codeword(721),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN722 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4337 downto 4332),
        Din0 => VN722_in0,
        Din1 => VN722_in1,
        Din2 => VN722_in2,
        Din3 => VN722_in3,
        Din4 => VN722_in4,
        Din5 => VN722_in5,
        VN2CN0_bit => VN_data_out(4332),
        VN2CN1_bit => VN_data_out(4333),
        VN2CN2_bit => VN_data_out(4334),
        VN2CN3_bit => VN_data_out(4335),
        VN2CN4_bit => VN_data_out(4336),
        VN2CN5_bit => VN_data_out(4337),
        VN2CN0_sign => VN_sign_out(4332),
        VN2CN1_sign => VN_sign_out(4333),
        VN2CN2_sign => VN_sign_out(4334),
        VN2CN3_sign => VN_sign_out(4335),
        VN2CN4_sign => VN_sign_out(4336),
        VN2CN5_sign => VN_sign_out(4337),
        codeword => codeword(722),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN723 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4343 downto 4338),
        Din0 => VN723_in0,
        Din1 => VN723_in1,
        Din2 => VN723_in2,
        Din3 => VN723_in3,
        Din4 => VN723_in4,
        Din5 => VN723_in5,
        VN2CN0_bit => VN_data_out(4338),
        VN2CN1_bit => VN_data_out(4339),
        VN2CN2_bit => VN_data_out(4340),
        VN2CN3_bit => VN_data_out(4341),
        VN2CN4_bit => VN_data_out(4342),
        VN2CN5_bit => VN_data_out(4343),
        VN2CN0_sign => VN_sign_out(4338),
        VN2CN1_sign => VN_sign_out(4339),
        VN2CN2_sign => VN_sign_out(4340),
        VN2CN3_sign => VN_sign_out(4341),
        VN2CN4_sign => VN_sign_out(4342),
        VN2CN5_sign => VN_sign_out(4343),
        codeword => codeword(723),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN724 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4349 downto 4344),
        Din0 => VN724_in0,
        Din1 => VN724_in1,
        Din2 => VN724_in2,
        Din3 => VN724_in3,
        Din4 => VN724_in4,
        Din5 => VN724_in5,
        VN2CN0_bit => VN_data_out(4344),
        VN2CN1_bit => VN_data_out(4345),
        VN2CN2_bit => VN_data_out(4346),
        VN2CN3_bit => VN_data_out(4347),
        VN2CN4_bit => VN_data_out(4348),
        VN2CN5_bit => VN_data_out(4349),
        VN2CN0_sign => VN_sign_out(4344),
        VN2CN1_sign => VN_sign_out(4345),
        VN2CN2_sign => VN_sign_out(4346),
        VN2CN3_sign => VN_sign_out(4347),
        VN2CN4_sign => VN_sign_out(4348),
        VN2CN5_sign => VN_sign_out(4349),
        codeword => codeword(724),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN725 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4355 downto 4350),
        Din0 => VN725_in0,
        Din1 => VN725_in1,
        Din2 => VN725_in2,
        Din3 => VN725_in3,
        Din4 => VN725_in4,
        Din5 => VN725_in5,
        VN2CN0_bit => VN_data_out(4350),
        VN2CN1_bit => VN_data_out(4351),
        VN2CN2_bit => VN_data_out(4352),
        VN2CN3_bit => VN_data_out(4353),
        VN2CN4_bit => VN_data_out(4354),
        VN2CN5_bit => VN_data_out(4355),
        VN2CN0_sign => VN_sign_out(4350),
        VN2CN1_sign => VN_sign_out(4351),
        VN2CN2_sign => VN_sign_out(4352),
        VN2CN3_sign => VN_sign_out(4353),
        VN2CN4_sign => VN_sign_out(4354),
        VN2CN5_sign => VN_sign_out(4355),
        codeword => codeword(725),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN726 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4361 downto 4356),
        Din0 => VN726_in0,
        Din1 => VN726_in1,
        Din2 => VN726_in2,
        Din3 => VN726_in3,
        Din4 => VN726_in4,
        Din5 => VN726_in5,
        VN2CN0_bit => VN_data_out(4356),
        VN2CN1_bit => VN_data_out(4357),
        VN2CN2_bit => VN_data_out(4358),
        VN2CN3_bit => VN_data_out(4359),
        VN2CN4_bit => VN_data_out(4360),
        VN2CN5_bit => VN_data_out(4361),
        VN2CN0_sign => VN_sign_out(4356),
        VN2CN1_sign => VN_sign_out(4357),
        VN2CN2_sign => VN_sign_out(4358),
        VN2CN3_sign => VN_sign_out(4359),
        VN2CN4_sign => VN_sign_out(4360),
        VN2CN5_sign => VN_sign_out(4361),
        codeword => codeword(726),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN727 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4367 downto 4362),
        Din0 => VN727_in0,
        Din1 => VN727_in1,
        Din2 => VN727_in2,
        Din3 => VN727_in3,
        Din4 => VN727_in4,
        Din5 => VN727_in5,
        VN2CN0_bit => VN_data_out(4362),
        VN2CN1_bit => VN_data_out(4363),
        VN2CN2_bit => VN_data_out(4364),
        VN2CN3_bit => VN_data_out(4365),
        VN2CN4_bit => VN_data_out(4366),
        VN2CN5_bit => VN_data_out(4367),
        VN2CN0_sign => VN_sign_out(4362),
        VN2CN1_sign => VN_sign_out(4363),
        VN2CN2_sign => VN_sign_out(4364),
        VN2CN3_sign => VN_sign_out(4365),
        VN2CN4_sign => VN_sign_out(4366),
        VN2CN5_sign => VN_sign_out(4367),
        codeword => codeword(727),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN728 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4373 downto 4368),
        Din0 => VN728_in0,
        Din1 => VN728_in1,
        Din2 => VN728_in2,
        Din3 => VN728_in3,
        Din4 => VN728_in4,
        Din5 => VN728_in5,
        VN2CN0_bit => VN_data_out(4368),
        VN2CN1_bit => VN_data_out(4369),
        VN2CN2_bit => VN_data_out(4370),
        VN2CN3_bit => VN_data_out(4371),
        VN2CN4_bit => VN_data_out(4372),
        VN2CN5_bit => VN_data_out(4373),
        VN2CN0_sign => VN_sign_out(4368),
        VN2CN1_sign => VN_sign_out(4369),
        VN2CN2_sign => VN_sign_out(4370),
        VN2CN3_sign => VN_sign_out(4371),
        VN2CN4_sign => VN_sign_out(4372),
        VN2CN5_sign => VN_sign_out(4373),
        codeword => codeword(728),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN729 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4379 downto 4374),
        Din0 => VN729_in0,
        Din1 => VN729_in1,
        Din2 => VN729_in2,
        Din3 => VN729_in3,
        Din4 => VN729_in4,
        Din5 => VN729_in5,
        VN2CN0_bit => VN_data_out(4374),
        VN2CN1_bit => VN_data_out(4375),
        VN2CN2_bit => VN_data_out(4376),
        VN2CN3_bit => VN_data_out(4377),
        VN2CN4_bit => VN_data_out(4378),
        VN2CN5_bit => VN_data_out(4379),
        VN2CN0_sign => VN_sign_out(4374),
        VN2CN1_sign => VN_sign_out(4375),
        VN2CN2_sign => VN_sign_out(4376),
        VN2CN3_sign => VN_sign_out(4377),
        VN2CN4_sign => VN_sign_out(4378),
        VN2CN5_sign => VN_sign_out(4379),
        codeword => codeword(729),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN730 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4385 downto 4380),
        Din0 => VN730_in0,
        Din1 => VN730_in1,
        Din2 => VN730_in2,
        Din3 => VN730_in3,
        Din4 => VN730_in4,
        Din5 => VN730_in5,
        VN2CN0_bit => VN_data_out(4380),
        VN2CN1_bit => VN_data_out(4381),
        VN2CN2_bit => VN_data_out(4382),
        VN2CN3_bit => VN_data_out(4383),
        VN2CN4_bit => VN_data_out(4384),
        VN2CN5_bit => VN_data_out(4385),
        VN2CN0_sign => VN_sign_out(4380),
        VN2CN1_sign => VN_sign_out(4381),
        VN2CN2_sign => VN_sign_out(4382),
        VN2CN3_sign => VN_sign_out(4383),
        VN2CN4_sign => VN_sign_out(4384),
        VN2CN5_sign => VN_sign_out(4385),
        codeword => codeword(730),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN731 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4391 downto 4386),
        Din0 => VN731_in0,
        Din1 => VN731_in1,
        Din2 => VN731_in2,
        Din3 => VN731_in3,
        Din4 => VN731_in4,
        Din5 => VN731_in5,
        VN2CN0_bit => VN_data_out(4386),
        VN2CN1_bit => VN_data_out(4387),
        VN2CN2_bit => VN_data_out(4388),
        VN2CN3_bit => VN_data_out(4389),
        VN2CN4_bit => VN_data_out(4390),
        VN2CN5_bit => VN_data_out(4391),
        VN2CN0_sign => VN_sign_out(4386),
        VN2CN1_sign => VN_sign_out(4387),
        VN2CN2_sign => VN_sign_out(4388),
        VN2CN3_sign => VN_sign_out(4389),
        VN2CN4_sign => VN_sign_out(4390),
        VN2CN5_sign => VN_sign_out(4391),
        codeword => codeword(731),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN732 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4397 downto 4392),
        Din0 => VN732_in0,
        Din1 => VN732_in1,
        Din2 => VN732_in2,
        Din3 => VN732_in3,
        Din4 => VN732_in4,
        Din5 => VN732_in5,
        VN2CN0_bit => VN_data_out(4392),
        VN2CN1_bit => VN_data_out(4393),
        VN2CN2_bit => VN_data_out(4394),
        VN2CN3_bit => VN_data_out(4395),
        VN2CN4_bit => VN_data_out(4396),
        VN2CN5_bit => VN_data_out(4397),
        VN2CN0_sign => VN_sign_out(4392),
        VN2CN1_sign => VN_sign_out(4393),
        VN2CN2_sign => VN_sign_out(4394),
        VN2CN3_sign => VN_sign_out(4395),
        VN2CN4_sign => VN_sign_out(4396),
        VN2CN5_sign => VN_sign_out(4397),
        codeword => codeword(732),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN733 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4403 downto 4398),
        Din0 => VN733_in0,
        Din1 => VN733_in1,
        Din2 => VN733_in2,
        Din3 => VN733_in3,
        Din4 => VN733_in4,
        Din5 => VN733_in5,
        VN2CN0_bit => VN_data_out(4398),
        VN2CN1_bit => VN_data_out(4399),
        VN2CN2_bit => VN_data_out(4400),
        VN2CN3_bit => VN_data_out(4401),
        VN2CN4_bit => VN_data_out(4402),
        VN2CN5_bit => VN_data_out(4403),
        VN2CN0_sign => VN_sign_out(4398),
        VN2CN1_sign => VN_sign_out(4399),
        VN2CN2_sign => VN_sign_out(4400),
        VN2CN3_sign => VN_sign_out(4401),
        VN2CN4_sign => VN_sign_out(4402),
        VN2CN5_sign => VN_sign_out(4403),
        codeword => codeword(733),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN734 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4409 downto 4404),
        Din0 => VN734_in0,
        Din1 => VN734_in1,
        Din2 => VN734_in2,
        Din3 => VN734_in3,
        Din4 => VN734_in4,
        Din5 => VN734_in5,
        VN2CN0_bit => VN_data_out(4404),
        VN2CN1_bit => VN_data_out(4405),
        VN2CN2_bit => VN_data_out(4406),
        VN2CN3_bit => VN_data_out(4407),
        VN2CN4_bit => VN_data_out(4408),
        VN2CN5_bit => VN_data_out(4409),
        VN2CN0_sign => VN_sign_out(4404),
        VN2CN1_sign => VN_sign_out(4405),
        VN2CN2_sign => VN_sign_out(4406),
        VN2CN3_sign => VN_sign_out(4407),
        VN2CN4_sign => VN_sign_out(4408),
        VN2CN5_sign => VN_sign_out(4409),
        codeword => codeword(734),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN735 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4415 downto 4410),
        Din0 => VN735_in0,
        Din1 => VN735_in1,
        Din2 => VN735_in2,
        Din3 => VN735_in3,
        Din4 => VN735_in4,
        Din5 => VN735_in5,
        VN2CN0_bit => VN_data_out(4410),
        VN2CN1_bit => VN_data_out(4411),
        VN2CN2_bit => VN_data_out(4412),
        VN2CN3_bit => VN_data_out(4413),
        VN2CN4_bit => VN_data_out(4414),
        VN2CN5_bit => VN_data_out(4415),
        VN2CN0_sign => VN_sign_out(4410),
        VN2CN1_sign => VN_sign_out(4411),
        VN2CN2_sign => VN_sign_out(4412),
        VN2CN3_sign => VN_sign_out(4413),
        VN2CN4_sign => VN_sign_out(4414),
        VN2CN5_sign => VN_sign_out(4415),
        codeword => codeword(735),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN736 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4421 downto 4416),
        Din0 => VN736_in0,
        Din1 => VN736_in1,
        Din2 => VN736_in2,
        Din3 => VN736_in3,
        Din4 => VN736_in4,
        Din5 => VN736_in5,
        VN2CN0_bit => VN_data_out(4416),
        VN2CN1_bit => VN_data_out(4417),
        VN2CN2_bit => VN_data_out(4418),
        VN2CN3_bit => VN_data_out(4419),
        VN2CN4_bit => VN_data_out(4420),
        VN2CN5_bit => VN_data_out(4421),
        VN2CN0_sign => VN_sign_out(4416),
        VN2CN1_sign => VN_sign_out(4417),
        VN2CN2_sign => VN_sign_out(4418),
        VN2CN3_sign => VN_sign_out(4419),
        VN2CN4_sign => VN_sign_out(4420),
        VN2CN5_sign => VN_sign_out(4421),
        codeword => codeword(736),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN737 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4427 downto 4422),
        Din0 => VN737_in0,
        Din1 => VN737_in1,
        Din2 => VN737_in2,
        Din3 => VN737_in3,
        Din4 => VN737_in4,
        Din5 => VN737_in5,
        VN2CN0_bit => VN_data_out(4422),
        VN2CN1_bit => VN_data_out(4423),
        VN2CN2_bit => VN_data_out(4424),
        VN2CN3_bit => VN_data_out(4425),
        VN2CN4_bit => VN_data_out(4426),
        VN2CN5_bit => VN_data_out(4427),
        VN2CN0_sign => VN_sign_out(4422),
        VN2CN1_sign => VN_sign_out(4423),
        VN2CN2_sign => VN_sign_out(4424),
        VN2CN3_sign => VN_sign_out(4425),
        VN2CN4_sign => VN_sign_out(4426),
        VN2CN5_sign => VN_sign_out(4427),
        codeword => codeword(737),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN738 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4433 downto 4428),
        Din0 => VN738_in0,
        Din1 => VN738_in1,
        Din2 => VN738_in2,
        Din3 => VN738_in3,
        Din4 => VN738_in4,
        Din5 => VN738_in5,
        VN2CN0_bit => VN_data_out(4428),
        VN2CN1_bit => VN_data_out(4429),
        VN2CN2_bit => VN_data_out(4430),
        VN2CN3_bit => VN_data_out(4431),
        VN2CN4_bit => VN_data_out(4432),
        VN2CN5_bit => VN_data_out(4433),
        VN2CN0_sign => VN_sign_out(4428),
        VN2CN1_sign => VN_sign_out(4429),
        VN2CN2_sign => VN_sign_out(4430),
        VN2CN3_sign => VN_sign_out(4431),
        VN2CN4_sign => VN_sign_out(4432),
        VN2CN5_sign => VN_sign_out(4433),
        codeword => codeword(738),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN739 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4439 downto 4434),
        Din0 => VN739_in0,
        Din1 => VN739_in1,
        Din2 => VN739_in2,
        Din3 => VN739_in3,
        Din4 => VN739_in4,
        Din5 => VN739_in5,
        VN2CN0_bit => VN_data_out(4434),
        VN2CN1_bit => VN_data_out(4435),
        VN2CN2_bit => VN_data_out(4436),
        VN2CN3_bit => VN_data_out(4437),
        VN2CN4_bit => VN_data_out(4438),
        VN2CN5_bit => VN_data_out(4439),
        VN2CN0_sign => VN_sign_out(4434),
        VN2CN1_sign => VN_sign_out(4435),
        VN2CN2_sign => VN_sign_out(4436),
        VN2CN3_sign => VN_sign_out(4437),
        VN2CN4_sign => VN_sign_out(4438),
        VN2CN5_sign => VN_sign_out(4439),
        codeword => codeword(739),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN740 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4445 downto 4440),
        Din0 => VN740_in0,
        Din1 => VN740_in1,
        Din2 => VN740_in2,
        Din3 => VN740_in3,
        Din4 => VN740_in4,
        Din5 => VN740_in5,
        VN2CN0_bit => VN_data_out(4440),
        VN2CN1_bit => VN_data_out(4441),
        VN2CN2_bit => VN_data_out(4442),
        VN2CN3_bit => VN_data_out(4443),
        VN2CN4_bit => VN_data_out(4444),
        VN2CN5_bit => VN_data_out(4445),
        VN2CN0_sign => VN_sign_out(4440),
        VN2CN1_sign => VN_sign_out(4441),
        VN2CN2_sign => VN_sign_out(4442),
        VN2CN3_sign => VN_sign_out(4443),
        VN2CN4_sign => VN_sign_out(4444),
        VN2CN5_sign => VN_sign_out(4445),
        codeword => codeword(740),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN741 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4451 downto 4446),
        Din0 => VN741_in0,
        Din1 => VN741_in1,
        Din2 => VN741_in2,
        Din3 => VN741_in3,
        Din4 => VN741_in4,
        Din5 => VN741_in5,
        VN2CN0_bit => VN_data_out(4446),
        VN2CN1_bit => VN_data_out(4447),
        VN2CN2_bit => VN_data_out(4448),
        VN2CN3_bit => VN_data_out(4449),
        VN2CN4_bit => VN_data_out(4450),
        VN2CN5_bit => VN_data_out(4451),
        VN2CN0_sign => VN_sign_out(4446),
        VN2CN1_sign => VN_sign_out(4447),
        VN2CN2_sign => VN_sign_out(4448),
        VN2CN3_sign => VN_sign_out(4449),
        VN2CN4_sign => VN_sign_out(4450),
        VN2CN5_sign => VN_sign_out(4451),
        codeword => codeword(741),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN742 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4457 downto 4452),
        Din0 => VN742_in0,
        Din1 => VN742_in1,
        Din2 => VN742_in2,
        Din3 => VN742_in3,
        Din4 => VN742_in4,
        Din5 => VN742_in5,
        VN2CN0_bit => VN_data_out(4452),
        VN2CN1_bit => VN_data_out(4453),
        VN2CN2_bit => VN_data_out(4454),
        VN2CN3_bit => VN_data_out(4455),
        VN2CN4_bit => VN_data_out(4456),
        VN2CN5_bit => VN_data_out(4457),
        VN2CN0_sign => VN_sign_out(4452),
        VN2CN1_sign => VN_sign_out(4453),
        VN2CN2_sign => VN_sign_out(4454),
        VN2CN3_sign => VN_sign_out(4455),
        VN2CN4_sign => VN_sign_out(4456),
        VN2CN5_sign => VN_sign_out(4457),
        codeword => codeword(742),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN743 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4463 downto 4458),
        Din0 => VN743_in0,
        Din1 => VN743_in1,
        Din2 => VN743_in2,
        Din3 => VN743_in3,
        Din4 => VN743_in4,
        Din5 => VN743_in5,
        VN2CN0_bit => VN_data_out(4458),
        VN2CN1_bit => VN_data_out(4459),
        VN2CN2_bit => VN_data_out(4460),
        VN2CN3_bit => VN_data_out(4461),
        VN2CN4_bit => VN_data_out(4462),
        VN2CN5_bit => VN_data_out(4463),
        VN2CN0_sign => VN_sign_out(4458),
        VN2CN1_sign => VN_sign_out(4459),
        VN2CN2_sign => VN_sign_out(4460),
        VN2CN3_sign => VN_sign_out(4461),
        VN2CN4_sign => VN_sign_out(4462),
        VN2CN5_sign => VN_sign_out(4463),
        codeword => codeword(743),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN744 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4469 downto 4464),
        Din0 => VN744_in0,
        Din1 => VN744_in1,
        Din2 => VN744_in2,
        Din3 => VN744_in3,
        Din4 => VN744_in4,
        Din5 => VN744_in5,
        VN2CN0_bit => VN_data_out(4464),
        VN2CN1_bit => VN_data_out(4465),
        VN2CN2_bit => VN_data_out(4466),
        VN2CN3_bit => VN_data_out(4467),
        VN2CN4_bit => VN_data_out(4468),
        VN2CN5_bit => VN_data_out(4469),
        VN2CN0_sign => VN_sign_out(4464),
        VN2CN1_sign => VN_sign_out(4465),
        VN2CN2_sign => VN_sign_out(4466),
        VN2CN3_sign => VN_sign_out(4467),
        VN2CN4_sign => VN_sign_out(4468),
        VN2CN5_sign => VN_sign_out(4469),
        codeword => codeword(744),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN745 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4475 downto 4470),
        Din0 => VN745_in0,
        Din1 => VN745_in1,
        Din2 => VN745_in2,
        Din3 => VN745_in3,
        Din4 => VN745_in4,
        Din5 => VN745_in5,
        VN2CN0_bit => VN_data_out(4470),
        VN2CN1_bit => VN_data_out(4471),
        VN2CN2_bit => VN_data_out(4472),
        VN2CN3_bit => VN_data_out(4473),
        VN2CN4_bit => VN_data_out(4474),
        VN2CN5_bit => VN_data_out(4475),
        VN2CN0_sign => VN_sign_out(4470),
        VN2CN1_sign => VN_sign_out(4471),
        VN2CN2_sign => VN_sign_out(4472),
        VN2CN3_sign => VN_sign_out(4473),
        VN2CN4_sign => VN_sign_out(4474),
        VN2CN5_sign => VN_sign_out(4475),
        codeword => codeword(745),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN746 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4481 downto 4476),
        Din0 => VN746_in0,
        Din1 => VN746_in1,
        Din2 => VN746_in2,
        Din3 => VN746_in3,
        Din4 => VN746_in4,
        Din5 => VN746_in5,
        VN2CN0_bit => VN_data_out(4476),
        VN2CN1_bit => VN_data_out(4477),
        VN2CN2_bit => VN_data_out(4478),
        VN2CN3_bit => VN_data_out(4479),
        VN2CN4_bit => VN_data_out(4480),
        VN2CN5_bit => VN_data_out(4481),
        VN2CN0_sign => VN_sign_out(4476),
        VN2CN1_sign => VN_sign_out(4477),
        VN2CN2_sign => VN_sign_out(4478),
        VN2CN3_sign => VN_sign_out(4479),
        VN2CN4_sign => VN_sign_out(4480),
        VN2CN5_sign => VN_sign_out(4481),
        codeword => codeword(746),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN747 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4487 downto 4482),
        Din0 => VN747_in0,
        Din1 => VN747_in1,
        Din2 => VN747_in2,
        Din3 => VN747_in3,
        Din4 => VN747_in4,
        Din5 => VN747_in5,
        VN2CN0_bit => VN_data_out(4482),
        VN2CN1_bit => VN_data_out(4483),
        VN2CN2_bit => VN_data_out(4484),
        VN2CN3_bit => VN_data_out(4485),
        VN2CN4_bit => VN_data_out(4486),
        VN2CN5_bit => VN_data_out(4487),
        VN2CN0_sign => VN_sign_out(4482),
        VN2CN1_sign => VN_sign_out(4483),
        VN2CN2_sign => VN_sign_out(4484),
        VN2CN3_sign => VN_sign_out(4485),
        VN2CN4_sign => VN_sign_out(4486),
        VN2CN5_sign => VN_sign_out(4487),
        codeword => codeword(747),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN748 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4493 downto 4488),
        Din0 => VN748_in0,
        Din1 => VN748_in1,
        Din2 => VN748_in2,
        Din3 => VN748_in3,
        Din4 => VN748_in4,
        Din5 => VN748_in5,
        VN2CN0_bit => VN_data_out(4488),
        VN2CN1_bit => VN_data_out(4489),
        VN2CN2_bit => VN_data_out(4490),
        VN2CN3_bit => VN_data_out(4491),
        VN2CN4_bit => VN_data_out(4492),
        VN2CN5_bit => VN_data_out(4493),
        VN2CN0_sign => VN_sign_out(4488),
        VN2CN1_sign => VN_sign_out(4489),
        VN2CN2_sign => VN_sign_out(4490),
        VN2CN3_sign => VN_sign_out(4491),
        VN2CN4_sign => VN_sign_out(4492),
        VN2CN5_sign => VN_sign_out(4493),
        codeword => codeword(748),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN749 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4499 downto 4494),
        Din0 => VN749_in0,
        Din1 => VN749_in1,
        Din2 => VN749_in2,
        Din3 => VN749_in3,
        Din4 => VN749_in4,
        Din5 => VN749_in5,
        VN2CN0_bit => VN_data_out(4494),
        VN2CN1_bit => VN_data_out(4495),
        VN2CN2_bit => VN_data_out(4496),
        VN2CN3_bit => VN_data_out(4497),
        VN2CN4_bit => VN_data_out(4498),
        VN2CN5_bit => VN_data_out(4499),
        VN2CN0_sign => VN_sign_out(4494),
        VN2CN1_sign => VN_sign_out(4495),
        VN2CN2_sign => VN_sign_out(4496),
        VN2CN3_sign => VN_sign_out(4497),
        VN2CN4_sign => VN_sign_out(4498),
        VN2CN5_sign => VN_sign_out(4499),
        codeword => codeword(749),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN750 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4505 downto 4500),
        Din0 => VN750_in0,
        Din1 => VN750_in1,
        Din2 => VN750_in2,
        Din3 => VN750_in3,
        Din4 => VN750_in4,
        Din5 => VN750_in5,
        VN2CN0_bit => VN_data_out(4500),
        VN2CN1_bit => VN_data_out(4501),
        VN2CN2_bit => VN_data_out(4502),
        VN2CN3_bit => VN_data_out(4503),
        VN2CN4_bit => VN_data_out(4504),
        VN2CN5_bit => VN_data_out(4505),
        VN2CN0_sign => VN_sign_out(4500),
        VN2CN1_sign => VN_sign_out(4501),
        VN2CN2_sign => VN_sign_out(4502),
        VN2CN3_sign => VN_sign_out(4503),
        VN2CN4_sign => VN_sign_out(4504),
        VN2CN5_sign => VN_sign_out(4505),
        codeword => codeword(750),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN751 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4511 downto 4506),
        Din0 => VN751_in0,
        Din1 => VN751_in1,
        Din2 => VN751_in2,
        Din3 => VN751_in3,
        Din4 => VN751_in4,
        Din5 => VN751_in5,
        VN2CN0_bit => VN_data_out(4506),
        VN2CN1_bit => VN_data_out(4507),
        VN2CN2_bit => VN_data_out(4508),
        VN2CN3_bit => VN_data_out(4509),
        VN2CN4_bit => VN_data_out(4510),
        VN2CN5_bit => VN_data_out(4511),
        VN2CN0_sign => VN_sign_out(4506),
        VN2CN1_sign => VN_sign_out(4507),
        VN2CN2_sign => VN_sign_out(4508),
        VN2CN3_sign => VN_sign_out(4509),
        VN2CN4_sign => VN_sign_out(4510),
        VN2CN5_sign => VN_sign_out(4511),
        codeword => codeword(751),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN752 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4517 downto 4512),
        Din0 => VN752_in0,
        Din1 => VN752_in1,
        Din2 => VN752_in2,
        Din3 => VN752_in3,
        Din4 => VN752_in4,
        Din5 => VN752_in5,
        VN2CN0_bit => VN_data_out(4512),
        VN2CN1_bit => VN_data_out(4513),
        VN2CN2_bit => VN_data_out(4514),
        VN2CN3_bit => VN_data_out(4515),
        VN2CN4_bit => VN_data_out(4516),
        VN2CN5_bit => VN_data_out(4517),
        VN2CN0_sign => VN_sign_out(4512),
        VN2CN1_sign => VN_sign_out(4513),
        VN2CN2_sign => VN_sign_out(4514),
        VN2CN3_sign => VN_sign_out(4515),
        VN2CN4_sign => VN_sign_out(4516),
        VN2CN5_sign => VN_sign_out(4517),
        codeword => codeword(752),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN753 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4523 downto 4518),
        Din0 => VN753_in0,
        Din1 => VN753_in1,
        Din2 => VN753_in2,
        Din3 => VN753_in3,
        Din4 => VN753_in4,
        Din5 => VN753_in5,
        VN2CN0_bit => VN_data_out(4518),
        VN2CN1_bit => VN_data_out(4519),
        VN2CN2_bit => VN_data_out(4520),
        VN2CN3_bit => VN_data_out(4521),
        VN2CN4_bit => VN_data_out(4522),
        VN2CN5_bit => VN_data_out(4523),
        VN2CN0_sign => VN_sign_out(4518),
        VN2CN1_sign => VN_sign_out(4519),
        VN2CN2_sign => VN_sign_out(4520),
        VN2CN3_sign => VN_sign_out(4521),
        VN2CN4_sign => VN_sign_out(4522),
        VN2CN5_sign => VN_sign_out(4523),
        codeword => codeword(753),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN754 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4529 downto 4524),
        Din0 => VN754_in0,
        Din1 => VN754_in1,
        Din2 => VN754_in2,
        Din3 => VN754_in3,
        Din4 => VN754_in4,
        Din5 => VN754_in5,
        VN2CN0_bit => VN_data_out(4524),
        VN2CN1_bit => VN_data_out(4525),
        VN2CN2_bit => VN_data_out(4526),
        VN2CN3_bit => VN_data_out(4527),
        VN2CN4_bit => VN_data_out(4528),
        VN2CN5_bit => VN_data_out(4529),
        VN2CN0_sign => VN_sign_out(4524),
        VN2CN1_sign => VN_sign_out(4525),
        VN2CN2_sign => VN_sign_out(4526),
        VN2CN3_sign => VN_sign_out(4527),
        VN2CN4_sign => VN_sign_out(4528),
        VN2CN5_sign => VN_sign_out(4529),
        codeword => codeword(754),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN755 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4535 downto 4530),
        Din0 => VN755_in0,
        Din1 => VN755_in1,
        Din2 => VN755_in2,
        Din3 => VN755_in3,
        Din4 => VN755_in4,
        Din5 => VN755_in5,
        VN2CN0_bit => VN_data_out(4530),
        VN2CN1_bit => VN_data_out(4531),
        VN2CN2_bit => VN_data_out(4532),
        VN2CN3_bit => VN_data_out(4533),
        VN2CN4_bit => VN_data_out(4534),
        VN2CN5_bit => VN_data_out(4535),
        VN2CN0_sign => VN_sign_out(4530),
        VN2CN1_sign => VN_sign_out(4531),
        VN2CN2_sign => VN_sign_out(4532),
        VN2CN3_sign => VN_sign_out(4533),
        VN2CN4_sign => VN_sign_out(4534),
        VN2CN5_sign => VN_sign_out(4535),
        codeword => codeword(755),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN756 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4541 downto 4536),
        Din0 => VN756_in0,
        Din1 => VN756_in1,
        Din2 => VN756_in2,
        Din3 => VN756_in3,
        Din4 => VN756_in4,
        Din5 => VN756_in5,
        VN2CN0_bit => VN_data_out(4536),
        VN2CN1_bit => VN_data_out(4537),
        VN2CN2_bit => VN_data_out(4538),
        VN2CN3_bit => VN_data_out(4539),
        VN2CN4_bit => VN_data_out(4540),
        VN2CN5_bit => VN_data_out(4541),
        VN2CN0_sign => VN_sign_out(4536),
        VN2CN1_sign => VN_sign_out(4537),
        VN2CN2_sign => VN_sign_out(4538),
        VN2CN3_sign => VN_sign_out(4539),
        VN2CN4_sign => VN_sign_out(4540),
        VN2CN5_sign => VN_sign_out(4541),
        codeword => codeword(756),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN757 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4547 downto 4542),
        Din0 => VN757_in0,
        Din1 => VN757_in1,
        Din2 => VN757_in2,
        Din3 => VN757_in3,
        Din4 => VN757_in4,
        Din5 => VN757_in5,
        VN2CN0_bit => VN_data_out(4542),
        VN2CN1_bit => VN_data_out(4543),
        VN2CN2_bit => VN_data_out(4544),
        VN2CN3_bit => VN_data_out(4545),
        VN2CN4_bit => VN_data_out(4546),
        VN2CN5_bit => VN_data_out(4547),
        VN2CN0_sign => VN_sign_out(4542),
        VN2CN1_sign => VN_sign_out(4543),
        VN2CN2_sign => VN_sign_out(4544),
        VN2CN3_sign => VN_sign_out(4545),
        VN2CN4_sign => VN_sign_out(4546),
        VN2CN5_sign => VN_sign_out(4547),
        codeword => codeword(757),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN758 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4553 downto 4548),
        Din0 => VN758_in0,
        Din1 => VN758_in1,
        Din2 => VN758_in2,
        Din3 => VN758_in3,
        Din4 => VN758_in4,
        Din5 => VN758_in5,
        VN2CN0_bit => VN_data_out(4548),
        VN2CN1_bit => VN_data_out(4549),
        VN2CN2_bit => VN_data_out(4550),
        VN2CN3_bit => VN_data_out(4551),
        VN2CN4_bit => VN_data_out(4552),
        VN2CN5_bit => VN_data_out(4553),
        VN2CN0_sign => VN_sign_out(4548),
        VN2CN1_sign => VN_sign_out(4549),
        VN2CN2_sign => VN_sign_out(4550),
        VN2CN3_sign => VN_sign_out(4551),
        VN2CN4_sign => VN_sign_out(4552),
        VN2CN5_sign => VN_sign_out(4553),
        codeword => codeword(758),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN759 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4559 downto 4554),
        Din0 => VN759_in0,
        Din1 => VN759_in1,
        Din2 => VN759_in2,
        Din3 => VN759_in3,
        Din4 => VN759_in4,
        Din5 => VN759_in5,
        VN2CN0_bit => VN_data_out(4554),
        VN2CN1_bit => VN_data_out(4555),
        VN2CN2_bit => VN_data_out(4556),
        VN2CN3_bit => VN_data_out(4557),
        VN2CN4_bit => VN_data_out(4558),
        VN2CN5_bit => VN_data_out(4559),
        VN2CN0_sign => VN_sign_out(4554),
        VN2CN1_sign => VN_sign_out(4555),
        VN2CN2_sign => VN_sign_out(4556),
        VN2CN3_sign => VN_sign_out(4557),
        VN2CN4_sign => VN_sign_out(4558),
        VN2CN5_sign => VN_sign_out(4559),
        codeword => codeword(759),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN760 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4565 downto 4560),
        Din0 => VN760_in0,
        Din1 => VN760_in1,
        Din2 => VN760_in2,
        Din3 => VN760_in3,
        Din4 => VN760_in4,
        Din5 => VN760_in5,
        VN2CN0_bit => VN_data_out(4560),
        VN2CN1_bit => VN_data_out(4561),
        VN2CN2_bit => VN_data_out(4562),
        VN2CN3_bit => VN_data_out(4563),
        VN2CN4_bit => VN_data_out(4564),
        VN2CN5_bit => VN_data_out(4565),
        VN2CN0_sign => VN_sign_out(4560),
        VN2CN1_sign => VN_sign_out(4561),
        VN2CN2_sign => VN_sign_out(4562),
        VN2CN3_sign => VN_sign_out(4563),
        VN2CN4_sign => VN_sign_out(4564),
        VN2CN5_sign => VN_sign_out(4565),
        codeword => codeword(760),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN761 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4571 downto 4566),
        Din0 => VN761_in0,
        Din1 => VN761_in1,
        Din2 => VN761_in2,
        Din3 => VN761_in3,
        Din4 => VN761_in4,
        Din5 => VN761_in5,
        VN2CN0_bit => VN_data_out(4566),
        VN2CN1_bit => VN_data_out(4567),
        VN2CN2_bit => VN_data_out(4568),
        VN2CN3_bit => VN_data_out(4569),
        VN2CN4_bit => VN_data_out(4570),
        VN2CN5_bit => VN_data_out(4571),
        VN2CN0_sign => VN_sign_out(4566),
        VN2CN1_sign => VN_sign_out(4567),
        VN2CN2_sign => VN_sign_out(4568),
        VN2CN3_sign => VN_sign_out(4569),
        VN2CN4_sign => VN_sign_out(4570),
        VN2CN5_sign => VN_sign_out(4571),
        codeword => codeword(761),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN762 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4577 downto 4572),
        Din0 => VN762_in0,
        Din1 => VN762_in1,
        Din2 => VN762_in2,
        Din3 => VN762_in3,
        Din4 => VN762_in4,
        Din5 => VN762_in5,
        VN2CN0_bit => VN_data_out(4572),
        VN2CN1_bit => VN_data_out(4573),
        VN2CN2_bit => VN_data_out(4574),
        VN2CN3_bit => VN_data_out(4575),
        VN2CN4_bit => VN_data_out(4576),
        VN2CN5_bit => VN_data_out(4577),
        VN2CN0_sign => VN_sign_out(4572),
        VN2CN1_sign => VN_sign_out(4573),
        VN2CN2_sign => VN_sign_out(4574),
        VN2CN3_sign => VN_sign_out(4575),
        VN2CN4_sign => VN_sign_out(4576),
        VN2CN5_sign => VN_sign_out(4577),
        codeword => codeword(762),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN763 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4583 downto 4578),
        Din0 => VN763_in0,
        Din1 => VN763_in1,
        Din2 => VN763_in2,
        Din3 => VN763_in3,
        Din4 => VN763_in4,
        Din5 => VN763_in5,
        VN2CN0_bit => VN_data_out(4578),
        VN2CN1_bit => VN_data_out(4579),
        VN2CN2_bit => VN_data_out(4580),
        VN2CN3_bit => VN_data_out(4581),
        VN2CN4_bit => VN_data_out(4582),
        VN2CN5_bit => VN_data_out(4583),
        VN2CN0_sign => VN_sign_out(4578),
        VN2CN1_sign => VN_sign_out(4579),
        VN2CN2_sign => VN_sign_out(4580),
        VN2CN3_sign => VN_sign_out(4581),
        VN2CN4_sign => VN_sign_out(4582),
        VN2CN5_sign => VN_sign_out(4583),
        codeword => codeword(763),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN764 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4589 downto 4584),
        Din0 => VN764_in0,
        Din1 => VN764_in1,
        Din2 => VN764_in2,
        Din3 => VN764_in3,
        Din4 => VN764_in4,
        Din5 => VN764_in5,
        VN2CN0_bit => VN_data_out(4584),
        VN2CN1_bit => VN_data_out(4585),
        VN2CN2_bit => VN_data_out(4586),
        VN2CN3_bit => VN_data_out(4587),
        VN2CN4_bit => VN_data_out(4588),
        VN2CN5_bit => VN_data_out(4589),
        VN2CN0_sign => VN_sign_out(4584),
        VN2CN1_sign => VN_sign_out(4585),
        VN2CN2_sign => VN_sign_out(4586),
        VN2CN3_sign => VN_sign_out(4587),
        VN2CN4_sign => VN_sign_out(4588),
        VN2CN5_sign => VN_sign_out(4589),
        codeword => codeword(764),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN765 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4595 downto 4590),
        Din0 => VN765_in0,
        Din1 => VN765_in1,
        Din2 => VN765_in2,
        Din3 => VN765_in3,
        Din4 => VN765_in4,
        Din5 => VN765_in5,
        VN2CN0_bit => VN_data_out(4590),
        VN2CN1_bit => VN_data_out(4591),
        VN2CN2_bit => VN_data_out(4592),
        VN2CN3_bit => VN_data_out(4593),
        VN2CN4_bit => VN_data_out(4594),
        VN2CN5_bit => VN_data_out(4595),
        VN2CN0_sign => VN_sign_out(4590),
        VN2CN1_sign => VN_sign_out(4591),
        VN2CN2_sign => VN_sign_out(4592),
        VN2CN3_sign => VN_sign_out(4593),
        VN2CN4_sign => VN_sign_out(4594),
        VN2CN5_sign => VN_sign_out(4595),
        codeword => codeword(765),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN766 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4601 downto 4596),
        Din0 => VN766_in0,
        Din1 => VN766_in1,
        Din2 => VN766_in2,
        Din3 => VN766_in3,
        Din4 => VN766_in4,
        Din5 => VN766_in5,
        VN2CN0_bit => VN_data_out(4596),
        VN2CN1_bit => VN_data_out(4597),
        VN2CN2_bit => VN_data_out(4598),
        VN2CN3_bit => VN_data_out(4599),
        VN2CN4_bit => VN_data_out(4600),
        VN2CN5_bit => VN_data_out(4601),
        VN2CN0_sign => VN_sign_out(4596),
        VN2CN1_sign => VN_sign_out(4597),
        VN2CN2_sign => VN_sign_out(4598),
        VN2CN3_sign => VN_sign_out(4599),
        VN2CN4_sign => VN_sign_out(4600),
        VN2CN5_sign => VN_sign_out(4601),
        codeword => codeword(766),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN767 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4607 downto 4602),
        Din0 => VN767_in0,
        Din1 => VN767_in1,
        Din2 => VN767_in2,
        Din3 => VN767_in3,
        Din4 => VN767_in4,
        Din5 => VN767_in5,
        VN2CN0_bit => VN_data_out(4602),
        VN2CN1_bit => VN_data_out(4603),
        VN2CN2_bit => VN_data_out(4604),
        VN2CN3_bit => VN_data_out(4605),
        VN2CN4_bit => VN_data_out(4606),
        VN2CN5_bit => VN_data_out(4607),
        VN2CN0_sign => VN_sign_out(4602),
        VN2CN1_sign => VN_sign_out(4603),
        VN2CN2_sign => VN_sign_out(4604),
        VN2CN3_sign => VN_sign_out(4605),
        VN2CN4_sign => VN_sign_out(4606),
        VN2CN5_sign => VN_sign_out(4607),
        codeword => codeword(767),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN768 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4613 downto 4608),
        Din0 => VN768_in0,
        Din1 => VN768_in1,
        Din2 => VN768_in2,
        Din3 => VN768_in3,
        Din4 => VN768_in4,
        Din5 => VN768_in5,
        VN2CN0_bit => VN_data_out(4608),
        VN2CN1_bit => VN_data_out(4609),
        VN2CN2_bit => VN_data_out(4610),
        VN2CN3_bit => VN_data_out(4611),
        VN2CN4_bit => VN_data_out(4612),
        VN2CN5_bit => VN_data_out(4613),
        VN2CN0_sign => VN_sign_out(4608),
        VN2CN1_sign => VN_sign_out(4609),
        VN2CN2_sign => VN_sign_out(4610),
        VN2CN3_sign => VN_sign_out(4611),
        VN2CN4_sign => VN_sign_out(4612),
        VN2CN5_sign => VN_sign_out(4613),
        codeword => codeword(768),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN769 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4619 downto 4614),
        Din0 => VN769_in0,
        Din1 => VN769_in1,
        Din2 => VN769_in2,
        Din3 => VN769_in3,
        Din4 => VN769_in4,
        Din5 => VN769_in5,
        VN2CN0_bit => VN_data_out(4614),
        VN2CN1_bit => VN_data_out(4615),
        VN2CN2_bit => VN_data_out(4616),
        VN2CN3_bit => VN_data_out(4617),
        VN2CN4_bit => VN_data_out(4618),
        VN2CN5_bit => VN_data_out(4619),
        VN2CN0_sign => VN_sign_out(4614),
        VN2CN1_sign => VN_sign_out(4615),
        VN2CN2_sign => VN_sign_out(4616),
        VN2CN3_sign => VN_sign_out(4617),
        VN2CN4_sign => VN_sign_out(4618),
        VN2CN5_sign => VN_sign_out(4619),
        codeword => codeword(769),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN770 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4625 downto 4620),
        Din0 => VN770_in0,
        Din1 => VN770_in1,
        Din2 => VN770_in2,
        Din3 => VN770_in3,
        Din4 => VN770_in4,
        Din5 => VN770_in5,
        VN2CN0_bit => VN_data_out(4620),
        VN2CN1_bit => VN_data_out(4621),
        VN2CN2_bit => VN_data_out(4622),
        VN2CN3_bit => VN_data_out(4623),
        VN2CN4_bit => VN_data_out(4624),
        VN2CN5_bit => VN_data_out(4625),
        VN2CN0_sign => VN_sign_out(4620),
        VN2CN1_sign => VN_sign_out(4621),
        VN2CN2_sign => VN_sign_out(4622),
        VN2CN3_sign => VN_sign_out(4623),
        VN2CN4_sign => VN_sign_out(4624),
        VN2CN5_sign => VN_sign_out(4625),
        codeword => codeword(770),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN771 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4631 downto 4626),
        Din0 => VN771_in0,
        Din1 => VN771_in1,
        Din2 => VN771_in2,
        Din3 => VN771_in3,
        Din4 => VN771_in4,
        Din5 => VN771_in5,
        VN2CN0_bit => VN_data_out(4626),
        VN2CN1_bit => VN_data_out(4627),
        VN2CN2_bit => VN_data_out(4628),
        VN2CN3_bit => VN_data_out(4629),
        VN2CN4_bit => VN_data_out(4630),
        VN2CN5_bit => VN_data_out(4631),
        VN2CN0_sign => VN_sign_out(4626),
        VN2CN1_sign => VN_sign_out(4627),
        VN2CN2_sign => VN_sign_out(4628),
        VN2CN3_sign => VN_sign_out(4629),
        VN2CN4_sign => VN_sign_out(4630),
        VN2CN5_sign => VN_sign_out(4631),
        codeword => codeword(771),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN772 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4637 downto 4632),
        Din0 => VN772_in0,
        Din1 => VN772_in1,
        Din2 => VN772_in2,
        Din3 => VN772_in3,
        Din4 => VN772_in4,
        Din5 => VN772_in5,
        VN2CN0_bit => VN_data_out(4632),
        VN2CN1_bit => VN_data_out(4633),
        VN2CN2_bit => VN_data_out(4634),
        VN2CN3_bit => VN_data_out(4635),
        VN2CN4_bit => VN_data_out(4636),
        VN2CN5_bit => VN_data_out(4637),
        VN2CN0_sign => VN_sign_out(4632),
        VN2CN1_sign => VN_sign_out(4633),
        VN2CN2_sign => VN_sign_out(4634),
        VN2CN3_sign => VN_sign_out(4635),
        VN2CN4_sign => VN_sign_out(4636),
        VN2CN5_sign => VN_sign_out(4637),
        codeword => codeword(772),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN773 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4643 downto 4638),
        Din0 => VN773_in0,
        Din1 => VN773_in1,
        Din2 => VN773_in2,
        Din3 => VN773_in3,
        Din4 => VN773_in4,
        Din5 => VN773_in5,
        VN2CN0_bit => VN_data_out(4638),
        VN2CN1_bit => VN_data_out(4639),
        VN2CN2_bit => VN_data_out(4640),
        VN2CN3_bit => VN_data_out(4641),
        VN2CN4_bit => VN_data_out(4642),
        VN2CN5_bit => VN_data_out(4643),
        VN2CN0_sign => VN_sign_out(4638),
        VN2CN1_sign => VN_sign_out(4639),
        VN2CN2_sign => VN_sign_out(4640),
        VN2CN3_sign => VN_sign_out(4641),
        VN2CN4_sign => VN_sign_out(4642),
        VN2CN5_sign => VN_sign_out(4643),
        codeword => codeword(773),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN774 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4649 downto 4644),
        Din0 => VN774_in0,
        Din1 => VN774_in1,
        Din2 => VN774_in2,
        Din3 => VN774_in3,
        Din4 => VN774_in4,
        Din5 => VN774_in5,
        VN2CN0_bit => VN_data_out(4644),
        VN2CN1_bit => VN_data_out(4645),
        VN2CN2_bit => VN_data_out(4646),
        VN2CN3_bit => VN_data_out(4647),
        VN2CN4_bit => VN_data_out(4648),
        VN2CN5_bit => VN_data_out(4649),
        VN2CN0_sign => VN_sign_out(4644),
        VN2CN1_sign => VN_sign_out(4645),
        VN2CN2_sign => VN_sign_out(4646),
        VN2CN3_sign => VN_sign_out(4647),
        VN2CN4_sign => VN_sign_out(4648),
        VN2CN5_sign => VN_sign_out(4649),
        codeword => codeword(774),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN775 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4655 downto 4650),
        Din0 => VN775_in0,
        Din1 => VN775_in1,
        Din2 => VN775_in2,
        Din3 => VN775_in3,
        Din4 => VN775_in4,
        Din5 => VN775_in5,
        VN2CN0_bit => VN_data_out(4650),
        VN2CN1_bit => VN_data_out(4651),
        VN2CN2_bit => VN_data_out(4652),
        VN2CN3_bit => VN_data_out(4653),
        VN2CN4_bit => VN_data_out(4654),
        VN2CN5_bit => VN_data_out(4655),
        VN2CN0_sign => VN_sign_out(4650),
        VN2CN1_sign => VN_sign_out(4651),
        VN2CN2_sign => VN_sign_out(4652),
        VN2CN3_sign => VN_sign_out(4653),
        VN2CN4_sign => VN_sign_out(4654),
        VN2CN5_sign => VN_sign_out(4655),
        codeword => codeword(775),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN776 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4661 downto 4656),
        Din0 => VN776_in0,
        Din1 => VN776_in1,
        Din2 => VN776_in2,
        Din3 => VN776_in3,
        Din4 => VN776_in4,
        Din5 => VN776_in5,
        VN2CN0_bit => VN_data_out(4656),
        VN2CN1_bit => VN_data_out(4657),
        VN2CN2_bit => VN_data_out(4658),
        VN2CN3_bit => VN_data_out(4659),
        VN2CN4_bit => VN_data_out(4660),
        VN2CN5_bit => VN_data_out(4661),
        VN2CN0_sign => VN_sign_out(4656),
        VN2CN1_sign => VN_sign_out(4657),
        VN2CN2_sign => VN_sign_out(4658),
        VN2CN3_sign => VN_sign_out(4659),
        VN2CN4_sign => VN_sign_out(4660),
        VN2CN5_sign => VN_sign_out(4661),
        codeword => codeword(776),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN777 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4667 downto 4662),
        Din0 => VN777_in0,
        Din1 => VN777_in1,
        Din2 => VN777_in2,
        Din3 => VN777_in3,
        Din4 => VN777_in4,
        Din5 => VN777_in5,
        VN2CN0_bit => VN_data_out(4662),
        VN2CN1_bit => VN_data_out(4663),
        VN2CN2_bit => VN_data_out(4664),
        VN2CN3_bit => VN_data_out(4665),
        VN2CN4_bit => VN_data_out(4666),
        VN2CN5_bit => VN_data_out(4667),
        VN2CN0_sign => VN_sign_out(4662),
        VN2CN1_sign => VN_sign_out(4663),
        VN2CN2_sign => VN_sign_out(4664),
        VN2CN3_sign => VN_sign_out(4665),
        VN2CN4_sign => VN_sign_out(4666),
        VN2CN5_sign => VN_sign_out(4667),
        codeword => codeword(777),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN778 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4673 downto 4668),
        Din0 => VN778_in0,
        Din1 => VN778_in1,
        Din2 => VN778_in2,
        Din3 => VN778_in3,
        Din4 => VN778_in4,
        Din5 => VN778_in5,
        VN2CN0_bit => VN_data_out(4668),
        VN2CN1_bit => VN_data_out(4669),
        VN2CN2_bit => VN_data_out(4670),
        VN2CN3_bit => VN_data_out(4671),
        VN2CN4_bit => VN_data_out(4672),
        VN2CN5_bit => VN_data_out(4673),
        VN2CN0_sign => VN_sign_out(4668),
        VN2CN1_sign => VN_sign_out(4669),
        VN2CN2_sign => VN_sign_out(4670),
        VN2CN3_sign => VN_sign_out(4671),
        VN2CN4_sign => VN_sign_out(4672),
        VN2CN5_sign => VN_sign_out(4673),
        codeword => codeword(778),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN779 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4679 downto 4674),
        Din0 => VN779_in0,
        Din1 => VN779_in1,
        Din2 => VN779_in2,
        Din3 => VN779_in3,
        Din4 => VN779_in4,
        Din5 => VN779_in5,
        VN2CN0_bit => VN_data_out(4674),
        VN2CN1_bit => VN_data_out(4675),
        VN2CN2_bit => VN_data_out(4676),
        VN2CN3_bit => VN_data_out(4677),
        VN2CN4_bit => VN_data_out(4678),
        VN2CN5_bit => VN_data_out(4679),
        VN2CN0_sign => VN_sign_out(4674),
        VN2CN1_sign => VN_sign_out(4675),
        VN2CN2_sign => VN_sign_out(4676),
        VN2CN3_sign => VN_sign_out(4677),
        VN2CN4_sign => VN_sign_out(4678),
        VN2CN5_sign => VN_sign_out(4679),
        codeword => codeword(779),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN780 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4685 downto 4680),
        Din0 => VN780_in0,
        Din1 => VN780_in1,
        Din2 => VN780_in2,
        Din3 => VN780_in3,
        Din4 => VN780_in4,
        Din5 => VN780_in5,
        VN2CN0_bit => VN_data_out(4680),
        VN2CN1_bit => VN_data_out(4681),
        VN2CN2_bit => VN_data_out(4682),
        VN2CN3_bit => VN_data_out(4683),
        VN2CN4_bit => VN_data_out(4684),
        VN2CN5_bit => VN_data_out(4685),
        VN2CN0_sign => VN_sign_out(4680),
        VN2CN1_sign => VN_sign_out(4681),
        VN2CN2_sign => VN_sign_out(4682),
        VN2CN3_sign => VN_sign_out(4683),
        VN2CN4_sign => VN_sign_out(4684),
        VN2CN5_sign => VN_sign_out(4685),
        codeword => codeword(780),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN781 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4691 downto 4686),
        Din0 => VN781_in0,
        Din1 => VN781_in1,
        Din2 => VN781_in2,
        Din3 => VN781_in3,
        Din4 => VN781_in4,
        Din5 => VN781_in5,
        VN2CN0_bit => VN_data_out(4686),
        VN2CN1_bit => VN_data_out(4687),
        VN2CN2_bit => VN_data_out(4688),
        VN2CN3_bit => VN_data_out(4689),
        VN2CN4_bit => VN_data_out(4690),
        VN2CN5_bit => VN_data_out(4691),
        VN2CN0_sign => VN_sign_out(4686),
        VN2CN1_sign => VN_sign_out(4687),
        VN2CN2_sign => VN_sign_out(4688),
        VN2CN3_sign => VN_sign_out(4689),
        VN2CN4_sign => VN_sign_out(4690),
        VN2CN5_sign => VN_sign_out(4691),
        codeword => codeword(781),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN782 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4697 downto 4692),
        Din0 => VN782_in0,
        Din1 => VN782_in1,
        Din2 => VN782_in2,
        Din3 => VN782_in3,
        Din4 => VN782_in4,
        Din5 => VN782_in5,
        VN2CN0_bit => VN_data_out(4692),
        VN2CN1_bit => VN_data_out(4693),
        VN2CN2_bit => VN_data_out(4694),
        VN2CN3_bit => VN_data_out(4695),
        VN2CN4_bit => VN_data_out(4696),
        VN2CN5_bit => VN_data_out(4697),
        VN2CN0_sign => VN_sign_out(4692),
        VN2CN1_sign => VN_sign_out(4693),
        VN2CN2_sign => VN_sign_out(4694),
        VN2CN3_sign => VN_sign_out(4695),
        VN2CN4_sign => VN_sign_out(4696),
        VN2CN5_sign => VN_sign_out(4697),
        codeword => codeword(782),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN783 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4703 downto 4698),
        Din0 => VN783_in0,
        Din1 => VN783_in1,
        Din2 => VN783_in2,
        Din3 => VN783_in3,
        Din4 => VN783_in4,
        Din5 => VN783_in5,
        VN2CN0_bit => VN_data_out(4698),
        VN2CN1_bit => VN_data_out(4699),
        VN2CN2_bit => VN_data_out(4700),
        VN2CN3_bit => VN_data_out(4701),
        VN2CN4_bit => VN_data_out(4702),
        VN2CN5_bit => VN_data_out(4703),
        VN2CN0_sign => VN_sign_out(4698),
        VN2CN1_sign => VN_sign_out(4699),
        VN2CN2_sign => VN_sign_out(4700),
        VN2CN3_sign => VN_sign_out(4701),
        VN2CN4_sign => VN_sign_out(4702),
        VN2CN5_sign => VN_sign_out(4703),
        codeword => codeword(783),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN784 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4709 downto 4704),
        Din0 => VN784_in0,
        Din1 => VN784_in1,
        Din2 => VN784_in2,
        Din3 => VN784_in3,
        Din4 => VN784_in4,
        Din5 => VN784_in5,
        VN2CN0_bit => VN_data_out(4704),
        VN2CN1_bit => VN_data_out(4705),
        VN2CN2_bit => VN_data_out(4706),
        VN2CN3_bit => VN_data_out(4707),
        VN2CN4_bit => VN_data_out(4708),
        VN2CN5_bit => VN_data_out(4709),
        VN2CN0_sign => VN_sign_out(4704),
        VN2CN1_sign => VN_sign_out(4705),
        VN2CN2_sign => VN_sign_out(4706),
        VN2CN3_sign => VN_sign_out(4707),
        VN2CN4_sign => VN_sign_out(4708),
        VN2CN5_sign => VN_sign_out(4709),
        codeword => codeword(784),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN785 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4715 downto 4710),
        Din0 => VN785_in0,
        Din1 => VN785_in1,
        Din2 => VN785_in2,
        Din3 => VN785_in3,
        Din4 => VN785_in4,
        Din5 => VN785_in5,
        VN2CN0_bit => VN_data_out(4710),
        VN2CN1_bit => VN_data_out(4711),
        VN2CN2_bit => VN_data_out(4712),
        VN2CN3_bit => VN_data_out(4713),
        VN2CN4_bit => VN_data_out(4714),
        VN2CN5_bit => VN_data_out(4715),
        VN2CN0_sign => VN_sign_out(4710),
        VN2CN1_sign => VN_sign_out(4711),
        VN2CN2_sign => VN_sign_out(4712),
        VN2CN3_sign => VN_sign_out(4713),
        VN2CN4_sign => VN_sign_out(4714),
        VN2CN5_sign => VN_sign_out(4715),
        codeword => codeword(785),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN786 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4721 downto 4716),
        Din0 => VN786_in0,
        Din1 => VN786_in1,
        Din2 => VN786_in2,
        Din3 => VN786_in3,
        Din4 => VN786_in4,
        Din5 => VN786_in5,
        VN2CN0_bit => VN_data_out(4716),
        VN2CN1_bit => VN_data_out(4717),
        VN2CN2_bit => VN_data_out(4718),
        VN2CN3_bit => VN_data_out(4719),
        VN2CN4_bit => VN_data_out(4720),
        VN2CN5_bit => VN_data_out(4721),
        VN2CN0_sign => VN_sign_out(4716),
        VN2CN1_sign => VN_sign_out(4717),
        VN2CN2_sign => VN_sign_out(4718),
        VN2CN3_sign => VN_sign_out(4719),
        VN2CN4_sign => VN_sign_out(4720),
        VN2CN5_sign => VN_sign_out(4721),
        codeword => codeword(786),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN787 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4727 downto 4722),
        Din0 => VN787_in0,
        Din1 => VN787_in1,
        Din2 => VN787_in2,
        Din3 => VN787_in3,
        Din4 => VN787_in4,
        Din5 => VN787_in5,
        VN2CN0_bit => VN_data_out(4722),
        VN2CN1_bit => VN_data_out(4723),
        VN2CN2_bit => VN_data_out(4724),
        VN2CN3_bit => VN_data_out(4725),
        VN2CN4_bit => VN_data_out(4726),
        VN2CN5_bit => VN_data_out(4727),
        VN2CN0_sign => VN_sign_out(4722),
        VN2CN1_sign => VN_sign_out(4723),
        VN2CN2_sign => VN_sign_out(4724),
        VN2CN3_sign => VN_sign_out(4725),
        VN2CN4_sign => VN_sign_out(4726),
        VN2CN5_sign => VN_sign_out(4727),
        codeword => codeword(787),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN788 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4733 downto 4728),
        Din0 => VN788_in0,
        Din1 => VN788_in1,
        Din2 => VN788_in2,
        Din3 => VN788_in3,
        Din4 => VN788_in4,
        Din5 => VN788_in5,
        VN2CN0_bit => VN_data_out(4728),
        VN2CN1_bit => VN_data_out(4729),
        VN2CN2_bit => VN_data_out(4730),
        VN2CN3_bit => VN_data_out(4731),
        VN2CN4_bit => VN_data_out(4732),
        VN2CN5_bit => VN_data_out(4733),
        VN2CN0_sign => VN_sign_out(4728),
        VN2CN1_sign => VN_sign_out(4729),
        VN2CN2_sign => VN_sign_out(4730),
        VN2CN3_sign => VN_sign_out(4731),
        VN2CN4_sign => VN_sign_out(4732),
        VN2CN5_sign => VN_sign_out(4733),
        codeword => codeword(788),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN789 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4739 downto 4734),
        Din0 => VN789_in0,
        Din1 => VN789_in1,
        Din2 => VN789_in2,
        Din3 => VN789_in3,
        Din4 => VN789_in4,
        Din5 => VN789_in5,
        VN2CN0_bit => VN_data_out(4734),
        VN2CN1_bit => VN_data_out(4735),
        VN2CN2_bit => VN_data_out(4736),
        VN2CN3_bit => VN_data_out(4737),
        VN2CN4_bit => VN_data_out(4738),
        VN2CN5_bit => VN_data_out(4739),
        VN2CN0_sign => VN_sign_out(4734),
        VN2CN1_sign => VN_sign_out(4735),
        VN2CN2_sign => VN_sign_out(4736),
        VN2CN3_sign => VN_sign_out(4737),
        VN2CN4_sign => VN_sign_out(4738),
        VN2CN5_sign => VN_sign_out(4739),
        codeword => codeword(789),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN790 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4745 downto 4740),
        Din0 => VN790_in0,
        Din1 => VN790_in1,
        Din2 => VN790_in2,
        Din3 => VN790_in3,
        Din4 => VN790_in4,
        Din5 => VN790_in5,
        VN2CN0_bit => VN_data_out(4740),
        VN2CN1_bit => VN_data_out(4741),
        VN2CN2_bit => VN_data_out(4742),
        VN2CN3_bit => VN_data_out(4743),
        VN2CN4_bit => VN_data_out(4744),
        VN2CN5_bit => VN_data_out(4745),
        VN2CN0_sign => VN_sign_out(4740),
        VN2CN1_sign => VN_sign_out(4741),
        VN2CN2_sign => VN_sign_out(4742),
        VN2CN3_sign => VN_sign_out(4743),
        VN2CN4_sign => VN_sign_out(4744),
        VN2CN5_sign => VN_sign_out(4745),
        codeword => codeword(790),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN791 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4751 downto 4746),
        Din0 => VN791_in0,
        Din1 => VN791_in1,
        Din2 => VN791_in2,
        Din3 => VN791_in3,
        Din4 => VN791_in4,
        Din5 => VN791_in5,
        VN2CN0_bit => VN_data_out(4746),
        VN2CN1_bit => VN_data_out(4747),
        VN2CN2_bit => VN_data_out(4748),
        VN2CN3_bit => VN_data_out(4749),
        VN2CN4_bit => VN_data_out(4750),
        VN2CN5_bit => VN_data_out(4751),
        VN2CN0_sign => VN_sign_out(4746),
        VN2CN1_sign => VN_sign_out(4747),
        VN2CN2_sign => VN_sign_out(4748),
        VN2CN3_sign => VN_sign_out(4749),
        VN2CN4_sign => VN_sign_out(4750),
        VN2CN5_sign => VN_sign_out(4751),
        codeword => codeword(791),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN792 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4757 downto 4752),
        Din0 => VN792_in0,
        Din1 => VN792_in1,
        Din2 => VN792_in2,
        Din3 => VN792_in3,
        Din4 => VN792_in4,
        Din5 => VN792_in5,
        VN2CN0_bit => VN_data_out(4752),
        VN2CN1_bit => VN_data_out(4753),
        VN2CN2_bit => VN_data_out(4754),
        VN2CN3_bit => VN_data_out(4755),
        VN2CN4_bit => VN_data_out(4756),
        VN2CN5_bit => VN_data_out(4757),
        VN2CN0_sign => VN_sign_out(4752),
        VN2CN1_sign => VN_sign_out(4753),
        VN2CN2_sign => VN_sign_out(4754),
        VN2CN3_sign => VN_sign_out(4755),
        VN2CN4_sign => VN_sign_out(4756),
        VN2CN5_sign => VN_sign_out(4757),
        codeword => codeword(792),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN793 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4763 downto 4758),
        Din0 => VN793_in0,
        Din1 => VN793_in1,
        Din2 => VN793_in2,
        Din3 => VN793_in3,
        Din4 => VN793_in4,
        Din5 => VN793_in5,
        VN2CN0_bit => VN_data_out(4758),
        VN2CN1_bit => VN_data_out(4759),
        VN2CN2_bit => VN_data_out(4760),
        VN2CN3_bit => VN_data_out(4761),
        VN2CN4_bit => VN_data_out(4762),
        VN2CN5_bit => VN_data_out(4763),
        VN2CN0_sign => VN_sign_out(4758),
        VN2CN1_sign => VN_sign_out(4759),
        VN2CN2_sign => VN_sign_out(4760),
        VN2CN3_sign => VN_sign_out(4761),
        VN2CN4_sign => VN_sign_out(4762),
        VN2CN5_sign => VN_sign_out(4763),
        codeword => codeword(793),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN794 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4769 downto 4764),
        Din0 => VN794_in0,
        Din1 => VN794_in1,
        Din2 => VN794_in2,
        Din3 => VN794_in3,
        Din4 => VN794_in4,
        Din5 => VN794_in5,
        VN2CN0_bit => VN_data_out(4764),
        VN2CN1_bit => VN_data_out(4765),
        VN2CN2_bit => VN_data_out(4766),
        VN2CN3_bit => VN_data_out(4767),
        VN2CN4_bit => VN_data_out(4768),
        VN2CN5_bit => VN_data_out(4769),
        VN2CN0_sign => VN_sign_out(4764),
        VN2CN1_sign => VN_sign_out(4765),
        VN2CN2_sign => VN_sign_out(4766),
        VN2CN3_sign => VN_sign_out(4767),
        VN2CN4_sign => VN_sign_out(4768),
        VN2CN5_sign => VN_sign_out(4769),
        codeword => codeword(794),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN795 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4775 downto 4770),
        Din0 => VN795_in0,
        Din1 => VN795_in1,
        Din2 => VN795_in2,
        Din3 => VN795_in3,
        Din4 => VN795_in4,
        Din5 => VN795_in5,
        VN2CN0_bit => VN_data_out(4770),
        VN2CN1_bit => VN_data_out(4771),
        VN2CN2_bit => VN_data_out(4772),
        VN2CN3_bit => VN_data_out(4773),
        VN2CN4_bit => VN_data_out(4774),
        VN2CN5_bit => VN_data_out(4775),
        VN2CN0_sign => VN_sign_out(4770),
        VN2CN1_sign => VN_sign_out(4771),
        VN2CN2_sign => VN_sign_out(4772),
        VN2CN3_sign => VN_sign_out(4773),
        VN2CN4_sign => VN_sign_out(4774),
        VN2CN5_sign => VN_sign_out(4775),
        codeword => codeword(795),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN796 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4781 downto 4776),
        Din0 => VN796_in0,
        Din1 => VN796_in1,
        Din2 => VN796_in2,
        Din3 => VN796_in3,
        Din4 => VN796_in4,
        Din5 => VN796_in5,
        VN2CN0_bit => VN_data_out(4776),
        VN2CN1_bit => VN_data_out(4777),
        VN2CN2_bit => VN_data_out(4778),
        VN2CN3_bit => VN_data_out(4779),
        VN2CN4_bit => VN_data_out(4780),
        VN2CN5_bit => VN_data_out(4781),
        VN2CN0_sign => VN_sign_out(4776),
        VN2CN1_sign => VN_sign_out(4777),
        VN2CN2_sign => VN_sign_out(4778),
        VN2CN3_sign => VN_sign_out(4779),
        VN2CN4_sign => VN_sign_out(4780),
        VN2CN5_sign => VN_sign_out(4781),
        codeword => codeword(796),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN797 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4787 downto 4782),
        Din0 => VN797_in0,
        Din1 => VN797_in1,
        Din2 => VN797_in2,
        Din3 => VN797_in3,
        Din4 => VN797_in4,
        Din5 => VN797_in5,
        VN2CN0_bit => VN_data_out(4782),
        VN2CN1_bit => VN_data_out(4783),
        VN2CN2_bit => VN_data_out(4784),
        VN2CN3_bit => VN_data_out(4785),
        VN2CN4_bit => VN_data_out(4786),
        VN2CN5_bit => VN_data_out(4787),
        VN2CN0_sign => VN_sign_out(4782),
        VN2CN1_sign => VN_sign_out(4783),
        VN2CN2_sign => VN_sign_out(4784),
        VN2CN3_sign => VN_sign_out(4785),
        VN2CN4_sign => VN_sign_out(4786),
        VN2CN5_sign => VN_sign_out(4787),
        codeword => codeword(797),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN798 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4793 downto 4788),
        Din0 => VN798_in0,
        Din1 => VN798_in1,
        Din2 => VN798_in2,
        Din3 => VN798_in3,
        Din4 => VN798_in4,
        Din5 => VN798_in5,
        VN2CN0_bit => VN_data_out(4788),
        VN2CN1_bit => VN_data_out(4789),
        VN2CN2_bit => VN_data_out(4790),
        VN2CN3_bit => VN_data_out(4791),
        VN2CN4_bit => VN_data_out(4792),
        VN2CN5_bit => VN_data_out(4793),
        VN2CN0_sign => VN_sign_out(4788),
        VN2CN1_sign => VN_sign_out(4789),
        VN2CN2_sign => VN_sign_out(4790),
        VN2CN3_sign => VN_sign_out(4791),
        VN2CN4_sign => VN_sign_out(4792),
        VN2CN5_sign => VN_sign_out(4793),
        codeword => codeword(798),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN799 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4799 downto 4794),
        Din0 => VN799_in0,
        Din1 => VN799_in1,
        Din2 => VN799_in2,
        Din3 => VN799_in3,
        Din4 => VN799_in4,
        Din5 => VN799_in5,
        VN2CN0_bit => VN_data_out(4794),
        VN2CN1_bit => VN_data_out(4795),
        VN2CN2_bit => VN_data_out(4796),
        VN2CN3_bit => VN_data_out(4797),
        VN2CN4_bit => VN_data_out(4798),
        VN2CN5_bit => VN_data_out(4799),
        VN2CN0_sign => VN_sign_out(4794),
        VN2CN1_sign => VN_sign_out(4795),
        VN2CN2_sign => VN_sign_out(4796),
        VN2CN3_sign => VN_sign_out(4797),
        VN2CN4_sign => VN_sign_out(4798),
        VN2CN5_sign => VN_sign_out(4799),
        codeword => codeword(799),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN800 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4805 downto 4800),
        Din0 => VN800_in0,
        Din1 => VN800_in1,
        Din2 => VN800_in2,
        Din3 => VN800_in3,
        Din4 => VN800_in4,
        Din5 => VN800_in5,
        VN2CN0_bit => VN_data_out(4800),
        VN2CN1_bit => VN_data_out(4801),
        VN2CN2_bit => VN_data_out(4802),
        VN2CN3_bit => VN_data_out(4803),
        VN2CN4_bit => VN_data_out(4804),
        VN2CN5_bit => VN_data_out(4805),
        VN2CN0_sign => VN_sign_out(4800),
        VN2CN1_sign => VN_sign_out(4801),
        VN2CN2_sign => VN_sign_out(4802),
        VN2CN3_sign => VN_sign_out(4803),
        VN2CN4_sign => VN_sign_out(4804),
        VN2CN5_sign => VN_sign_out(4805),
        codeword => codeword(800),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN801 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4811 downto 4806),
        Din0 => VN801_in0,
        Din1 => VN801_in1,
        Din2 => VN801_in2,
        Din3 => VN801_in3,
        Din4 => VN801_in4,
        Din5 => VN801_in5,
        VN2CN0_bit => VN_data_out(4806),
        VN2CN1_bit => VN_data_out(4807),
        VN2CN2_bit => VN_data_out(4808),
        VN2CN3_bit => VN_data_out(4809),
        VN2CN4_bit => VN_data_out(4810),
        VN2CN5_bit => VN_data_out(4811),
        VN2CN0_sign => VN_sign_out(4806),
        VN2CN1_sign => VN_sign_out(4807),
        VN2CN2_sign => VN_sign_out(4808),
        VN2CN3_sign => VN_sign_out(4809),
        VN2CN4_sign => VN_sign_out(4810),
        VN2CN5_sign => VN_sign_out(4811),
        codeword => codeword(801),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN802 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4817 downto 4812),
        Din0 => VN802_in0,
        Din1 => VN802_in1,
        Din2 => VN802_in2,
        Din3 => VN802_in3,
        Din4 => VN802_in4,
        Din5 => VN802_in5,
        VN2CN0_bit => VN_data_out(4812),
        VN2CN1_bit => VN_data_out(4813),
        VN2CN2_bit => VN_data_out(4814),
        VN2CN3_bit => VN_data_out(4815),
        VN2CN4_bit => VN_data_out(4816),
        VN2CN5_bit => VN_data_out(4817),
        VN2CN0_sign => VN_sign_out(4812),
        VN2CN1_sign => VN_sign_out(4813),
        VN2CN2_sign => VN_sign_out(4814),
        VN2CN3_sign => VN_sign_out(4815),
        VN2CN4_sign => VN_sign_out(4816),
        VN2CN5_sign => VN_sign_out(4817),
        codeword => codeword(802),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN803 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4823 downto 4818),
        Din0 => VN803_in0,
        Din1 => VN803_in1,
        Din2 => VN803_in2,
        Din3 => VN803_in3,
        Din4 => VN803_in4,
        Din5 => VN803_in5,
        VN2CN0_bit => VN_data_out(4818),
        VN2CN1_bit => VN_data_out(4819),
        VN2CN2_bit => VN_data_out(4820),
        VN2CN3_bit => VN_data_out(4821),
        VN2CN4_bit => VN_data_out(4822),
        VN2CN5_bit => VN_data_out(4823),
        VN2CN0_sign => VN_sign_out(4818),
        VN2CN1_sign => VN_sign_out(4819),
        VN2CN2_sign => VN_sign_out(4820),
        VN2CN3_sign => VN_sign_out(4821),
        VN2CN4_sign => VN_sign_out(4822),
        VN2CN5_sign => VN_sign_out(4823),
        codeword => codeword(803),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN804 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4829 downto 4824),
        Din0 => VN804_in0,
        Din1 => VN804_in1,
        Din2 => VN804_in2,
        Din3 => VN804_in3,
        Din4 => VN804_in4,
        Din5 => VN804_in5,
        VN2CN0_bit => VN_data_out(4824),
        VN2CN1_bit => VN_data_out(4825),
        VN2CN2_bit => VN_data_out(4826),
        VN2CN3_bit => VN_data_out(4827),
        VN2CN4_bit => VN_data_out(4828),
        VN2CN5_bit => VN_data_out(4829),
        VN2CN0_sign => VN_sign_out(4824),
        VN2CN1_sign => VN_sign_out(4825),
        VN2CN2_sign => VN_sign_out(4826),
        VN2CN3_sign => VN_sign_out(4827),
        VN2CN4_sign => VN_sign_out(4828),
        VN2CN5_sign => VN_sign_out(4829),
        codeword => codeword(804),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN805 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4835 downto 4830),
        Din0 => VN805_in0,
        Din1 => VN805_in1,
        Din2 => VN805_in2,
        Din3 => VN805_in3,
        Din4 => VN805_in4,
        Din5 => VN805_in5,
        VN2CN0_bit => VN_data_out(4830),
        VN2CN1_bit => VN_data_out(4831),
        VN2CN2_bit => VN_data_out(4832),
        VN2CN3_bit => VN_data_out(4833),
        VN2CN4_bit => VN_data_out(4834),
        VN2CN5_bit => VN_data_out(4835),
        VN2CN0_sign => VN_sign_out(4830),
        VN2CN1_sign => VN_sign_out(4831),
        VN2CN2_sign => VN_sign_out(4832),
        VN2CN3_sign => VN_sign_out(4833),
        VN2CN4_sign => VN_sign_out(4834),
        VN2CN5_sign => VN_sign_out(4835),
        codeword => codeword(805),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN806 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4841 downto 4836),
        Din0 => VN806_in0,
        Din1 => VN806_in1,
        Din2 => VN806_in2,
        Din3 => VN806_in3,
        Din4 => VN806_in4,
        Din5 => VN806_in5,
        VN2CN0_bit => VN_data_out(4836),
        VN2CN1_bit => VN_data_out(4837),
        VN2CN2_bit => VN_data_out(4838),
        VN2CN3_bit => VN_data_out(4839),
        VN2CN4_bit => VN_data_out(4840),
        VN2CN5_bit => VN_data_out(4841),
        VN2CN0_sign => VN_sign_out(4836),
        VN2CN1_sign => VN_sign_out(4837),
        VN2CN2_sign => VN_sign_out(4838),
        VN2CN3_sign => VN_sign_out(4839),
        VN2CN4_sign => VN_sign_out(4840),
        VN2CN5_sign => VN_sign_out(4841),
        codeword => codeword(806),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN807 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4847 downto 4842),
        Din0 => VN807_in0,
        Din1 => VN807_in1,
        Din2 => VN807_in2,
        Din3 => VN807_in3,
        Din4 => VN807_in4,
        Din5 => VN807_in5,
        VN2CN0_bit => VN_data_out(4842),
        VN2CN1_bit => VN_data_out(4843),
        VN2CN2_bit => VN_data_out(4844),
        VN2CN3_bit => VN_data_out(4845),
        VN2CN4_bit => VN_data_out(4846),
        VN2CN5_bit => VN_data_out(4847),
        VN2CN0_sign => VN_sign_out(4842),
        VN2CN1_sign => VN_sign_out(4843),
        VN2CN2_sign => VN_sign_out(4844),
        VN2CN3_sign => VN_sign_out(4845),
        VN2CN4_sign => VN_sign_out(4846),
        VN2CN5_sign => VN_sign_out(4847),
        codeword => codeword(807),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN808 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4853 downto 4848),
        Din0 => VN808_in0,
        Din1 => VN808_in1,
        Din2 => VN808_in2,
        Din3 => VN808_in3,
        Din4 => VN808_in4,
        Din5 => VN808_in5,
        VN2CN0_bit => VN_data_out(4848),
        VN2CN1_bit => VN_data_out(4849),
        VN2CN2_bit => VN_data_out(4850),
        VN2CN3_bit => VN_data_out(4851),
        VN2CN4_bit => VN_data_out(4852),
        VN2CN5_bit => VN_data_out(4853),
        VN2CN0_sign => VN_sign_out(4848),
        VN2CN1_sign => VN_sign_out(4849),
        VN2CN2_sign => VN_sign_out(4850),
        VN2CN3_sign => VN_sign_out(4851),
        VN2CN4_sign => VN_sign_out(4852),
        VN2CN5_sign => VN_sign_out(4853),
        codeword => codeword(808),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN809 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4859 downto 4854),
        Din0 => VN809_in0,
        Din1 => VN809_in1,
        Din2 => VN809_in2,
        Din3 => VN809_in3,
        Din4 => VN809_in4,
        Din5 => VN809_in5,
        VN2CN0_bit => VN_data_out(4854),
        VN2CN1_bit => VN_data_out(4855),
        VN2CN2_bit => VN_data_out(4856),
        VN2CN3_bit => VN_data_out(4857),
        VN2CN4_bit => VN_data_out(4858),
        VN2CN5_bit => VN_data_out(4859),
        VN2CN0_sign => VN_sign_out(4854),
        VN2CN1_sign => VN_sign_out(4855),
        VN2CN2_sign => VN_sign_out(4856),
        VN2CN3_sign => VN_sign_out(4857),
        VN2CN4_sign => VN_sign_out(4858),
        VN2CN5_sign => VN_sign_out(4859),
        codeword => codeword(809),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN810 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4865 downto 4860),
        Din0 => VN810_in0,
        Din1 => VN810_in1,
        Din2 => VN810_in2,
        Din3 => VN810_in3,
        Din4 => VN810_in4,
        Din5 => VN810_in5,
        VN2CN0_bit => VN_data_out(4860),
        VN2CN1_bit => VN_data_out(4861),
        VN2CN2_bit => VN_data_out(4862),
        VN2CN3_bit => VN_data_out(4863),
        VN2CN4_bit => VN_data_out(4864),
        VN2CN5_bit => VN_data_out(4865),
        VN2CN0_sign => VN_sign_out(4860),
        VN2CN1_sign => VN_sign_out(4861),
        VN2CN2_sign => VN_sign_out(4862),
        VN2CN3_sign => VN_sign_out(4863),
        VN2CN4_sign => VN_sign_out(4864),
        VN2CN5_sign => VN_sign_out(4865),
        codeword => codeword(810),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN811 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4871 downto 4866),
        Din0 => VN811_in0,
        Din1 => VN811_in1,
        Din2 => VN811_in2,
        Din3 => VN811_in3,
        Din4 => VN811_in4,
        Din5 => VN811_in5,
        VN2CN0_bit => VN_data_out(4866),
        VN2CN1_bit => VN_data_out(4867),
        VN2CN2_bit => VN_data_out(4868),
        VN2CN3_bit => VN_data_out(4869),
        VN2CN4_bit => VN_data_out(4870),
        VN2CN5_bit => VN_data_out(4871),
        VN2CN0_sign => VN_sign_out(4866),
        VN2CN1_sign => VN_sign_out(4867),
        VN2CN2_sign => VN_sign_out(4868),
        VN2CN3_sign => VN_sign_out(4869),
        VN2CN4_sign => VN_sign_out(4870),
        VN2CN5_sign => VN_sign_out(4871),
        codeword => codeword(811),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN812 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4877 downto 4872),
        Din0 => VN812_in0,
        Din1 => VN812_in1,
        Din2 => VN812_in2,
        Din3 => VN812_in3,
        Din4 => VN812_in4,
        Din5 => VN812_in5,
        VN2CN0_bit => VN_data_out(4872),
        VN2CN1_bit => VN_data_out(4873),
        VN2CN2_bit => VN_data_out(4874),
        VN2CN3_bit => VN_data_out(4875),
        VN2CN4_bit => VN_data_out(4876),
        VN2CN5_bit => VN_data_out(4877),
        VN2CN0_sign => VN_sign_out(4872),
        VN2CN1_sign => VN_sign_out(4873),
        VN2CN2_sign => VN_sign_out(4874),
        VN2CN3_sign => VN_sign_out(4875),
        VN2CN4_sign => VN_sign_out(4876),
        VN2CN5_sign => VN_sign_out(4877),
        codeword => codeword(812),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN813 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4883 downto 4878),
        Din0 => VN813_in0,
        Din1 => VN813_in1,
        Din2 => VN813_in2,
        Din3 => VN813_in3,
        Din4 => VN813_in4,
        Din5 => VN813_in5,
        VN2CN0_bit => VN_data_out(4878),
        VN2CN1_bit => VN_data_out(4879),
        VN2CN2_bit => VN_data_out(4880),
        VN2CN3_bit => VN_data_out(4881),
        VN2CN4_bit => VN_data_out(4882),
        VN2CN5_bit => VN_data_out(4883),
        VN2CN0_sign => VN_sign_out(4878),
        VN2CN1_sign => VN_sign_out(4879),
        VN2CN2_sign => VN_sign_out(4880),
        VN2CN3_sign => VN_sign_out(4881),
        VN2CN4_sign => VN_sign_out(4882),
        VN2CN5_sign => VN_sign_out(4883),
        codeword => codeword(813),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN814 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4889 downto 4884),
        Din0 => VN814_in0,
        Din1 => VN814_in1,
        Din2 => VN814_in2,
        Din3 => VN814_in3,
        Din4 => VN814_in4,
        Din5 => VN814_in5,
        VN2CN0_bit => VN_data_out(4884),
        VN2CN1_bit => VN_data_out(4885),
        VN2CN2_bit => VN_data_out(4886),
        VN2CN3_bit => VN_data_out(4887),
        VN2CN4_bit => VN_data_out(4888),
        VN2CN5_bit => VN_data_out(4889),
        VN2CN0_sign => VN_sign_out(4884),
        VN2CN1_sign => VN_sign_out(4885),
        VN2CN2_sign => VN_sign_out(4886),
        VN2CN3_sign => VN_sign_out(4887),
        VN2CN4_sign => VN_sign_out(4888),
        VN2CN5_sign => VN_sign_out(4889),
        codeword => codeword(814),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN815 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4895 downto 4890),
        Din0 => VN815_in0,
        Din1 => VN815_in1,
        Din2 => VN815_in2,
        Din3 => VN815_in3,
        Din4 => VN815_in4,
        Din5 => VN815_in5,
        VN2CN0_bit => VN_data_out(4890),
        VN2CN1_bit => VN_data_out(4891),
        VN2CN2_bit => VN_data_out(4892),
        VN2CN3_bit => VN_data_out(4893),
        VN2CN4_bit => VN_data_out(4894),
        VN2CN5_bit => VN_data_out(4895),
        VN2CN0_sign => VN_sign_out(4890),
        VN2CN1_sign => VN_sign_out(4891),
        VN2CN2_sign => VN_sign_out(4892),
        VN2CN3_sign => VN_sign_out(4893),
        VN2CN4_sign => VN_sign_out(4894),
        VN2CN5_sign => VN_sign_out(4895),
        codeword => codeword(815),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN816 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4901 downto 4896),
        Din0 => VN816_in0,
        Din1 => VN816_in1,
        Din2 => VN816_in2,
        Din3 => VN816_in3,
        Din4 => VN816_in4,
        Din5 => VN816_in5,
        VN2CN0_bit => VN_data_out(4896),
        VN2CN1_bit => VN_data_out(4897),
        VN2CN2_bit => VN_data_out(4898),
        VN2CN3_bit => VN_data_out(4899),
        VN2CN4_bit => VN_data_out(4900),
        VN2CN5_bit => VN_data_out(4901),
        VN2CN0_sign => VN_sign_out(4896),
        VN2CN1_sign => VN_sign_out(4897),
        VN2CN2_sign => VN_sign_out(4898),
        VN2CN3_sign => VN_sign_out(4899),
        VN2CN4_sign => VN_sign_out(4900),
        VN2CN5_sign => VN_sign_out(4901),
        codeword => codeword(816),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN817 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4907 downto 4902),
        Din0 => VN817_in0,
        Din1 => VN817_in1,
        Din2 => VN817_in2,
        Din3 => VN817_in3,
        Din4 => VN817_in4,
        Din5 => VN817_in5,
        VN2CN0_bit => VN_data_out(4902),
        VN2CN1_bit => VN_data_out(4903),
        VN2CN2_bit => VN_data_out(4904),
        VN2CN3_bit => VN_data_out(4905),
        VN2CN4_bit => VN_data_out(4906),
        VN2CN5_bit => VN_data_out(4907),
        VN2CN0_sign => VN_sign_out(4902),
        VN2CN1_sign => VN_sign_out(4903),
        VN2CN2_sign => VN_sign_out(4904),
        VN2CN3_sign => VN_sign_out(4905),
        VN2CN4_sign => VN_sign_out(4906),
        VN2CN5_sign => VN_sign_out(4907),
        codeword => codeword(817),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN818 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4913 downto 4908),
        Din0 => VN818_in0,
        Din1 => VN818_in1,
        Din2 => VN818_in2,
        Din3 => VN818_in3,
        Din4 => VN818_in4,
        Din5 => VN818_in5,
        VN2CN0_bit => VN_data_out(4908),
        VN2CN1_bit => VN_data_out(4909),
        VN2CN2_bit => VN_data_out(4910),
        VN2CN3_bit => VN_data_out(4911),
        VN2CN4_bit => VN_data_out(4912),
        VN2CN5_bit => VN_data_out(4913),
        VN2CN0_sign => VN_sign_out(4908),
        VN2CN1_sign => VN_sign_out(4909),
        VN2CN2_sign => VN_sign_out(4910),
        VN2CN3_sign => VN_sign_out(4911),
        VN2CN4_sign => VN_sign_out(4912),
        VN2CN5_sign => VN_sign_out(4913),
        codeword => codeword(818),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN819 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4919 downto 4914),
        Din0 => VN819_in0,
        Din1 => VN819_in1,
        Din2 => VN819_in2,
        Din3 => VN819_in3,
        Din4 => VN819_in4,
        Din5 => VN819_in5,
        VN2CN0_bit => VN_data_out(4914),
        VN2CN1_bit => VN_data_out(4915),
        VN2CN2_bit => VN_data_out(4916),
        VN2CN3_bit => VN_data_out(4917),
        VN2CN4_bit => VN_data_out(4918),
        VN2CN5_bit => VN_data_out(4919),
        VN2CN0_sign => VN_sign_out(4914),
        VN2CN1_sign => VN_sign_out(4915),
        VN2CN2_sign => VN_sign_out(4916),
        VN2CN3_sign => VN_sign_out(4917),
        VN2CN4_sign => VN_sign_out(4918),
        VN2CN5_sign => VN_sign_out(4919),
        codeword => codeword(819),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN820 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4925 downto 4920),
        Din0 => VN820_in0,
        Din1 => VN820_in1,
        Din2 => VN820_in2,
        Din3 => VN820_in3,
        Din4 => VN820_in4,
        Din5 => VN820_in5,
        VN2CN0_bit => VN_data_out(4920),
        VN2CN1_bit => VN_data_out(4921),
        VN2CN2_bit => VN_data_out(4922),
        VN2CN3_bit => VN_data_out(4923),
        VN2CN4_bit => VN_data_out(4924),
        VN2CN5_bit => VN_data_out(4925),
        VN2CN0_sign => VN_sign_out(4920),
        VN2CN1_sign => VN_sign_out(4921),
        VN2CN2_sign => VN_sign_out(4922),
        VN2CN3_sign => VN_sign_out(4923),
        VN2CN4_sign => VN_sign_out(4924),
        VN2CN5_sign => VN_sign_out(4925),
        codeword => codeword(820),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN821 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4931 downto 4926),
        Din0 => VN821_in0,
        Din1 => VN821_in1,
        Din2 => VN821_in2,
        Din3 => VN821_in3,
        Din4 => VN821_in4,
        Din5 => VN821_in5,
        VN2CN0_bit => VN_data_out(4926),
        VN2CN1_bit => VN_data_out(4927),
        VN2CN2_bit => VN_data_out(4928),
        VN2CN3_bit => VN_data_out(4929),
        VN2CN4_bit => VN_data_out(4930),
        VN2CN5_bit => VN_data_out(4931),
        VN2CN0_sign => VN_sign_out(4926),
        VN2CN1_sign => VN_sign_out(4927),
        VN2CN2_sign => VN_sign_out(4928),
        VN2CN3_sign => VN_sign_out(4929),
        VN2CN4_sign => VN_sign_out(4930),
        VN2CN5_sign => VN_sign_out(4931),
        codeword => codeword(821),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN822 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4937 downto 4932),
        Din0 => VN822_in0,
        Din1 => VN822_in1,
        Din2 => VN822_in2,
        Din3 => VN822_in3,
        Din4 => VN822_in4,
        Din5 => VN822_in5,
        VN2CN0_bit => VN_data_out(4932),
        VN2CN1_bit => VN_data_out(4933),
        VN2CN2_bit => VN_data_out(4934),
        VN2CN3_bit => VN_data_out(4935),
        VN2CN4_bit => VN_data_out(4936),
        VN2CN5_bit => VN_data_out(4937),
        VN2CN0_sign => VN_sign_out(4932),
        VN2CN1_sign => VN_sign_out(4933),
        VN2CN2_sign => VN_sign_out(4934),
        VN2CN3_sign => VN_sign_out(4935),
        VN2CN4_sign => VN_sign_out(4936),
        VN2CN5_sign => VN_sign_out(4937),
        codeword => codeword(822),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN823 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4943 downto 4938),
        Din0 => VN823_in0,
        Din1 => VN823_in1,
        Din2 => VN823_in2,
        Din3 => VN823_in3,
        Din4 => VN823_in4,
        Din5 => VN823_in5,
        VN2CN0_bit => VN_data_out(4938),
        VN2CN1_bit => VN_data_out(4939),
        VN2CN2_bit => VN_data_out(4940),
        VN2CN3_bit => VN_data_out(4941),
        VN2CN4_bit => VN_data_out(4942),
        VN2CN5_bit => VN_data_out(4943),
        VN2CN0_sign => VN_sign_out(4938),
        VN2CN1_sign => VN_sign_out(4939),
        VN2CN2_sign => VN_sign_out(4940),
        VN2CN3_sign => VN_sign_out(4941),
        VN2CN4_sign => VN_sign_out(4942),
        VN2CN5_sign => VN_sign_out(4943),
        codeword => codeword(823),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN824 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4949 downto 4944),
        Din0 => VN824_in0,
        Din1 => VN824_in1,
        Din2 => VN824_in2,
        Din3 => VN824_in3,
        Din4 => VN824_in4,
        Din5 => VN824_in5,
        VN2CN0_bit => VN_data_out(4944),
        VN2CN1_bit => VN_data_out(4945),
        VN2CN2_bit => VN_data_out(4946),
        VN2CN3_bit => VN_data_out(4947),
        VN2CN4_bit => VN_data_out(4948),
        VN2CN5_bit => VN_data_out(4949),
        VN2CN0_sign => VN_sign_out(4944),
        VN2CN1_sign => VN_sign_out(4945),
        VN2CN2_sign => VN_sign_out(4946),
        VN2CN3_sign => VN_sign_out(4947),
        VN2CN4_sign => VN_sign_out(4948),
        VN2CN5_sign => VN_sign_out(4949),
        codeword => codeword(824),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN825 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4955 downto 4950),
        Din0 => VN825_in0,
        Din1 => VN825_in1,
        Din2 => VN825_in2,
        Din3 => VN825_in3,
        Din4 => VN825_in4,
        Din5 => VN825_in5,
        VN2CN0_bit => VN_data_out(4950),
        VN2CN1_bit => VN_data_out(4951),
        VN2CN2_bit => VN_data_out(4952),
        VN2CN3_bit => VN_data_out(4953),
        VN2CN4_bit => VN_data_out(4954),
        VN2CN5_bit => VN_data_out(4955),
        VN2CN0_sign => VN_sign_out(4950),
        VN2CN1_sign => VN_sign_out(4951),
        VN2CN2_sign => VN_sign_out(4952),
        VN2CN3_sign => VN_sign_out(4953),
        VN2CN4_sign => VN_sign_out(4954),
        VN2CN5_sign => VN_sign_out(4955),
        codeword => codeword(825),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN826 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4961 downto 4956),
        Din0 => VN826_in0,
        Din1 => VN826_in1,
        Din2 => VN826_in2,
        Din3 => VN826_in3,
        Din4 => VN826_in4,
        Din5 => VN826_in5,
        VN2CN0_bit => VN_data_out(4956),
        VN2CN1_bit => VN_data_out(4957),
        VN2CN2_bit => VN_data_out(4958),
        VN2CN3_bit => VN_data_out(4959),
        VN2CN4_bit => VN_data_out(4960),
        VN2CN5_bit => VN_data_out(4961),
        VN2CN0_sign => VN_sign_out(4956),
        VN2CN1_sign => VN_sign_out(4957),
        VN2CN2_sign => VN_sign_out(4958),
        VN2CN3_sign => VN_sign_out(4959),
        VN2CN4_sign => VN_sign_out(4960),
        VN2CN5_sign => VN_sign_out(4961),
        codeword => codeword(826),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN827 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4967 downto 4962),
        Din0 => VN827_in0,
        Din1 => VN827_in1,
        Din2 => VN827_in2,
        Din3 => VN827_in3,
        Din4 => VN827_in4,
        Din5 => VN827_in5,
        VN2CN0_bit => VN_data_out(4962),
        VN2CN1_bit => VN_data_out(4963),
        VN2CN2_bit => VN_data_out(4964),
        VN2CN3_bit => VN_data_out(4965),
        VN2CN4_bit => VN_data_out(4966),
        VN2CN5_bit => VN_data_out(4967),
        VN2CN0_sign => VN_sign_out(4962),
        VN2CN1_sign => VN_sign_out(4963),
        VN2CN2_sign => VN_sign_out(4964),
        VN2CN3_sign => VN_sign_out(4965),
        VN2CN4_sign => VN_sign_out(4966),
        VN2CN5_sign => VN_sign_out(4967),
        codeword => codeword(827),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN828 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4973 downto 4968),
        Din0 => VN828_in0,
        Din1 => VN828_in1,
        Din2 => VN828_in2,
        Din3 => VN828_in3,
        Din4 => VN828_in4,
        Din5 => VN828_in5,
        VN2CN0_bit => VN_data_out(4968),
        VN2CN1_bit => VN_data_out(4969),
        VN2CN2_bit => VN_data_out(4970),
        VN2CN3_bit => VN_data_out(4971),
        VN2CN4_bit => VN_data_out(4972),
        VN2CN5_bit => VN_data_out(4973),
        VN2CN0_sign => VN_sign_out(4968),
        VN2CN1_sign => VN_sign_out(4969),
        VN2CN2_sign => VN_sign_out(4970),
        VN2CN3_sign => VN_sign_out(4971),
        VN2CN4_sign => VN_sign_out(4972),
        VN2CN5_sign => VN_sign_out(4973),
        codeword => codeword(828),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN829 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4979 downto 4974),
        Din0 => VN829_in0,
        Din1 => VN829_in1,
        Din2 => VN829_in2,
        Din3 => VN829_in3,
        Din4 => VN829_in4,
        Din5 => VN829_in5,
        VN2CN0_bit => VN_data_out(4974),
        VN2CN1_bit => VN_data_out(4975),
        VN2CN2_bit => VN_data_out(4976),
        VN2CN3_bit => VN_data_out(4977),
        VN2CN4_bit => VN_data_out(4978),
        VN2CN5_bit => VN_data_out(4979),
        VN2CN0_sign => VN_sign_out(4974),
        VN2CN1_sign => VN_sign_out(4975),
        VN2CN2_sign => VN_sign_out(4976),
        VN2CN3_sign => VN_sign_out(4977),
        VN2CN4_sign => VN_sign_out(4978),
        VN2CN5_sign => VN_sign_out(4979),
        codeword => codeword(829),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN830 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4985 downto 4980),
        Din0 => VN830_in0,
        Din1 => VN830_in1,
        Din2 => VN830_in2,
        Din3 => VN830_in3,
        Din4 => VN830_in4,
        Din5 => VN830_in5,
        VN2CN0_bit => VN_data_out(4980),
        VN2CN1_bit => VN_data_out(4981),
        VN2CN2_bit => VN_data_out(4982),
        VN2CN3_bit => VN_data_out(4983),
        VN2CN4_bit => VN_data_out(4984),
        VN2CN5_bit => VN_data_out(4985),
        VN2CN0_sign => VN_sign_out(4980),
        VN2CN1_sign => VN_sign_out(4981),
        VN2CN2_sign => VN_sign_out(4982),
        VN2CN3_sign => VN_sign_out(4983),
        VN2CN4_sign => VN_sign_out(4984),
        VN2CN5_sign => VN_sign_out(4985),
        codeword => codeword(830),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN831 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4991 downto 4986),
        Din0 => VN831_in0,
        Din1 => VN831_in1,
        Din2 => VN831_in2,
        Din3 => VN831_in3,
        Din4 => VN831_in4,
        Din5 => VN831_in5,
        VN2CN0_bit => VN_data_out(4986),
        VN2CN1_bit => VN_data_out(4987),
        VN2CN2_bit => VN_data_out(4988),
        VN2CN3_bit => VN_data_out(4989),
        VN2CN4_bit => VN_data_out(4990),
        VN2CN5_bit => VN_data_out(4991),
        VN2CN0_sign => VN_sign_out(4986),
        VN2CN1_sign => VN_sign_out(4987),
        VN2CN2_sign => VN_sign_out(4988),
        VN2CN3_sign => VN_sign_out(4989),
        VN2CN4_sign => VN_sign_out(4990),
        VN2CN5_sign => VN_sign_out(4991),
        codeword => codeword(831),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN832 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(4997 downto 4992),
        Din0 => VN832_in0,
        Din1 => VN832_in1,
        Din2 => VN832_in2,
        Din3 => VN832_in3,
        Din4 => VN832_in4,
        Din5 => VN832_in5,
        VN2CN0_bit => VN_data_out(4992),
        VN2CN1_bit => VN_data_out(4993),
        VN2CN2_bit => VN_data_out(4994),
        VN2CN3_bit => VN_data_out(4995),
        VN2CN4_bit => VN_data_out(4996),
        VN2CN5_bit => VN_data_out(4997),
        VN2CN0_sign => VN_sign_out(4992),
        VN2CN1_sign => VN_sign_out(4993),
        VN2CN2_sign => VN_sign_out(4994),
        VN2CN3_sign => VN_sign_out(4995),
        VN2CN4_sign => VN_sign_out(4996),
        VN2CN5_sign => VN_sign_out(4997),
        codeword => codeword(832),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN833 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5003 downto 4998),
        Din0 => VN833_in0,
        Din1 => VN833_in1,
        Din2 => VN833_in2,
        Din3 => VN833_in3,
        Din4 => VN833_in4,
        Din5 => VN833_in5,
        VN2CN0_bit => VN_data_out(4998),
        VN2CN1_bit => VN_data_out(4999),
        VN2CN2_bit => VN_data_out(5000),
        VN2CN3_bit => VN_data_out(5001),
        VN2CN4_bit => VN_data_out(5002),
        VN2CN5_bit => VN_data_out(5003),
        VN2CN0_sign => VN_sign_out(4998),
        VN2CN1_sign => VN_sign_out(4999),
        VN2CN2_sign => VN_sign_out(5000),
        VN2CN3_sign => VN_sign_out(5001),
        VN2CN4_sign => VN_sign_out(5002),
        VN2CN5_sign => VN_sign_out(5003),
        codeword => codeword(833),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN834 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5009 downto 5004),
        Din0 => VN834_in0,
        Din1 => VN834_in1,
        Din2 => VN834_in2,
        Din3 => VN834_in3,
        Din4 => VN834_in4,
        Din5 => VN834_in5,
        VN2CN0_bit => VN_data_out(5004),
        VN2CN1_bit => VN_data_out(5005),
        VN2CN2_bit => VN_data_out(5006),
        VN2CN3_bit => VN_data_out(5007),
        VN2CN4_bit => VN_data_out(5008),
        VN2CN5_bit => VN_data_out(5009),
        VN2CN0_sign => VN_sign_out(5004),
        VN2CN1_sign => VN_sign_out(5005),
        VN2CN2_sign => VN_sign_out(5006),
        VN2CN3_sign => VN_sign_out(5007),
        VN2CN4_sign => VN_sign_out(5008),
        VN2CN5_sign => VN_sign_out(5009),
        codeword => codeword(834),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN835 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5015 downto 5010),
        Din0 => VN835_in0,
        Din1 => VN835_in1,
        Din2 => VN835_in2,
        Din3 => VN835_in3,
        Din4 => VN835_in4,
        Din5 => VN835_in5,
        VN2CN0_bit => VN_data_out(5010),
        VN2CN1_bit => VN_data_out(5011),
        VN2CN2_bit => VN_data_out(5012),
        VN2CN3_bit => VN_data_out(5013),
        VN2CN4_bit => VN_data_out(5014),
        VN2CN5_bit => VN_data_out(5015),
        VN2CN0_sign => VN_sign_out(5010),
        VN2CN1_sign => VN_sign_out(5011),
        VN2CN2_sign => VN_sign_out(5012),
        VN2CN3_sign => VN_sign_out(5013),
        VN2CN4_sign => VN_sign_out(5014),
        VN2CN5_sign => VN_sign_out(5015),
        codeword => codeword(835),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN836 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5021 downto 5016),
        Din0 => VN836_in0,
        Din1 => VN836_in1,
        Din2 => VN836_in2,
        Din3 => VN836_in3,
        Din4 => VN836_in4,
        Din5 => VN836_in5,
        VN2CN0_bit => VN_data_out(5016),
        VN2CN1_bit => VN_data_out(5017),
        VN2CN2_bit => VN_data_out(5018),
        VN2CN3_bit => VN_data_out(5019),
        VN2CN4_bit => VN_data_out(5020),
        VN2CN5_bit => VN_data_out(5021),
        VN2CN0_sign => VN_sign_out(5016),
        VN2CN1_sign => VN_sign_out(5017),
        VN2CN2_sign => VN_sign_out(5018),
        VN2CN3_sign => VN_sign_out(5019),
        VN2CN4_sign => VN_sign_out(5020),
        VN2CN5_sign => VN_sign_out(5021),
        codeword => codeword(836),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN837 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5027 downto 5022),
        Din0 => VN837_in0,
        Din1 => VN837_in1,
        Din2 => VN837_in2,
        Din3 => VN837_in3,
        Din4 => VN837_in4,
        Din5 => VN837_in5,
        VN2CN0_bit => VN_data_out(5022),
        VN2CN1_bit => VN_data_out(5023),
        VN2CN2_bit => VN_data_out(5024),
        VN2CN3_bit => VN_data_out(5025),
        VN2CN4_bit => VN_data_out(5026),
        VN2CN5_bit => VN_data_out(5027),
        VN2CN0_sign => VN_sign_out(5022),
        VN2CN1_sign => VN_sign_out(5023),
        VN2CN2_sign => VN_sign_out(5024),
        VN2CN3_sign => VN_sign_out(5025),
        VN2CN4_sign => VN_sign_out(5026),
        VN2CN5_sign => VN_sign_out(5027),
        codeword => codeword(837),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN838 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5033 downto 5028),
        Din0 => VN838_in0,
        Din1 => VN838_in1,
        Din2 => VN838_in2,
        Din3 => VN838_in3,
        Din4 => VN838_in4,
        Din5 => VN838_in5,
        VN2CN0_bit => VN_data_out(5028),
        VN2CN1_bit => VN_data_out(5029),
        VN2CN2_bit => VN_data_out(5030),
        VN2CN3_bit => VN_data_out(5031),
        VN2CN4_bit => VN_data_out(5032),
        VN2CN5_bit => VN_data_out(5033),
        VN2CN0_sign => VN_sign_out(5028),
        VN2CN1_sign => VN_sign_out(5029),
        VN2CN2_sign => VN_sign_out(5030),
        VN2CN3_sign => VN_sign_out(5031),
        VN2CN4_sign => VN_sign_out(5032),
        VN2CN5_sign => VN_sign_out(5033),
        codeword => codeword(838),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN839 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5039 downto 5034),
        Din0 => VN839_in0,
        Din1 => VN839_in1,
        Din2 => VN839_in2,
        Din3 => VN839_in3,
        Din4 => VN839_in4,
        Din5 => VN839_in5,
        VN2CN0_bit => VN_data_out(5034),
        VN2CN1_bit => VN_data_out(5035),
        VN2CN2_bit => VN_data_out(5036),
        VN2CN3_bit => VN_data_out(5037),
        VN2CN4_bit => VN_data_out(5038),
        VN2CN5_bit => VN_data_out(5039),
        VN2CN0_sign => VN_sign_out(5034),
        VN2CN1_sign => VN_sign_out(5035),
        VN2CN2_sign => VN_sign_out(5036),
        VN2CN3_sign => VN_sign_out(5037),
        VN2CN4_sign => VN_sign_out(5038),
        VN2CN5_sign => VN_sign_out(5039),
        codeword => codeword(839),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN840 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5045 downto 5040),
        Din0 => VN840_in0,
        Din1 => VN840_in1,
        Din2 => VN840_in2,
        Din3 => VN840_in3,
        Din4 => VN840_in4,
        Din5 => VN840_in5,
        VN2CN0_bit => VN_data_out(5040),
        VN2CN1_bit => VN_data_out(5041),
        VN2CN2_bit => VN_data_out(5042),
        VN2CN3_bit => VN_data_out(5043),
        VN2CN4_bit => VN_data_out(5044),
        VN2CN5_bit => VN_data_out(5045),
        VN2CN0_sign => VN_sign_out(5040),
        VN2CN1_sign => VN_sign_out(5041),
        VN2CN2_sign => VN_sign_out(5042),
        VN2CN3_sign => VN_sign_out(5043),
        VN2CN4_sign => VN_sign_out(5044),
        VN2CN5_sign => VN_sign_out(5045),
        codeword => codeword(840),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN841 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5051 downto 5046),
        Din0 => VN841_in0,
        Din1 => VN841_in1,
        Din2 => VN841_in2,
        Din3 => VN841_in3,
        Din4 => VN841_in4,
        Din5 => VN841_in5,
        VN2CN0_bit => VN_data_out(5046),
        VN2CN1_bit => VN_data_out(5047),
        VN2CN2_bit => VN_data_out(5048),
        VN2CN3_bit => VN_data_out(5049),
        VN2CN4_bit => VN_data_out(5050),
        VN2CN5_bit => VN_data_out(5051),
        VN2CN0_sign => VN_sign_out(5046),
        VN2CN1_sign => VN_sign_out(5047),
        VN2CN2_sign => VN_sign_out(5048),
        VN2CN3_sign => VN_sign_out(5049),
        VN2CN4_sign => VN_sign_out(5050),
        VN2CN5_sign => VN_sign_out(5051),
        codeword => codeword(841),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN842 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5057 downto 5052),
        Din0 => VN842_in0,
        Din1 => VN842_in1,
        Din2 => VN842_in2,
        Din3 => VN842_in3,
        Din4 => VN842_in4,
        Din5 => VN842_in5,
        VN2CN0_bit => VN_data_out(5052),
        VN2CN1_bit => VN_data_out(5053),
        VN2CN2_bit => VN_data_out(5054),
        VN2CN3_bit => VN_data_out(5055),
        VN2CN4_bit => VN_data_out(5056),
        VN2CN5_bit => VN_data_out(5057),
        VN2CN0_sign => VN_sign_out(5052),
        VN2CN1_sign => VN_sign_out(5053),
        VN2CN2_sign => VN_sign_out(5054),
        VN2CN3_sign => VN_sign_out(5055),
        VN2CN4_sign => VN_sign_out(5056),
        VN2CN5_sign => VN_sign_out(5057),
        codeword => codeword(842),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN843 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5063 downto 5058),
        Din0 => VN843_in0,
        Din1 => VN843_in1,
        Din2 => VN843_in2,
        Din3 => VN843_in3,
        Din4 => VN843_in4,
        Din5 => VN843_in5,
        VN2CN0_bit => VN_data_out(5058),
        VN2CN1_bit => VN_data_out(5059),
        VN2CN2_bit => VN_data_out(5060),
        VN2CN3_bit => VN_data_out(5061),
        VN2CN4_bit => VN_data_out(5062),
        VN2CN5_bit => VN_data_out(5063),
        VN2CN0_sign => VN_sign_out(5058),
        VN2CN1_sign => VN_sign_out(5059),
        VN2CN2_sign => VN_sign_out(5060),
        VN2CN3_sign => VN_sign_out(5061),
        VN2CN4_sign => VN_sign_out(5062),
        VN2CN5_sign => VN_sign_out(5063),
        codeword => codeword(843),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN844 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5069 downto 5064),
        Din0 => VN844_in0,
        Din1 => VN844_in1,
        Din2 => VN844_in2,
        Din3 => VN844_in3,
        Din4 => VN844_in4,
        Din5 => VN844_in5,
        VN2CN0_bit => VN_data_out(5064),
        VN2CN1_bit => VN_data_out(5065),
        VN2CN2_bit => VN_data_out(5066),
        VN2CN3_bit => VN_data_out(5067),
        VN2CN4_bit => VN_data_out(5068),
        VN2CN5_bit => VN_data_out(5069),
        VN2CN0_sign => VN_sign_out(5064),
        VN2CN1_sign => VN_sign_out(5065),
        VN2CN2_sign => VN_sign_out(5066),
        VN2CN3_sign => VN_sign_out(5067),
        VN2CN4_sign => VN_sign_out(5068),
        VN2CN5_sign => VN_sign_out(5069),
        codeword => codeword(844),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN845 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5075 downto 5070),
        Din0 => VN845_in0,
        Din1 => VN845_in1,
        Din2 => VN845_in2,
        Din3 => VN845_in3,
        Din4 => VN845_in4,
        Din5 => VN845_in5,
        VN2CN0_bit => VN_data_out(5070),
        VN2CN1_bit => VN_data_out(5071),
        VN2CN2_bit => VN_data_out(5072),
        VN2CN3_bit => VN_data_out(5073),
        VN2CN4_bit => VN_data_out(5074),
        VN2CN5_bit => VN_data_out(5075),
        VN2CN0_sign => VN_sign_out(5070),
        VN2CN1_sign => VN_sign_out(5071),
        VN2CN2_sign => VN_sign_out(5072),
        VN2CN3_sign => VN_sign_out(5073),
        VN2CN4_sign => VN_sign_out(5074),
        VN2CN5_sign => VN_sign_out(5075),
        codeword => codeword(845),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN846 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5081 downto 5076),
        Din0 => VN846_in0,
        Din1 => VN846_in1,
        Din2 => VN846_in2,
        Din3 => VN846_in3,
        Din4 => VN846_in4,
        Din5 => VN846_in5,
        VN2CN0_bit => VN_data_out(5076),
        VN2CN1_bit => VN_data_out(5077),
        VN2CN2_bit => VN_data_out(5078),
        VN2CN3_bit => VN_data_out(5079),
        VN2CN4_bit => VN_data_out(5080),
        VN2CN5_bit => VN_data_out(5081),
        VN2CN0_sign => VN_sign_out(5076),
        VN2CN1_sign => VN_sign_out(5077),
        VN2CN2_sign => VN_sign_out(5078),
        VN2CN3_sign => VN_sign_out(5079),
        VN2CN4_sign => VN_sign_out(5080),
        VN2CN5_sign => VN_sign_out(5081),
        codeword => codeword(846),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN847 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5087 downto 5082),
        Din0 => VN847_in0,
        Din1 => VN847_in1,
        Din2 => VN847_in2,
        Din3 => VN847_in3,
        Din4 => VN847_in4,
        Din5 => VN847_in5,
        VN2CN0_bit => VN_data_out(5082),
        VN2CN1_bit => VN_data_out(5083),
        VN2CN2_bit => VN_data_out(5084),
        VN2CN3_bit => VN_data_out(5085),
        VN2CN4_bit => VN_data_out(5086),
        VN2CN5_bit => VN_data_out(5087),
        VN2CN0_sign => VN_sign_out(5082),
        VN2CN1_sign => VN_sign_out(5083),
        VN2CN2_sign => VN_sign_out(5084),
        VN2CN3_sign => VN_sign_out(5085),
        VN2CN4_sign => VN_sign_out(5086),
        VN2CN5_sign => VN_sign_out(5087),
        codeword => codeword(847),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN848 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5093 downto 5088),
        Din0 => VN848_in0,
        Din1 => VN848_in1,
        Din2 => VN848_in2,
        Din3 => VN848_in3,
        Din4 => VN848_in4,
        Din5 => VN848_in5,
        VN2CN0_bit => VN_data_out(5088),
        VN2CN1_bit => VN_data_out(5089),
        VN2CN2_bit => VN_data_out(5090),
        VN2CN3_bit => VN_data_out(5091),
        VN2CN4_bit => VN_data_out(5092),
        VN2CN5_bit => VN_data_out(5093),
        VN2CN0_sign => VN_sign_out(5088),
        VN2CN1_sign => VN_sign_out(5089),
        VN2CN2_sign => VN_sign_out(5090),
        VN2CN3_sign => VN_sign_out(5091),
        VN2CN4_sign => VN_sign_out(5092),
        VN2CN5_sign => VN_sign_out(5093),
        codeword => codeword(848),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN849 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5099 downto 5094),
        Din0 => VN849_in0,
        Din1 => VN849_in1,
        Din2 => VN849_in2,
        Din3 => VN849_in3,
        Din4 => VN849_in4,
        Din5 => VN849_in5,
        VN2CN0_bit => VN_data_out(5094),
        VN2CN1_bit => VN_data_out(5095),
        VN2CN2_bit => VN_data_out(5096),
        VN2CN3_bit => VN_data_out(5097),
        VN2CN4_bit => VN_data_out(5098),
        VN2CN5_bit => VN_data_out(5099),
        VN2CN0_sign => VN_sign_out(5094),
        VN2CN1_sign => VN_sign_out(5095),
        VN2CN2_sign => VN_sign_out(5096),
        VN2CN3_sign => VN_sign_out(5097),
        VN2CN4_sign => VN_sign_out(5098),
        VN2CN5_sign => VN_sign_out(5099),
        codeword => codeword(849),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN850 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5105 downto 5100),
        Din0 => VN850_in0,
        Din1 => VN850_in1,
        Din2 => VN850_in2,
        Din3 => VN850_in3,
        Din4 => VN850_in4,
        Din5 => VN850_in5,
        VN2CN0_bit => VN_data_out(5100),
        VN2CN1_bit => VN_data_out(5101),
        VN2CN2_bit => VN_data_out(5102),
        VN2CN3_bit => VN_data_out(5103),
        VN2CN4_bit => VN_data_out(5104),
        VN2CN5_bit => VN_data_out(5105),
        VN2CN0_sign => VN_sign_out(5100),
        VN2CN1_sign => VN_sign_out(5101),
        VN2CN2_sign => VN_sign_out(5102),
        VN2CN3_sign => VN_sign_out(5103),
        VN2CN4_sign => VN_sign_out(5104),
        VN2CN5_sign => VN_sign_out(5105),
        codeword => codeword(850),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN851 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5111 downto 5106),
        Din0 => VN851_in0,
        Din1 => VN851_in1,
        Din2 => VN851_in2,
        Din3 => VN851_in3,
        Din4 => VN851_in4,
        Din5 => VN851_in5,
        VN2CN0_bit => VN_data_out(5106),
        VN2CN1_bit => VN_data_out(5107),
        VN2CN2_bit => VN_data_out(5108),
        VN2CN3_bit => VN_data_out(5109),
        VN2CN4_bit => VN_data_out(5110),
        VN2CN5_bit => VN_data_out(5111),
        VN2CN0_sign => VN_sign_out(5106),
        VN2CN1_sign => VN_sign_out(5107),
        VN2CN2_sign => VN_sign_out(5108),
        VN2CN3_sign => VN_sign_out(5109),
        VN2CN4_sign => VN_sign_out(5110),
        VN2CN5_sign => VN_sign_out(5111),
        codeword => codeword(851),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN852 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5117 downto 5112),
        Din0 => VN852_in0,
        Din1 => VN852_in1,
        Din2 => VN852_in2,
        Din3 => VN852_in3,
        Din4 => VN852_in4,
        Din5 => VN852_in5,
        VN2CN0_bit => VN_data_out(5112),
        VN2CN1_bit => VN_data_out(5113),
        VN2CN2_bit => VN_data_out(5114),
        VN2CN3_bit => VN_data_out(5115),
        VN2CN4_bit => VN_data_out(5116),
        VN2CN5_bit => VN_data_out(5117),
        VN2CN0_sign => VN_sign_out(5112),
        VN2CN1_sign => VN_sign_out(5113),
        VN2CN2_sign => VN_sign_out(5114),
        VN2CN3_sign => VN_sign_out(5115),
        VN2CN4_sign => VN_sign_out(5116),
        VN2CN5_sign => VN_sign_out(5117),
        codeword => codeword(852),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN853 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5123 downto 5118),
        Din0 => VN853_in0,
        Din1 => VN853_in1,
        Din2 => VN853_in2,
        Din3 => VN853_in3,
        Din4 => VN853_in4,
        Din5 => VN853_in5,
        VN2CN0_bit => VN_data_out(5118),
        VN2CN1_bit => VN_data_out(5119),
        VN2CN2_bit => VN_data_out(5120),
        VN2CN3_bit => VN_data_out(5121),
        VN2CN4_bit => VN_data_out(5122),
        VN2CN5_bit => VN_data_out(5123),
        VN2CN0_sign => VN_sign_out(5118),
        VN2CN1_sign => VN_sign_out(5119),
        VN2CN2_sign => VN_sign_out(5120),
        VN2CN3_sign => VN_sign_out(5121),
        VN2CN4_sign => VN_sign_out(5122),
        VN2CN5_sign => VN_sign_out(5123),
        codeword => codeword(853),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN854 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5129 downto 5124),
        Din0 => VN854_in0,
        Din1 => VN854_in1,
        Din2 => VN854_in2,
        Din3 => VN854_in3,
        Din4 => VN854_in4,
        Din5 => VN854_in5,
        VN2CN0_bit => VN_data_out(5124),
        VN2CN1_bit => VN_data_out(5125),
        VN2CN2_bit => VN_data_out(5126),
        VN2CN3_bit => VN_data_out(5127),
        VN2CN4_bit => VN_data_out(5128),
        VN2CN5_bit => VN_data_out(5129),
        VN2CN0_sign => VN_sign_out(5124),
        VN2CN1_sign => VN_sign_out(5125),
        VN2CN2_sign => VN_sign_out(5126),
        VN2CN3_sign => VN_sign_out(5127),
        VN2CN4_sign => VN_sign_out(5128),
        VN2CN5_sign => VN_sign_out(5129),
        codeword => codeword(854),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN855 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5135 downto 5130),
        Din0 => VN855_in0,
        Din1 => VN855_in1,
        Din2 => VN855_in2,
        Din3 => VN855_in3,
        Din4 => VN855_in4,
        Din5 => VN855_in5,
        VN2CN0_bit => VN_data_out(5130),
        VN2CN1_bit => VN_data_out(5131),
        VN2CN2_bit => VN_data_out(5132),
        VN2CN3_bit => VN_data_out(5133),
        VN2CN4_bit => VN_data_out(5134),
        VN2CN5_bit => VN_data_out(5135),
        VN2CN0_sign => VN_sign_out(5130),
        VN2CN1_sign => VN_sign_out(5131),
        VN2CN2_sign => VN_sign_out(5132),
        VN2CN3_sign => VN_sign_out(5133),
        VN2CN4_sign => VN_sign_out(5134),
        VN2CN5_sign => VN_sign_out(5135),
        codeword => codeword(855),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN856 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5141 downto 5136),
        Din0 => VN856_in0,
        Din1 => VN856_in1,
        Din2 => VN856_in2,
        Din3 => VN856_in3,
        Din4 => VN856_in4,
        Din5 => VN856_in5,
        VN2CN0_bit => VN_data_out(5136),
        VN2CN1_bit => VN_data_out(5137),
        VN2CN2_bit => VN_data_out(5138),
        VN2CN3_bit => VN_data_out(5139),
        VN2CN4_bit => VN_data_out(5140),
        VN2CN5_bit => VN_data_out(5141),
        VN2CN0_sign => VN_sign_out(5136),
        VN2CN1_sign => VN_sign_out(5137),
        VN2CN2_sign => VN_sign_out(5138),
        VN2CN3_sign => VN_sign_out(5139),
        VN2CN4_sign => VN_sign_out(5140),
        VN2CN5_sign => VN_sign_out(5141),
        codeword => codeword(856),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN857 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5147 downto 5142),
        Din0 => VN857_in0,
        Din1 => VN857_in1,
        Din2 => VN857_in2,
        Din3 => VN857_in3,
        Din4 => VN857_in4,
        Din5 => VN857_in5,
        VN2CN0_bit => VN_data_out(5142),
        VN2CN1_bit => VN_data_out(5143),
        VN2CN2_bit => VN_data_out(5144),
        VN2CN3_bit => VN_data_out(5145),
        VN2CN4_bit => VN_data_out(5146),
        VN2CN5_bit => VN_data_out(5147),
        VN2CN0_sign => VN_sign_out(5142),
        VN2CN1_sign => VN_sign_out(5143),
        VN2CN2_sign => VN_sign_out(5144),
        VN2CN3_sign => VN_sign_out(5145),
        VN2CN4_sign => VN_sign_out(5146),
        VN2CN5_sign => VN_sign_out(5147),
        codeword => codeword(857),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN858 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5153 downto 5148),
        Din0 => VN858_in0,
        Din1 => VN858_in1,
        Din2 => VN858_in2,
        Din3 => VN858_in3,
        Din4 => VN858_in4,
        Din5 => VN858_in5,
        VN2CN0_bit => VN_data_out(5148),
        VN2CN1_bit => VN_data_out(5149),
        VN2CN2_bit => VN_data_out(5150),
        VN2CN3_bit => VN_data_out(5151),
        VN2CN4_bit => VN_data_out(5152),
        VN2CN5_bit => VN_data_out(5153),
        VN2CN0_sign => VN_sign_out(5148),
        VN2CN1_sign => VN_sign_out(5149),
        VN2CN2_sign => VN_sign_out(5150),
        VN2CN3_sign => VN_sign_out(5151),
        VN2CN4_sign => VN_sign_out(5152),
        VN2CN5_sign => VN_sign_out(5153),
        codeword => codeword(858),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN859 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5159 downto 5154),
        Din0 => VN859_in0,
        Din1 => VN859_in1,
        Din2 => VN859_in2,
        Din3 => VN859_in3,
        Din4 => VN859_in4,
        Din5 => VN859_in5,
        VN2CN0_bit => VN_data_out(5154),
        VN2CN1_bit => VN_data_out(5155),
        VN2CN2_bit => VN_data_out(5156),
        VN2CN3_bit => VN_data_out(5157),
        VN2CN4_bit => VN_data_out(5158),
        VN2CN5_bit => VN_data_out(5159),
        VN2CN0_sign => VN_sign_out(5154),
        VN2CN1_sign => VN_sign_out(5155),
        VN2CN2_sign => VN_sign_out(5156),
        VN2CN3_sign => VN_sign_out(5157),
        VN2CN4_sign => VN_sign_out(5158),
        VN2CN5_sign => VN_sign_out(5159),
        codeword => codeword(859),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN860 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5165 downto 5160),
        Din0 => VN860_in0,
        Din1 => VN860_in1,
        Din2 => VN860_in2,
        Din3 => VN860_in3,
        Din4 => VN860_in4,
        Din5 => VN860_in5,
        VN2CN0_bit => VN_data_out(5160),
        VN2CN1_bit => VN_data_out(5161),
        VN2CN2_bit => VN_data_out(5162),
        VN2CN3_bit => VN_data_out(5163),
        VN2CN4_bit => VN_data_out(5164),
        VN2CN5_bit => VN_data_out(5165),
        VN2CN0_sign => VN_sign_out(5160),
        VN2CN1_sign => VN_sign_out(5161),
        VN2CN2_sign => VN_sign_out(5162),
        VN2CN3_sign => VN_sign_out(5163),
        VN2CN4_sign => VN_sign_out(5164),
        VN2CN5_sign => VN_sign_out(5165),
        codeword => codeword(860),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN861 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5171 downto 5166),
        Din0 => VN861_in0,
        Din1 => VN861_in1,
        Din2 => VN861_in2,
        Din3 => VN861_in3,
        Din4 => VN861_in4,
        Din5 => VN861_in5,
        VN2CN0_bit => VN_data_out(5166),
        VN2CN1_bit => VN_data_out(5167),
        VN2CN2_bit => VN_data_out(5168),
        VN2CN3_bit => VN_data_out(5169),
        VN2CN4_bit => VN_data_out(5170),
        VN2CN5_bit => VN_data_out(5171),
        VN2CN0_sign => VN_sign_out(5166),
        VN2CN1_sign => VN_sign_out(5167),
        VN2CN2_sign => VN_sign_out(5168),
        VN2CN3_sign => VN_sign_out(5169),
        VN2CN4_sign => VN_sign_out(5170),
        VN2CN5_sign => VN_sign_out(5171),
        codeword => codeword(861),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN862 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5177 downto 5172),
        Din0 => VN862_in0,
        Din1 => VN862_in1,
        Din2 => VN862_in2,
        Din3 => VN862_in3,
        Din4 => VN862_in4,
        Din5 => VN862_in5,
        VN2CN0_bit => VN_data_out(5172),
        VN2CN1_bit => VN_data_out(5173),
        VN2CN2_bit => VN_data_out(5174),
        VN2CN3_bit => VN_data_out(5175),
        VN2CN4_bit => VN_data_out(5176),
        VN2CN5_bit => VN_data_out(5177),
        VN2CN0_sign => VN_sign_out(5172),
        VN2CN1_sign => VN_sign_out(5173),
        VN2CN2_sign => VN_sign_out(5174),
        VN2CN3_sign => VN_sign_out(5175),
        VN2CN4_sign => VN_sign_out(5176),
        VN2CN5_sign => VN_sign_out(5177),
        codeword => codeword(862),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN863 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5183 downto 5178),
        Din0 => VN863_in0,
        Din1 => VN863_in1,
        Din2 => VN863_in2,
        Din3 => VN863_in3,
        Din4 => VN863_in4,
        Din5 => VN863_in5,
        VN2CN0_bit => VN_data_out(5178),
        VN2CN1_bit => VN_data_out(5179),
        VN2CN2_bit => VN_data_out(5180),
        VN2CN3_bit => VN_data_out(5181),
        VN2CN4_bit => VN_data_out(5182),
        VN2CN5_bit => VN_data_out(5183),
        VN2CN0_sign => VN_sign_out(5178),
        VN2CN1_sign => VN_sign_out(5179),
        VN2CN2_sign => VN_sign_out(5180),
        VN2CN3_sign => VN_sign_out(5181),
        VN2CN4_sign => VN_sign_out(5182),
        VN2CN5_sign => VN_sign_out(5183),
        codeword => codeword(863),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN864 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5189 downto 5184),
        Din0 => VN864_in0,
        Din1 => VN864_in1,
        Din2 => VN864_in2,
        Din3 => VN864_in3,
        Din4 => VN864_in4,
        Din5 => VN864_in5,
        VN2CN0_bit => VN_data_out(5184),
        VN2CN1_bit => VN_data_out(5185),
        VN2CN2_bit => VN_data_out(5186),
        VN2CN3_bit => VN_data_out(5187),
        VN2CN4_bit => VN_data_out(5188),
        VN2CN5_bit => VN_data_out(5189),
        VN2CN0_sign => VN_sign_out(5184),
        VN2CN1_sign => VN_sign_out(5185),
        VN2CN2_sign => VN_sign_out(5186),
        VN2CN3_sign => VN_sign_out(5187),
        VN2CN4_sign => VN_sign_out(5188),
        VN2CN5_sign => VN_sign_out(5189),
        codeword => codeword(864),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN865 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5195 downto 5190),
        Din0 => VN865_in0,
        Din1 => VN865_in1,
        Din2 => VN865_in2,
        Din3 => VN865_in3,
        Din4 => VN865_in4,
        Din5 => VN865_in5,
        VN2CN0_bit => VN_data_out(5190),
        VN2CN1_bit => VN_data_out(5191),
        VN2CN2_bit => VN_data_out(5192),
        VN2CN3_bit => VN_data_out(5193),
        VN2CN4_bit => VN_data_out(5194),
        VN2CN5_bit => VN_data_out(5195),
        VN2CN0_sign => VN_sign_out(5190),
        VN2CN1_sign => VN_sign_out(5191),
        VN2CN2_sign => VN_sign_out(5192),
        VN2CN3_sign => VN_sign_out(5193),
        VN2CN4_sign => VN_sign_out(5194),
        VN2CN5_sign => VN_sign_out(5195),
        codeword => codeword(865),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN866 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5201 downto 5196),
        Din0 => VN866_in0,
        Din1 => VN866_in1,
        Din2 => VN866_in2,
        Din3 => VN866_in3,
        Din4 => VN866_in4,
        Din5 => VN866_in5,
        VN2CN0_bit => VN_data_out(5196),
        VN2CN1_bit => VN_data_out(5197),
        VN2CN2_bit => VN_data_out(5198),
        VN2CN3_bit => VN_data_out(5199),
        VN2CN4_bit => VN_data_out(5200),
        VN2CN5_bit => VN_data_out(5201),
        VN2CN0_sign => VN_sign_out(5196),
        VN2CN1_sign => VN_sign_out(5197),
        VN2CN2_sign => VN_sign_out(5198),
        VN2CN3_sign => VN_sign_out(5199),
        VN2CN4_sign => VN_sign_out(5200),
        VN2CN5_sign => VN_sign_out(5201),
        codeword => codeword(866),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN867 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5207 downto 5202),
        Din0 => VN867_in0,
        Din1 => VN867_in1,
        Din2 => VN867_in2,
        Din3 => VN867_in3,
        Din4 => VN867_in4,
        Din5 => VN867_in5,
        VN2CN0_bit => VN_data_out(5202),
        VN2CN1_bit => VN_data_out(5203),
        VN2CN2_bit => VN_data_out(5204),
        VN2CN3_bit => VN_data_out(5205),
        VN2CN4_bit => VN_data_out(5206),
        VN2CN5_bit => VN_data_out(5207),
        VN2CN0_sign => VN_sign_out(5202),
        VN2CN1_sign => VN_sign_out(5203),
        VN2CN2_sign => VN_sign_out(5204),
        VN2CN3_sign => VN_sign_out(5205),
        VN2CN4_sign => VN_sign_out(5206),
        VN2CN5_sign => VN_sign_out(5207),
        codeword => codeword(867),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN868 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5213 downto 5208),
        Din0 => VN868_in0,
        Din1 => VN868_in1,
        Din2 => VN868_in2,
        Din3 => VN868_in3,
        Din4 => VN868_in4,
        Din5 => VN868_in5,
        VN2CN0_bit => VN_data_out(5208),
        VN2CN1_bit => VN_data_out(5209),
        VN2CN2_bit => VN_data_out(5210),
        VN2CN3_bit => VN_data_out(5211),
        VN2CN4_bit => VN_data_out(5212),
        VN2CN5_bit => VN_data_out(5213),
        VN2CN0_sign => VN_sign_out(5208),
        VN2CN1_sign => VN_sign_out(5209),
        VN2CN2_sign => VN_sign_out(5210),
        VN2CN3_sign => VN_sign_out(5211),
        VN2CN4_sign => VN_sign_out(5212),
        VN2CN5_sign => VN_sign_out(5213),
        codeword => codeword(868),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN869 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5219 downto 5214),
        Din0 => VN869_in0,
        Din1 => VN869_in1,
        Din2 => VN869_in2,
        Din3 => VN869_in3,
        Din4 => VN869_in4,
        Din5 => VN869_in5,
        VN2CN0_bit => VN_data_out(5214),
        VN2CN1_bit => VN_data_out(5215),
        VN2CN2_bit => VN_data_out(5216),
        VN2CN3_bit => VN_data_out(5217),
        VN2CN4_bit => VN_data_out(5218),
        VN2CN5_bit => VN_data_out(5219),
        VN2CN0_sign => VN_sign_out(5214),
        VN2CN1_sign => VN_sign_out(5215),
        VN2CN2_sign => VN_sign_out(5216),
        VN2CN3_sign => VN_sign_out(5217),
        VN2CN4_sign => VN_sign_out(5218),
        VN2CN5_sign => VN_sign_out(5219),
        codeword => codeword(869),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN870 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5225 downto 5220),
        Din0 => VN870_in0,
        Din1 => VN870_in1,
        Din2 => VN870_in2,
        Din3 => VN870_in3,
        Din4 => VN870_in4,
        Din5 => VN870_in5,
        VN2CN0_bit => VN_data_out(5220),
        VN2CN1_bit => VN_data_out(5221),
        VN2CN2_bit => VN_data_out(5222),
        VN2CN3_bit => VN_data_out(5223),
        VN2CN4_bit => VN_data_out(5224),
        VN2CN5_bit => VN_data_out(5225),
        VN2CN0_sign => VN_sign_out(5220),
        VN2CN1_sign => VN_sign_out(5221),
        VN2CN2_sign => VN_sign_out(5222),
        VN2CN3_sign => VN_sign_out(5223),
        VN2CN4_sign => VN_sign_out(5224),
        VN2CN5_sign => VN_sign_out(5225),
        codeword => codeword(870),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN871 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5231 downto 5226),
        Din0 => VN871_in0,
        Din1 => VN871_in1,
        Din2 => VN871_in2,
        Din3 => VN871_in3,
        Din4 => VN871_in4,
        Din5 => VN871_in5,
        VN2CN0_bit => VN_data_out(5226),
        VN2CN1_bit => VN_data_out(5227),
        VN2CN2_bit => VN_data_out(5228),
        VN2CN3_bit => VN_data_out(5229),
        VN2CN4_bit => VN_data_out(5230),
        VN2CN5_bit => VN_data_out(5231),
        VN2CN0_sign => VN_sign_out(5226),
        VN2CN1_sign => VN_sign_out(5227),
        VN2CN2_sign => VN_sign_out(5228),
        VN2CN3_sign => VN_sign_out(5229),
        VN2CN4_sign => VN_sign_out(5230),
        VN2CN5_sign => VN_sign_out(5231),
        codeword => codeword(871),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN872 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5237 downto 5232),
        Din0 => VN872_in0,
        Din1 => VN872_in1,
        Din2 => VN872_in2,
        Din3 => VN872_in3,
        Din4 => VN872_in4,
        Din5 => VN872_in5,
        VN2CN0_bit => VN_data_out(5232),
        VN2CN1_bit => VN_data_out(5233),
        VN2CN2_bit => VN_data_out(5234),
        VN2CN3_bit => VN_data_out(5235),
        VN2CN4_bit => VN_data_out(5236),
        VN2CN5_bit => VN_data_out(5237),
        VN2CN0_sign => VN_sign_out(5232),
        VN2CN1_sign => VN_sign_out(5233),
        VN2CN2_sign => VN_sign_out(5234),
        VN2CN3_sign => VN_sign_out(5235),
        VN2CN4_sign => VN_sign_out(5236),
        VN2CN5_sign => VN_sign_out(5237),
        codeword => codeword(872),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN873 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5243 downto 5238),
        Din0 => VN873_in0,
        Din1 => VN873_in1,
        Din2 => VN873_in2,
        Din3 => VN873_in3,
        Din4 => VN873_in4,
        Din5 => VN873_in5,
        VN2CN0_bit => VN_data_out(5238),
        VN2CN1_bit => VN_data_out(5239),
        VN2CN2_bit => VN_data_out(5240),
        VN2CN3_bit => VN_data_out(5241),
        VN2CN4_bit => VN_data_out(5242),
        VN2CN5_bit => VN_data_out(5243),
        VN2CN0_sign => VN_sign_out(5238),
        VN2CN1_sign => VN_sign_out(5239),
        VN2CN2_sign => VN_sign_out(5240),
        VN2CN3_sign => VN_sign_out(5241),
        VN2CN4_sign => VN_sign_out(5242),
        VN2CN5_sign => VN_sign_out(5243),
        codeword => codeword(873),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN874 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5249 downto 5244),
        Din0 => VN874_in0,
        Din1 => VN874_in1,
        Din2 => VN874_in2,
        Din3 => VN874_in3,
        Din4 => VN874_in4,
        Din5 => VN874_in5,
        VN2CN0_bit => VN_data_out(5244),
        VN2CN1_bit => VN_data_out(5245),
        VN2CN2_bit => VN_data_out(5246),
        VN2CN3_bit => VN_data_out(5247),
        VN2CN4_bit => VN_data_out(5248),
        VN2CN5_bit => VN_data_out(5249),
        VN2CN0_sign => VN_sign_out(5244),
        VN2CN1_sign => VN_sign_out(5245),
        VN2CN2_sign => VN_sign_out(5246),
        VN2CN3_sign => VN_sign_out(5247),
        VN2CN4_sign => VN_sign_out(5248),
        VN2CN5_sign => VN_sign_out(5249),
        codeword => codeword(874),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN875 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5255 downto 5250),
        Din0 => VN875_in0,
        Din1 => VN875_in1,
        Din2 => VN875_in2,
        Din3 => VN875_in3,
        Din4 => VN875_in4,
        Din5 => VN875_in5,
        VN2CN0_bit => VN_data_out(5250),
        VN2CN1_bit => VN_data_out(5251),
        VN2CN2_bit => VN_data_out(5252),
        VN2CN3_bit => VN_data_out(5253),
        VN2CN4_bit => VN_data_out(5254),
        VN2CN5_bit => VN_data_out(5255),
        VN2CN0_sign => VN_sign_out(5250),
        VN2CN1_sign => VN_sign_out(5251),
        VN2CN2_sign => VN_sign_out(5252),
        VN2CN3_sign => VN_sign_out(5253),
        VN2CN4_sign => VN_sign_out(5254),
        VN2CN5_sign => VN_sign_out(5255),
        codeword => codeword(875),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN876 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5261 downto 5256),
        Din0 => VN876_in0,
        Din1 => VN876_in1,
        Din2 => VN876_in2,
        Din3 => VN876_in3,
        Din4 => VN876_in4,
        Din5 => VN876_in5,
        VN2CN0_bit => VN_data_out(5256),
        VN2CN1_bit => VN_data_out(5257),
        VN2CN2_bit => VN_data_out(5258),
        VN2CN3_bit => VN_data_out(5259),
        VN2CN4_bit => VN_data_out(5260),
        VN2CN5_bit => VN_data_out(5261),
        VN2CN0_sign => VN_sign_out(5256),
        VN2CN1_sign => VN_sign_out(5257),
        VN2CN2_sign => VN_sign_out(5258),
        VN2CN3_sign => VN_sign_out(5259),
        VN2CN4_sign => VN_sign_out(5260),
        VN2CN5_sign => VN_sign_out(5261),
        codeword => codeword(876),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN877 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5267 downto 5262),
        Din0 => VN877_in0,
        Din1 => VN877_in1,
        Din2 => VN877_in2,
        Din3 => VN877_in3,
        Din4 => VN877_in4,
        Din5 => VN877_in5,
        VN2CN0_bit => VN_data_out(5262),
        VN2CN1_bit => VN_data_out(5263),
        VN2CN2_bit => VN_data_out(5264),
        VN2CN3_bit => VN_data_out(5265),
        VN2CN4_bit => VN_data_out(5266),
        VN2CN5_bit => VN_data_out(5267),
        VN2CN0_sign => VN_sign_out(5262),
        VN2CN1_sign => VN_sign_out(5263),
        VN2CN2_sign => VN_sign_out(5264),
        VN2CN3_sign => VN_sign_out(5265),
        VN2CN4_sign => VN_sign_out(5266),
        VN2CN5_sign => VN_sign_out(5267),
        codeword => codeword(877),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN878 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5273 downto 5268),
        Din0 => VN878_in0,
        Din1 => VN878_in1,
        Din2 => VN878_in2,
        Din3 => VN878_in3,
        Din4 => VN878_in4,
        Din5 => VN878_in5,
        VN2CN0_bit => VN_data_out(5268),
        VN2CN1_bit => VN_data_out(5269),
        VN2CN2_bit => VN_data_out(5270),
        VN2CN3_bit => VN_data_out(5271),
        VN2CN4_bit => VN_data_out(5272),
        VN2CN5_bit => VN_data_out(5273),
        VN2CN0_sign => VN_sign_out(5268),
        VN2CN1_sign => VN_sign_out(5269),
        VN2CN2_sign => VN_sign_out(5270),
        VN2CN3_sign => VN_sign_out(5271),
        VN2CN4_sign => VN_sign_out(5272),
        VN2CN5_sign => VN_sign_out(5273),
        codeword => codeword(878),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN879 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5279 downto 5274),
        Din0 => VN879_in0,
        Din1 => VN879_in1,
        Din2 => VN879_in2,
        Din3 => VN879_in3,
        Din4 => VN879_in4,
        Din5 => VN879_in5,
        VN2CN0_bit => VN_data_out(5274),
        VN2CN1_bit => VN_data_out(5275),
        VN2CN2_bit => VN_data_out(5276),
        VN2CN3_bit => VN_data_out(5277),
        VN2CN4_bit => VN_data_out(5278),
        VN2CN5_bit => VN_data_out(5279),
        VN2CN0_sign => VN_sign_out(5274),
        VN2CN1_sign => VN_sign_out(5275),
        VN2CN2_sign => VN_sign_out(5276),
        VN2CN3_sign => VN_sign_out(5277),
        VN2CN4_sign => VN_sign_out(5278),
        VN2CN5_sign => VN_sign_out(5279),
        codeword => codeword(879),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN880 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5285 downto 5280),
        Din0 => VN880_in0,
        Din1 => VN880_in1,
        Din2 => VN880_in2,
        Din3 => VN880_in3,
        Din4 => VN880_in4,
        Din5 => VN880_in5,
        VN2CN0_bit => VN_data_out(5280),
        VN2CN1_bit => VN_data_out(5281),
        VN2CN2_bit => VN_data_out(5282),
        VN2CN3_bit => VN_data_out(5283),
        VN2CN4_bit => VN_data_out(5284),
        VN2CN5_bit => VN_data_out(5285),
        VN2CN0_sign => VN_sign_out(5280),
        VN2CN1_sign => VN_sign_out(5281),
        VN2CN2_sign => VN_sign_out(5282),
        VN2CN3_sign => VN_sign_out(5283),
        VN2CN4_sign => VN_sign_out(5284),
        VN2CN5_sign => VN_sign_out(5285),
        codeword => codeword(880),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN881 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5291 downto 5286),
        Din0 => VN881_in0,
        Din1 => VN881_in1,
        Din2 => VN881_in2,
        Din3 => VN881_in3,
        Din4 => VN881_in4,
        Din5 => VN881_in5,
        VN2CN0_bit => VN_data_out(5286),
        VN2CN1_bit => VN_data_out(5287),
        VN2CN2_bit => VN_data_out(5288),
        VN2CN3_bit => VN_data_out(5289),
        VN2CN4_bit => VN_data_out(5290),
        VN2CN5_bit => VN_data_out(5291),
        VN2CN0_sign => VN_sign_out(5286),
        VN2CN1_sign => VN_sign_out(5287),
        VN2CN2_sign => VN_sign_out(5288),
        VN2CN3_sign => VN_sign_out(5289),
        VN2CN4_sign => VN_sign_out(5290),
        VN2CN5_sign => VN_sign_out(5291),
        codeword => codeword(881),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN882 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5297 downto 5292),
        Din0 => VN882_in0,
        Din1 => VN882_in1,
        Din2 => VN882_in2,
        Din3 => VN882_in3,
        Din4 => VN882_in4,
        Din5 => VN882_in5,
        VN2CN0_bit => VN_data_out(5292),
        VN2CN1_bit => VN_data_out(5293),
        VN2CN2_bit => VN_data_out(5294),
        VN2CN3_bit => VN_data_out(5295),
        VN2CN4_bit => VN_data_out(5296),
        VN2CN5_bit => VN_data_out(5297),
        VN2CN0_sign => VN_sign_out(5292),
        VN2CN1_sign => VN_sign_out(5293),
        VN2CN2_sign => VN_sign_out(5294),
        VN2CN3_sign => VN_sign_out(5295),
        VN2CN4_sign => VN_sign_out(5296),
        VN2CN5_sign => VN_sign_out(5297),
        codeword => codeword(882),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN883 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5303 downto 5298),
        Din0 => VN883_in0,
        Din1 => VN883_in1,
        Din2 => VN883_in2,
        Din3 => VN883_in3,
        Din4 => VN883_in4,
        Din5 => VN883_in5,
        VN2CN0_bit => VN_data_out(5298),
        VN2CN1_bit => VN_data_out(5299),
        VN2CN2_bit => VN_data_out(5300),
        VN2CN3_bit => VN_data_out(5301),
        VN2CN4_bit => VN_data_out(5302),
        VN2CN5_bit => VN_data_out(5303),
        VN2CN0_sign => VN_sign_out(5298),
        VN2CN1_sign => VN_sign_out(5299),
        VN2CN2_sign => VN_sign_out(5300),
        VN2CN3_sign => VN_sign_out(5301),
        VN2CN4_sign => VN_sign_out(5302),
        VN2CN5_sign => VN_sign_out(5303),
        codeword => codeword(883),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN884 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5309 downto 5304),
        Din0 => VN884_in0,
        Din1 => VN884_in1,
        Din2 => VN884_in2,
        Din3 => VN884_in3,
        Din4 => VN884_in4,
        Din5 => VN884_in5,
        VN2CN0_bit => VN_data_out(5304),
        VN2CN1_bit => VN_data_out(5305),
        VN2CN2_bit => VN_data_out(5306),
        VN2CN3_bit => VN_data_out(5307),
        VN2CN4_bit => VN_data_out(5308),
        VN2CN5_bit => VN_data_out(5309),
        VN2CN0_sign => VN_sign_out(5304),
        VN2CN1_sign => VN_sign_out(5305),
        VN2CN2_sign => VN_sign_out(5306),
        VN2CN3_sign => VN_sign_out(5307),
        VN2CN4_sign => VN_sign_out(5308),
        VN2CN5_sign => VN_sign_out(5309),
        codeword => codeword(884),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN885 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5315 downto 5310),
        Din0 => VN885_in0,
        Din1 => VN885_in1,
        Din2 => VN885_in2,
        Din3 => VN885_in3,
        Din4 => VN885_in4,
        Din5 => VN885_in5,
        VN2CN0_bit => VN_data_out(5310),
        VN2CN1_bit => VN_data_out(5311),
        VN2CN2_bit => VN_data_out(5312),
        VN2CN3_bit => VN_data_out(5313),
        VN2CN4_bit => VN_data_out(5314),
        VN2CN5_bit => VN_data_out(5315),
        VN2CN0_sign => VN_sign_out(5310),
        VN2CN1_sign => VN_sign_out(5311),
        VN2CN2_sign => VN_sign_out(5312),
        VN2CN3_sign => VN_sign_out(5313),
        VN2CN4_sign => VN_sign_out(5314),
        VN2CN5_sign => VN_sign_out(5315),
        codeword => codeword(885),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN886 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5321 downto 5316),
        Din0 => VN886_in0,
        Din1 => VN886_in1,
        Din2 => VN886_in2,
        Din3 => VN886_in3,
        Din4 => VN886_in4,
        Din5 => VN886_in5,
        VN2CN0_bit => VN_data_out(5316),
        VN2CN1_bit => VN_data_out(5317),
        VN2CN2_bit => VN_data_out(5318),
        VN2CN3_bit => VN_data_out(5319),
        VN2CN4_bit => VN_data_out(5320),
        VN2CN5_bit => VN_data_out(5321),
        VN2CN0_sign => VN_sign_out(5316),
        VN2CN1_sign => VN_sign_out(5317),
        VN2CN2_sign => VN_sign_out(5318),
        VN2CN3_sign => VN_sign_out(5319),
        VN2CN4_sign => VN_sign_out(5320),
        VN2CN5_sign => VN_sign_out(5321),
        codeword => codeword(886),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN887 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5327 downto 5322),
        Din0 => VN887_in0,
        Din1 => VN887_in1,
        Din2 => VN887_in2,
        Din3 => VN887_in3,
        Din4 => VN887_in4,
        Din5 => VN887_in5,
        VN2CN0_bit => VN_data_out(5322),
        VN2CN1_bit => VN_data_out(5323),
        VN2CN2_bit => VN_data_out(5324),
        VN2CN3_bit => VN_data_out(5325),
        VN2CN4_bit => VN_data_out(5326),
        VN2CN5_bit => VN_data_out(5327),
        VN2CN0_sign => VN_sign_out(5322),
        VN2CN1_sign => VN_sign_out(5323),
        VN2CN2_sign => VN_sign_out(5324),
        VN2CN3_sign => VN_sign_out(5325),
        VN2CN4_sign => VN_sign_out(5326),
        VN2CN5_sign => VN_sign_out(5327),
        codeword => codeword(887),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN888 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5333 downto 5328),
        Din0 => VN888_in0,
        Din1 => VN888_in1,
        Din2 => VN888_in2,
        Din3 => VN888_in3,
        Din4 => VN888_in4,
        Din5 => VN888_in5,
        VN2CN0_bit => VN_data_out(5328),
        VN2CN1_bit => VN_data_out(5329),
        VN2CN2_bit => VN_data_out(5330),
        VN2CN3_bit => VN_data_out(5331),
        VN2CN4_bit => VN_data_out(5332),
        VN2CN5_bit => VN_data_out(5333),
        VN2CN0_sign => VN_sign_out(5328),
        VN2CN1_sign => VN_sign_out(5329),
        VN2CN2_sign => VN_sign_out(5330),
        VN2CN3_sign => VN_sign_out(5331),
        VN2CN4_sign => VN_sign_out(5332),
        VN2CN5_sign => VN_sign_out(5333),
        codeword => codeword(888),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN889 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5339 downto 5334),
        Din0 => VN889_in0,
        Din1 => VN889_in1,
        Din2 => VN889_in2,
        Din3 => VN889_in3,
        Din4 => VN889_in4,
        Din5 => VN889_in5,
        VN2CN0_bit => VN_data_out(5334),
        VN2CN1_bit => VN_data_out(5335),
        VN2CN2_bit => VN_data_out(5336),
        VN2CN3_bit => VN_data_out(5337),
        VN2CN4_bit => VN_data_out(5338),
        VN2CN5_bit => VN_data_out(5339),
        VN2CN0_sign => VN_sign_out(5334),
        VN2CN1_sign => VN_sign_out(5335),
        VN2CN2_sign => VN_sign_out(5336),
        VN2CN3_sign => VN_sign_out(5337),
        VN2CN4_sign => VN_sign_out(5338),
        VN2CN5_sign => VN_sign_out(5339),
        codeword => codeword(889),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN890 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5345 downto 5340),
        Din0 => VN890_in0,
        Din1 => VN890_in1,
        Din2 => VN890_in2,
        Din3 => VN890_in3,
        Din4 => VN890_in4,
        Din5 => VN890_in5,
        VN2CN0_bit => VN_data_out(5340),
        VN2CN1_bit => VN_data_out(5341),
        VN2CN2_bit => VN_data_out(5342),
        VN2CN3_bit => VN_data_out(5343),
        VN2CN4_bit => VN_data_out(5344),
        VN2CN5_bit => VN_data_out(5345),
        VN2CN0_sign => VN_sign_out(5340),
        VN2CN1_sign => VN_sign_out(5341),
        VN2CN2_sign => VN_sign_out(5342),
        VN2CN3_sign => VN_sign_out(5343),
        VN2CN4_sign => VN_sign_out(5344),
        VN2CN5_sign => VN_sign_out(5345),
        codeword => codeword(890),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN891 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5351 downto 5346),
        Din0 => VN891_in0,
        Din1 => VN891_in1,
        Din2 => VN891_in2,
        Din3 => VN891_in3,
        Din4 => VN891_in4,
        Din5 => VN891_in5,
        VN2CN0_bit => VN_data_out(5346),
        VN2CN1_bit => VN_data_out(5347),
        VN2CN2_bit => VN_data_out(5348),
        VN2CN3_bit => VN_data_out(5349),
        VN2CN4_bit => VN_data_out(5350),
        VN2CN5_bit => VN_data_out(5351),
        VN2CN0_sign => VN_sign_out(5346),
        VN2CN1_sign => VN_sign_out(5347),
        VN2CN2_sign => VN_sign_out(5348),
        VN2CN3_sign => VN_sign_out(5349),
        VN2CN4_sign => VN_sign_out(5350),
        VN2CN5_sign => VN_sign_out(5351),
        codeword => codeword(891),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN892 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5357 downto 5352),
        Din0 => VN892_in0,
        Din1 => VN892_in1,
        Din2 => VN892_in2,
        Din3 => VN892_in3,
        Din4 => VN892_in4,
        Din5 => VN892_in5,
        VN2CN0_bit => VN_data_out(5352),
        VN2CN1_bit => VN_data_out(5353),
        VN2CN2_bit => VN_data_out(5354),
        VN2CN3_bit => VN_data_out(5355),
        VN2CN4_bit => VN_data_out(5356),
        VN2CN5_bit => VN_data_out(5357),
        VN2CN0_sign => VN_sign_out(5352),
        VN2CN1_sign => VN_sign_out(5353),
        VN2CN2_sign => VN_sign_out(5354),
        VN2CN3_sign => VN_sign_out(5355),
        VN2CN4_sign => VN_sign_out(5356),
        VN2CN5_sign => VN_sign_out(5357),
        codeword => codeword(892),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN893 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5363 downto 5358),
        Din0 => VN893_in0,
        Din1 => VN893_in1,
        Din2 => VN893_in2,
        Din3 => VN893_in3,
        Din4 => VN893_in4,
        Din5 => VN893_in5,
        VN2CN0_bit => VN_data_out(5358),
        VN2CN1_bit => VN_data_out(5359),
        VN2CN2_bit => VN_data_out(5360),
        VN2CN3_bit => VN_data_out(5361),
        VN2CN4_bit => VN_data_out(5362),
        VN2CN5_bit => VN_data_out(5363),
        VN2CN0_sign => VN_sign_out(5358),
        VN2CN1_sign => VN_sign_out(5359),
        VN2CN2_sign => VN_sign_out(5360),
        VN2CN3_sign => VN_sign_out(5361),
        VN2CN4_sign => VN_sign_out(5362),
        VN2CN5_sign => VN_sign_out(5363),
        codeword => codeword(893),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN894 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5369 downto 5364),
        Din0 => VN894_in0,
        Din1 => VN894_in1,
        Din2 => VN894_in2,
        Din3 => VN894_in3,
        Din4 => VN894_in4,
        Din5 => VN894_in5,
        VN2CN0_bit => VN_data_out(5364),
        VN2CN1_bit => VN_data_out(5365),
        VN2CN2_bit => VN_data_out(5366),
        VN2CN3_bit => VN_data_out(5367),
        VN2CN4_bit => VN_data_out(5368),
        VN2CN5_bit => VN_data_out(5369),
        VN2CN0_sign => VN_sign_out(5364),
        VN2CN1_sign => VN_sign_out(5365),
        VN2CN2_sign => VN_sign_out(5366),
        VN2CN3_sign => VN_sign_out(5367),
        VN2CN4_sign => VN_sign_out(5368),
        VN2CN5_sign => VN_sign_out(5369),
        codeword => codeword(894),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN895 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5375 downto 5370),
        Din0 => VN895_in0,
        Din1 => VN895_in1,
        Din2 => VN895_in2,
        Din3 => VN895_in3,
        Din4 => VN895_in4,
        Din5 => VN895_in5,
        VN2CN0_bit => VN_data_out(5370),
        VN2CN1_bit => VN_data_out(5371),
        VN2CN2_bit => VN_data_out(5372),
        VN2CN3_bit => VN_data_out(5373),
        VN2CN4_bit => VN_data_out(5374),
        VN2CN5_bit => VN_data_out(5375),
        VN2CN0_sign => VN_sign_out(5370),
        VN2CN1_sign => VN_sign_out(5371),
        VN2CN2_sign => VN_sign_out(5372),
        VN2CN3_sign => VN_sign_out(5373),
        VN2CN4_sign => VN_sign_out(5374),
        VN2CN5_sign => VN_sign_out(5375),
        codeword => codeword(895),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN896 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5381 downto 5376),
        Din0 => VN896_in0,
        Din1 => VN896_in1,
        Din2 => VN896_in2,
        Din3 => VN896_in3,
        Din4 => VN896_in4,
        Din5 => VN896_in5,
        VN2CN0_bit => VN_data_out(5376),
        VN2CN1_bit => VN_data_out(5377),
        VN2CN2_bit => VN_data_out(5378),
        VN2CN3_bit => VN_data_out(5379),
        VN2CN4_bit => VN_data_out(5380),
        VN2CN5_bit => VN_data_out(5381),
        VN2CN0_sign => VN_sign_out(5376),
        VN2CN1_sign => VN_sign_out(5377),
        VN2CN2_sign => VN_sign_out(5378),
        VN2CN3_sign => VN_sign_out(5379),
        VN2CN4_sign => VN_sign_out(5380),
        VN2CN5_sign => VN_sign_out(5381),
        codeword => codeword(896),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN897 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5387 downto 5382),
        Din0 => VN897_in0,
        Din1 => VN897_in1,
        Din2 => VN897_in2,
        Din3 => VN897_in3,
        Din4 => VN897_in4,
        Din5 => VN897_in5,
        VN2CN0_bit => VN_data_out(5382),
        VN2CN1_bit => VN_data_out(5383),
        VN2CN2_bit => VN_data_out(5384),
        VN2CN3_bit => VN_data_out(5385),
        VN2CN4_bit => VN_data_out(5386),
        VN2CN5_bit => VN_data_out(5387),
        VN2CN0_sign => VN_sign_out(5382),
        VN2CN1_sign => VN_sign_out(5383),
        VN2CN2_sign => VN_sign_out(5384),
        VN2CN3_sign => VN_sign_out(5385),
        VN2CN4_sign => VN_sign_out(5386),
        VN2CN5_sign => VN_sign_out(5387),
        codeword => codeword(897),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN898 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5393 downto 5388),
        Din0 => VN898_in0,
        Din1 => VN898_in1,
        Din2 => VN898_in2,
        Din3 => VN898_in3,
        Din4 => VN898_in4,
        Din5 => VN898_in5,
        VN2CN0_bit => VN_data_out(5388),
        VN2CN1_bit => VN_data_out(5389),
        VN2CN2_bit => VN_data_out(5390),
        VN2CN3_bit => VN_data_out(5391),
        VN2CN4_bit => VN_data_out(5392),
        VN2CN5_bit => VN_data_out(5393),
        VN2CN0_sign => VN_sign_out(5388),
        VN2CN1_sign => VN_sign_out(5389),
        VN2CN2_sign => VN_sign_out(5390),
        VN2CN3_sign => VN_sign_out(5391),
        VN2CN4_sign => VN_sign_out(5392),
        VN2CN5_sign => VN_sign_out(5393),
        codeword => codeword(898),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN899 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5399 downto 5394),
        Din0 => VN899_in0,
        Din1 => VN899_in1,
        Din2 => VN899_in2,
        Din3 => VN899_in3,
        Din4 => VN899_in4,
        Din5 => VN899_in5,
        VN2CN0_bit => VN_data_out(5394),
        VN2CN1_bit => VN_data_out(5395),
        VN2CN2_bit => VN_data_out(5396),
        VN2CN3_bit => VN_data_out(5397),
        VN2CN4_bit => VN_data_out(5398),
        VN2CN5_bit => VN_data_out(5399),
        VN2CN0_sign => VN_sign_out(5394),
        VN2CN1_sign => VN_sign_out(5395),
        VN2CN2_sign => VN_sign_out(5396),
        VN2CN3_sign => VN_sign_out(5397),
        VN2CN4_sign => VN_sign_out(5398),
        VN2CN5_sign => VN_sign_out(5399),
        codeword => codeword(899),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN900 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5405 downto 5400),
        Din0 => VN900_in0,
        Din1 => VN900_in1,
        Din2 => VN900_in2,
        Din3 => VN900_in3,
        Din4 => VN900_in4,
        Din5 => VN900_in5,
        VN2CN0_bit => VN_data_out(5400),
        VN2CN1_bit => VN_data_out(5401),
        VN2CN2_bit => VN_data_out(5402),
        VN2CN3_bit => VN_data_out(5403),
        VN2CN4_bit => VN_data_out(5404),
        VN2CN5_bit => VN_data_out(5405),
        VN2CN0_sign => VN_sign_out(5400),
        VN2CN1_sign => VN_sign_out(5401),
        VN2CN2_sign => VN_sign_out(5402),
        VN2CN3_sign => VN_sign_out(5403),
        VN2CN4_sign => VN_sign_out(5404),
        VN2CN5_sign => VN_sign_out(5405),
        codeword => codeword(900),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN901 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5411 downto 5406),
        Din0 => VN901_in0,
        Din1 => VN901_in1,
        Din2 => VN901_in2,
        Din3 => VN901_in3,
        Din4 => VN901_in4,
        Din5 => VN901_in5,
        VN2CN0_bit => VN_data_out(5406),
        VN2CN1_bit => VN_data_out(5407),
        VN2CN2_bit => VN_data_out(5408),
        VN2CN3_bit => VN_data_out(5409),
        VN2CN4_bit => VN_data_out(5410),
        VN2CN5_bit => VN_data_out(5411),
        VN2CN0_sign => VN_sign_out(5406),
        VN2CN1_sign => VN_sign_out(5407),
        VN2CN2_sign => VN_sign_out(5408),
        VN2CN3_sign => VN_sign_out(5409),
        VN2CN4_sign => VN_sign_out(5410),
        VN2CN5_sign => VN_sign_out(5411),
        codeword => codeword(901),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN902 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5417 downto 5412),
        Din0 => VN902_in0,
        Din1 => VN902_in1,
        Din2 => VN902_in2,
        Din3 => VN902_in3,
        Din4 => VN902_in4,
        Din5 => VN902_in5,
        VN2CN0_bit => VN_data_out(5412),
        VN2CN1_bit => VN_data_out(5413),
        VN2CN2_bit => VN_data_out(5414),
        VN2CN3_bit => VN_data_out(5415),
        VN2CN4_bit => VN_data_out(5416),
        VN2CN5_bit => VN_data_out(5417),
        VN2CN0_sign => VN_sign_out(5412),
        VN2CN1_sign => VN_sign_out(5413),
        VN2CN2_sign => VN_sign_out(5414),
        VN2CN3_sign => VN_sign_out(5415),
        VN2CN4_sign => VN_sign_out(5416),
        VN2CN5_sign => VN_sign_out(5417),
        codeword => codeword(902),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN903 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5423 downto 5418),
        Din0 => VN903_in0,
        Din1 => VN903_in1,
        Din2 => VN903_in2,
        Din3 => VN903_in3,
        Din4 => VN903_in4,
        Din5 => VN903_in5,
        VN2CN0_bit => VN_data_out(5418),
        VN2CN1_bit => VN_data_out(5419),
        VN2CN2_bit => VN_data_out(5420),
        VN2CN3_bit => VN_data_out(5421),
        VN2CN4_bit => VN_data_out(5422),
        VN2CN5_bit => VN_data_out(5423),
        VN2CN0_sign => VN_sign_out(5418),
        VN2CN1_sign => VN_sign_out(5419),
        VN2CN2_sign => VN_sign_out(5420),
        VN2CN3_sign => VN_sign_out(5421),
        VN2CN4_sign => VN_sign_out(5422),
        VN2CN5_sign => VN_sign_out(5423),
        codeword => codeword(903),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN904 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5429 downto 5424),
        Din0 => VN904_in0,
        Din1 => VN904_in1,
        Din2 => VN904_in2,
        Din3 => VN904_in3,
        Din4 => VN904_in4,
        Din5 => VN904_in5,
        VN2CN0_bit => VN_data_out(5424),
        VN2CN1_bit => VN_data_out(5425),
        VN2CN2_bit => VN_data_out(5426),
        VN2CN3_bit => VN_data_out(5427),
        VN2CN4_bit => VN_data_out(5428),
        VN2CN5_bit => VN_data_out(5429),
        VN2CN0_sign => VN_sign_out(5424),
        VN2CN1_sign => VN_sign_out(5425),
        VN2CN2_sign => VN_sign_out(5426),
        VN2CN3_sign => VN_sign_out(5427),
        VN2CN4_sign => VN_sign_out(5428),
        VN2CN5_sign => VN_sign_out(5429),
        codeword => codeword(904),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN905 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5435 downto 5430),
        Din0 => VN905_in0,
        Din1 => VN905_in1,
        Din2 => VN905_in2,
        Din3 => VN905_in3,
        Din4 => VN905_in4,
        Din5 => VN905_in5,
        VN2CN0_bit => VN_data_out(5430),
        VN2CN1_bit => VN_data_out(5431),
        VN2CN2_bit => VN_data_out(5432),
        VN2CN3_bit => VN_data_out(5433),
        VN2CN4_bit => VN_data_out(5434),
        VN2CN5_bit => VN_data_out(5435),
        VN2CN0_sign => VN_sign_out(5430),
        VN2CN1_sign => VN_sign_out(5431),
        VN2CN2_sign => VN_sign_out(5432),
        VN2CN3_sign => VN_sign_out(5433),
        VN2CN4_sign => VN_sign_out(5434),
        VN2CN5_sign => VN_sign_out(5435),
        codeword => codeword(905),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN906 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5441 downto 5436),
        Din0 => VN906_in0,
        Din1 => VN906_in1,
        Din2 => VN906_in2,
        Din3 => VN906_in3,
        Din4 => VN906_in4,
        Din5 => VN906_in5,
        VN2CN0_bit => VN_data_out(5436),
        VN2CN1_bit => VN_data_out(5437),
        VN2CN2_bit => VN_data_out(5438),
        VN2CN3_bit => VN_data_out(5439),
        VN2CN4_bit => VN_data_out(5440),
        VN2CN5_bit => VN_data_out(5441),
        VN2CN0_sign => VN_sign_out(5436),
        VN2CN1_sign => VN_sign_out(5437),
        VN2CN2_sign => VN_sign_out(5438),
        VN2CN3_sign => VN_sign_out(5439),
        VN2CN4_sign => VN_sign_out(5440),
        VN2CN5_sign => VN_sign_out(5441),
        codeword => codeword(906),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN907 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5447 downto 5442),
        Din0 => VN907_in0,
        Din1 => VN907_in1,
        Din2 => VN907_in2,
        Din3 => VN907_in3,
        Din4 => VN907_in4,
        Din5 => VN907_in5,
        VN2CN0_bit => VN_data_out(5442),
        VN2CN1_bit => VN_data_out(5443),
        VN2CN2_bit => VN_data_out(5444),
        VN2CN3_bit => VN_data_out(5445),
        VN2CN4_bit => VN_data_out(5446),
        VN2CN5_bit => VN_data_out(5447),
        VN2CN0_sign => VN_sign_out(5442),
        VN2CN1_sign => VN_sign_out(5443),
        VN2CN2_sign => VN_sign_out(5444),
        VN2CN3_sign => VN_sign_out(5445),
        VN2CN4_sign => VN_sign_out(5446),
        VN2CN5_sign => VN_sign_out(5447),
        codeword => codeword(907),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN908 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5453 downto 5448),
        Din0 => VN908_in0,
        Din1 => VN908_in1,
        Din2 => VN908_in2,
        Din3 => VN908_in3,
        Din4 => VN908_in4,
        Din5 => VN908_in5,
        VN2CN0_bit => VN_data_out(5448),
        VN2CN1_bit => VN_data_out(5449),
        VN2CN2_bit => VN_data_out(5450),
        VN2CN3_bit => VN_data_out(5451),
        VN2CN4_bit => VN_data_out(5452),
        VN2CN5_bit => VN_data_out(5453),
        VN2CN0_sign => VN_sign_out(5448),
        VN2CN1_sign => VN_sign_out(5449),
        VN2CN2_sign => VN_sign_out(5450),
        VN2CN3_sign => VN_sign_out(5451),
        VN2CN4_sign => VN_sign_out(5452),
        VN2CN5_sign => VN_sign_out(5453),
        codeword => codeword(908),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN909 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5459 downto 5454),
        Din0 => VN909_in0,
        Din1 => VN909_in1,
        Din2 => VN909_in2,
        Din3 => VN909_in3,
        Din4 => VN909_in4,
        Din5 => VN909_in5,
        VN2CN0_bit => VN_data_out(5454),
        VN2CN1_bit => VN_data_out(5455),
        VN2CN2_bit => VN_data_out(5456),
        VN2CN3_bit => VN_data_out(5457),
        VN2CN4_bit => VN_data_out(5458),
        VN2CN5_bit => VN_data_out(5459),
        VN2CN0_sign => VN_sign_out(5454),
        VN2CN1_sign => VN_sign_out(5455),
        VN2CN2_sign => VN_sign_out(5456),
        VN2CN3_sign => VN_sign_out(5457),
        VN2CN4_sign => VN_sign_out(5458),
        VN2CN5_sign => VN_sign_out(5459),
        codeword => codeword(909),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN910 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5465 downto 5460),
        Din0 => VN910_in0,
        Din1 => VN910_in1,
        Din2 => VN910_in2,
        Din3 => VN910_in3,
        Din4 => VN910_in4,
        Din5 => VN910_in5,
        VN2CN0_bit => VN_data_out(5460),
        VN2CN1_bit => VN_data_out(5461),
        VN2CN2_bit => VN_data_out(5462),
        VN2CN3_bit => VN_data_out(5463),
        VN2CN4_bit => VN_data_out(5464),
        VN2CN5_bit => VN_data_out(5465),
        VN2CN0_sign => VN_sign_out(5460),
        VN2CN1_sign => VN_sign_out(5461),
        VN2CN2_sign => VN_sign_out(5462),
        VN2CN3_sign => VN_sign_out(5463),
        VN2CN4_sign => VN_sign_out(5464),
        VN2CN5_sign => VN_sign_out(5465),
        codeword => codeword(910),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN911 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5471 downto 5466),
        Din0 => VN911_in0,
        Din1 => VN911_in1,
        Din2 => VN911_in2,
        Din3 => VN911_in3,
        Din4 => VN911_in4,
        Din5 => VN911_in5,
        VN2CN0_bit => VN_data_out(5466),
        VN2CN1_bit => VN_data_out(5467),
        VN2CN2_bit => VN_data_out(5468),
        VN2CN3_bit => VN_data_out(5469),
        VN2CN4_bit => VN_data_out(5470),
        VN2CN5_bit => VN_data_out(5471),
        VN2CN0_sign => VN_sign_out(5466),
        VN2CN1_sign => VN_sign_out(5467),
        VN2CN2_sign => VN_sign_out(5468),
        VN2CN3_sign => VN_sign_out(5469),
        VN2CN4_sign => VN_sign_out(5470),
        VN2CN5_sign => VN_sign_out(5471),
        codeword => codeword(911),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN912 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5477 downto 5472),
        Din0 => VN912_in0,
        Din1 => VN912_in1,
        Din2 => VN912_in2,
        Din3 => VN912_in3,
        Din4 => VN912_in4,
        Din5 => VN912_in5,
        VN2CN0_bit => VN_data_out(5472),
        VN2CN1_bit => VN_data_out(5473),
        VN2CN2_bit => VN_data_out(5474),
        VN2CN3_bit => VN_data_out(5475),
        VN2CN4_bit => VN_data_out(5476),
        VN2CN5_bit => VN_data_out(5477),
        VN2CN0_sign => VN_sign_out(5472),
        VN2CN1_sign => VN_sign_out(5473),
        VN2CN2_sign => VN_sign_out(5474),
        VN2CN3_sign => VN_sign_out(5475),
        VN2CN4_sign => VN_sign_out(5476),
        VN2CN5_sign => VN_sign_out(5477),
        codeword => codeword(912),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN913 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5483 downto 5478),
        Din0 => VN913_in0,
        Din1 => VN913_in1,
        Din2 => VN913_in2,
        Din3 => VN913_in3,
        Din4 => VN913_in4,
        Din5 => VN913_in5,
        VN2CN0_bit => VN_data_out(5478),
        VN2CN1_bit => VN_data_out(5479),
        VN2CN2_bit => VN_data_out(5480),
        VN2CN3_bit => VN_data_out(5481),
        VN2CN4_bit => VN_data_out(5482),
        VN2CN5_bit => VN_data_out(5483),
        VN2CN0_sign => VN_sign_out(5478),
        VN2CN1_sign => VN_sign_out(5479),
        VN2CN2_sign => VN_sign_out(5480),
        VN2CN3_sign => VN_sign_out(5481),
        VN2CN4_sign => VN_sign_out(5482),
        VN2CN5_sign => VN_sign_out(5483),
        codeword => codeword(913),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN914 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5489 downto 5484),
        Din0 => VN914_in0,
        Din1 => VN914_in1,
        Din2 => VN914_in2,
        Din3 => VN914_in3,
        Din4 => VN914_in4,
        Din5 => VN914_in5,
        VN2CN0_bit => VN_data_out(5484),
        VN2CN1_bit => VN_data_out(5485),
        VN2CN2_bit => VN_data_out(5486),
        VN2CN3_bit => VN_data_out(5487),
        VN2CN4_bit => VN_data_out(5488),
        VN2CN5_bit => VN_data_out(5489),
        VN2CN0_sign => VN_sign_out(5484),
        VN2CN1_sign => VN_sign_out(5485),
        VN2CN2_sign => VN_sign_out(5486),
        VN2CN3_sign => VN_sign_out(5487),
        VN2CN4_sign => VN_sign_out(5488),
        VN2CN5_sign => VN_sign_out(5489),
        codeword => codeword(914),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN915 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5495 downto 5490),
        Din0 => VN915_in0,
        Din1 => VN915_in1,
        Din2 => VN915_in2,
        Din3 => VN915_in3,
        Din4 => VN915_in4,
        Din5 => VN915_in5,
        VN2CN0_bit => VN_data_out(5490),
        VN2CN1_bit => VN_data_out(5491),
        VN2CN2_bit => VN_data_out(5492),
        VN2CN3_bit => VN_data_out(5493),
        VN2CN4_bit => VN_data_out(5494),
        VN2CN5_bit => VN_data_out(5495),
        VN2CN0_sign => VN_sign_out(5490),
        VN2CN1_sign => VN_sign_out(5491),
        VN2CN2_sign => VN_sign_out(5492),
        VN2CN3_sign => VN_sign_out(5493),
        VN2CN4_sign => VN_sign_out(5494),
        VN2CN5_sign => VN_sign_out(5495),
        codeword => codeword(915),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN916 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5501 downto 5496),
        Din0 => VN916_in0,
        Din1 => VN916_in1,
        Din2 => VN916_in2,
        Din3 => VN916_in3,
        Din4 => VN916_in4,
        Din5 => VN916_in5,
        VN2CN0_bit => VN_data_out(5496),
        VN2CN1_bit => VN_data_out(5497),
        VN2CN2_bit => VN_data_out(5498),
        VN2CN3_bit => VN_data_out(5499),
        VN2CN4_bit => VN_data_out(5500),
        VN2CN5_bit => VN_data_out(5501),
        VN2CN0_sign => VN_sign_out(5496),
        VN2CN1_sign => VN_sign_out(5497),
        VN2CN2_sign => VN_sign_out(5498),
        VN2CN3_sign => VN_sign_out(5499),
        VN2CN4_sign => VN_sign_out(5500),
        VN2CN5_sign => VN_sign_out(5501),
        codeword => codeword(916),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN917 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5507 downto 5502),
        Din0 => VN917_in0,
        Din1 => VN917_in1,
        Din2 => VN917_in2,
        Din3 => VN917_in3,
        Din4 => VN917_in4,
        Din5 => VN917_in5,
        VN2CN0_bit => VN_data_out(5502),
        VN2CN1_bit => VN_data_out(5503),
        VN2CN2_bit => VN_data_out(5504),
        VN2CN3_bit => VN_data_out(5505),
        VN2CN4_bit => VN_data_out(5506),
        VN2CN5_bit => VN_data_out(5507),
        VN2CN0_sign => VN_sign_out(5502),
        VN2CN1_sign => VN_sign_out(5503),
        VN2CN2_sign => VN_sign_out(5504),
        VN2CN3_sign => VN_sign_out(5505),
        VN2CN4_sign => VN_sign_out(5506),
        VN2CN5_sign => VN_sign_out(5507),
        codeword => codeword(917),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN918 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5513 downto 5508),
        Din0 => VN918_in0,
        Din1 => VN918_in1,
        Din2 => VN918_in2,
        Din3 => VN918_in3,
        Din4 => VN918_in4,
        Din5 => VN918_in5,
        VN2CN0_bit => VN_data_out(5508),
        VN2CN1_bit => VN_data_out(5509),
        VN2CN2_bit => VN_data_out(5510),
        VN2CN3_bit => VN_data_out(5511),
        VN2CN4_bit => VN_data_out(5512),
        VN2CN5_bit => VN_data_out(5513),
        VN2CN0_sign => VN_sign_out(5508),
        VN2CN1_sign => VN_sign_out(5509),
        VN2CN2_sign => VN_sign_out(5510),
        VN2CN3_sign => VN_sign_out(5511),
        VN2CN4_sign => VN_sign_out(5512),
        VN2CN5_sign => VN_sign_out(5513),
        codeword => codeword(918),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN919 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5519 downto 5514),
        Din0 => VN919_in0,
        Din1 => VN919_in1,
        Din2 => VN919_in2,
        Din3 => VN919_in3,
        Din4 => VN919_in4,
        Din5 => VN919_in5,
        VN2CN0_bit => VN_data_out(5514),
        VN2CN1_bit => VN_data_out(5515),
        VN2CN2_bit => VN_data_out(5516),
        VN2CN3_bit => VN_data_out(5517),
        VN2CN4_bit => VN_data_out(5518),
        VN2CN5_bit => VN_data_out(5519),
        VN2CN0_sign => VN_sign_out(5514),
        VN2CN1_sign => VN_sign_out(5515),
        VN2CN2_sign => VN_sign_out(5516),
        VN2CN3_sign => VN_sign_out(5517),
        VN2CN4_sign => VN_sign_out(5518),
        VN2CN5_sign => VN_sign_out(5519),
        codeword => codeword(919),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN920 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5525 downto 5520),
        Din0 => VN920_in0,
        Din1 => VN920_in1,
        Din2 => VN920_in2,
        Din3 => VN920_in3,
        Din4 => VN920_in4,
        Din5 => VN920_in5,
        VN2CN0_bit => VN_data_out(5520),
        VN2CN1_bit => VN_data_out(5521),
        VN2CN2_bit => VN_data_out(5522),
        VN2CN3_bit => VN_data_out(5523),
        VN2CN4_bit => VN_data_out(5524),
        VN2CN5_bit => VN_data_out(5525),
        VN2CN0_sign => VN_sign_out(5520),
        VN2CN1_sign => VN_sign_out(5521),
        VN2CN2_sign => VN_sign_out(5522),
        VN2CN3_sign => VN_sign_out(5523),
        VN2CN4_sign => VN_sign_out(5524),
        VN2CN5_sign => VN_sign_out(5525),
        codeword => codeword(920),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN921 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5531 downto 5526),
        Din0 => VN921_in0,
        Din1 => VN921_in1,
        Din2 => VN921_in2,
        Din3 => VN921_in3,
        Din4 => VN921_in4,
        Din5 => VN921_in5,
        VN2CN0_bit => VN_data_out(5526),
        VN2CN1_bit => VN_data_out(5527),
        VN2CN2_bit => VN_data_out(5528),
        VN2CN3_bit => VN_data_out(5529),
        VN2CN4_bit => VN_data_out(5530),
        VN2CN5_bit => VN_data_out(5531),
        VN2CN0_sign => VN_sign_out(5526),
        VN2CN1_sign => VN_sign_out(5527),
        VN2CN2_sign => VN_sign_out(5528),
        VN2CN3_sign => VN_sign_out(5529),
        VN2CN4_sign => VN_sign_out(5530),
        VN2CN5_sign => VN_sign_out(5531),
        codeword => codeword(921),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN922 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5537 downto 5532),
        Din0 => VN922_in0,
        Din1 => VN922_in1,
        Din2 => VN922_in2,
        Din3 => VN922_in3,
        Din4 => VN922_in4,
        Din5 => VN922_in5,
        VN2CN0_bit => VN_data_out(5532),
        VN2CN1_bit => VN_data_out(5533),
        VN2CN2_bit => VN_data_out(5534),
        VN2CN3_bit => VN_data_out(5535),
        VN2CN4_bit => VN_data_out(5536),
        VN2CN5_bit => VN_data_out(5537),
        VN2CN0_sign => VN_sign_out(5532),
        VN2CN1_sign => VN_sign_out(5533),
        VN2CN2_sign => VN_sign_out(5534),
        VN2CN3_sign => VN_sign_out(5535),
        VN2CN4_sign => VN_sign_out(5536),
        VN2CN5_sign => VN_sign_out(5537),
        codeword => codeword(922),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN923 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5543 downto 5538),
        Din0 => VN923_in0,
        Din1 => VN923_in1,
        Din2 => VN923_in2,
        Din3 => VN923_in3,
        Din4 => VN923_in4,
        Din5 => VN923_in5,
        VN2CN0_bit => VN_data_out(5538),
        VN2CN1_bit => VN_data_out(5539),
        VN2CN2_bit => VN_data_out(5540),
        VN2CN3_bit => VN_data_out(5541),
        VN2CN4_bit => VN_data_out(5542),
        VN2CN5_bit => VN_data_out(5543),
        VN2CN0_sign => VN_sign_out(5538),
        VN2CN1_sign => VN_sign_out(5539),
        VN2CN2_sign => VN_sign_out(5540),
        VN2CN3_sign => VN_sign_out(5541),
        VN2CN4_sign => VN_sign_out(5542),
        VN2CN5_sign => VN_sign_out(5543),
        codeword => codeword(923),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN924 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5549 downto 5544),
        Din0 => VN924_in0,
        Din1 => VN924_in1,
        Din2 => VN924_in2,
        Din3 => VN924_in3,
        Din4 => VN924_in4,
        Din5 => VN924_in5,
        VN2CN0_bit => VN_data_out(5544),
        VN2CN1_bit => VN_data_out(5545),
        VN2CN2_bit => VN_data_out(5546),
        VN2CN3_bit => VN_data_out(5547),
        VN2CN4_bit => VN_data_out(5548),
        VN2CN5_bit => VN_data_out(5549),
        VN2CN0_sign => VN_sign_out(5544),
        VN2CN1_sign => VN_sign_out(5545),
        VN2CN2_sign => VN_sign_out(5546),
        VN2CN3_sign => VN_sign_out(5547),
        VN2CN4_sign => VN_sign_out(5548),
        VN2CN5_sign => VN_sign_out(5549),
        codeword => codeword(924),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN925 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5555 downto 5550),
        Din0 => VN925_in0,
        Din1 => VN925_in1,
        Din2 => VN925_in2,
        Din3 => VN925_in3,
        Din4 => VN925_in4,
        Din5 => VN925_in5,
        VN2CN0_bit => VN_data_out(5550),
        VN2CN1_bit => VN_data_out(5551),
        VN2CN2_bit => VN_data_out(5552),
        VN2CN3_bit => VN_data_out(5553),
        VN2CN4_bit => VN_data_out(5554),
        VN2CN5_bit => VN_data_out(5555),
        VN2CN0_sign => VN_sign_out(5550),
        VN2CN1_sign => VN_sign_out(5551),
        VN2CN2_sign => VN_sign_out(5552),
        VN2CN3_sign => VN_sign_out(5553),
        VN2CN4_sign => VN_sign_out(5554),
        VN2CN5_sign => VN_sign_out(5555),
        codeword => codeword(925),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN926 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5561 downto 5556),
        Din0 => VN926_in0,
        Din1 => VN926_in1,
        Din2 => VN926_in2,
        Din3 => VN926_in3,
        Din4 => VN926_in4,
        Din5 => VN926_in5,
        VN2CN0_bit => VN_data_out(5556),
        VN2CN1_bit => VN_data_out(5557),
        VN2CN2_bit => VN_data_out(5558),
        VN2CN3_bit => VN_data_out(5559),
        VN2CN4_bit => VN_data_out(5560),
        VN2CN5_bit => VN_data_out(5561),
        VN2CN0_sign => VN_sign_out(5556),
        VN2CN1_sign => VN_sign_out(5557),
        VN2CN2_sign => VN_sign_out(5558),
        VN2CN3_sign => VN_sign_out(5559),
        VN2CN4_sign => VN_sign_out(5560),
        VN2CN5_sign => VN_sign_out(5561),
        codeword => codeword(926),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN927 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5567 downto 5562),
        Din0 => VN927_in0,
        Din1 => VN927_in1,
        Din2 => VN927_in2,
        Din3 => VN927_in3,
        Din4 => VN927_in4,
        Din5 => VN927_in5,
        VN2CN0_bit => VN_data_out(5562),
        VN2CN1_bit => VN_data_out(5563),
        VN2CN2_bit => VN_data_out(5564),
        VN2CN3_bit => VN_data_out(5565),
        VN2CN4_bit => VN_data_out(5566),
        VN2CN5_bit => VN_data_out(5567),
        VN2CN0_sign => VN_sign_out(5562),
        VN2CN1_sign => VN_sign_out(5563),
        VN2CN2_sign => VN_sign_out(5564),
        VN2CN3_sign => VN_sign_out(5565),
        VN2CN4_sign => VN_sign_out(5566),
        VN2CN5_sign => VN_sign_out(5567),
        codeword => codeword(927),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN928 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5573 downto 5568),
        Din0 => VN928_in0,
        Din1 => VN928_in1,
        Din2 => VN928_in2,
        Din3 => VN928_in3,
        Din4 => VN928_in4,
        Din5 => VN928_in5,
        VN2CN0_bit => VN_data_out(5568),
        VN2CN1_bit => VN_data_out(5569),
        VN2CN2_bit => VN_data_out(5570),
        VN2CN3_bit => VN_data_out(5571),
        VN2CN4_bit => VN_data_out(5572),
        VN2CN5_bit => VN_data_out(5573),
        VN2CN0_sign => VN_sign_out(5568),
        VN2CN1_sign => VN_sign_out(5569),
        VN2CN2_sign => VN_sign_out(5570),
        VN2CN3_sign => VN_sign_out(5571),
        VN2CN4_sign => VN_sign_out(5572),
        VN2CN5_sign => VN_sign_out(5573),
        codeword => codeword(928),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN929 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5579 downto 5574),
        Din0 => VN929_in0,
        Din1 => VN929_in1,
        Din2 => VN929_in2,
        Din3 => VN929_in3,
        Din4 => VN929_in4,
        Din5 => VN929_in5,
        VN2CN0_bit => VN_data_out(5574),
        VN2CN1_bit => VN_data_out(5575),
        VN2CN2_bit => VN_data_out(5576),
        VN2CN3_bit => VN_data_out(5577),
        VN2CN4_bit => VN_data_out(5578),
        VN2CN5_bit => VN_data_out(5579),
        VN2CN0_sign => VN_sign_out(5574),
        VN2CN1_sign => VN_sign_out(5575),
        VN2CN2_sign => VN_sign_out(5576),
        VN2CN3_sign => VN_sign_out(5577),
        VN2CN4_sign => VN_sign_out(5578),
        VN2CN5_sign => VN_sign_out(5579),
        codeword => codeword(929),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN930 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5585 downto 5580),
        Din0 => VN930_in0,
        Din1 => VN930_in1,
        Din2 => VN930_in2,
        Din3 => VN930_in3,
        Din4 => VN930_in4,
        Din5 => VN930_in5,
        VN2CN0_bit => VN_data_out(5580),
        VN2CN1_bit => VN_data_out(5581),
        VN2CN2_bit => VN_data_out(5582),
        VN2CN3_bit => VN_data_out(5583),
        VN2CN4_bit => VN_data_out(5584),
        VN2CN5_bit => VN_data_out(5585),
        VN2CN0_sign => VN_sign_out(5580),
        VN2CN1_sign => VN_sign_out(5581),
        VN2CN2_sign => VN_sign_out(5582),
        VN2CN3_sign => VN_sign_out(5583),
        VN2CN4_sign => VN_sign_out(5584),
        VN2CN5_sign => VN_sign_out(5585),
        codeword => codeword(930),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN931 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5591 downto 5586),
        Din0 => VN931_in0,
        Din1 => VN931_in1,
        Din2 => VN931_in2,
        Din3 => VN931_in3,
        Din4 => VN931_in4,
        Din5 => VN931_in5,
        VN2CN0_bit => VN_data_out(5586),
        VN2CN1_bit => VN_data_out(5587),
        VN2CN2_bit => VN_data_out(5588),
        VN2CN3_bit => VN_data_out(5589),
        VN2CN4_bit => VN_data_out(5590),
        VN2CN5_bit => VN_data_out(5591),
        VN2CN0_sign => VN_sign_out(5586),
        VN2CN1_sign => VN_sign_out(5587),
        VN2CN2_sign => VN_sign_out(5588),
        VN2CN3_sign => VN_sign_out(5589),
        VN2CN4_sign => VN_sign_out(5590),
        VN2CN5_sign => VN_sign_out(5591),
        codeword => codeword(931),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN932 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5597 downto 5592),
        Din0 => VN932_in0,
        Din1 => VN932_in1,
        Din2 => VN932_in2,
        Din3 => VN932_in3,
        Din4 => VN932_in4,
        Din5 => VN932_in5,
        VN2CN0_bit => VN_data_out(5592),
        VN2CN1_bit => VN_data_out(5593),
        VN2CN2_bit => VN_data_out(5594),
        VN2CN3_bit => VN_data_out(5595),
        VN2CN4_bit => VN_data_out(5596),
        VN2CN5_bit => VN_data_out(5597),
        VN2CN0_sign => VN_sign_out(5592),
        VN2CN1_sign => VN_sign_out(5593),
        VN2CN2_sign => VN_sign_out(5594),
        VN2CN3_sign => VN_sign_out(5595),
        VN2CN4_sign => VN_sign_out(5596),
        VN2CN5_sign => VN_sign_out(5597),
        codeword => codeword(932),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN933 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5603 downto 5598),
        Din0 => VN933_in0,
        Din1 => VN933_in1,
        Din2 => VN933_in2,
        Din3 => VN933_in3,
        Din4 => VN933_in4,
        Din5 => VN933_in5,
        VN2CN0_bit => VN_data_out(5598),
        VN2CN1_bit => VN_data_out(5599),
        VN2CN2_bit => VN_data_out(5600),
        VN2CN3_bit => VN_data_out(5601),
        VN2CN4_bit => VN_data_out(5602),
        VN2CN5_bit => VN_data_out(5603),
        VN2CN0_sign => VN_sign_out(5598),
        VN2CN1_sign => VN_sign_out(5599),
        VN2CN2_sign => VN_sign_out(5600),
        VN2CN3_sign => VN_sign_out(5601),
        VN2CN4_sign => VN_sign_out(5602),
        VN2CN5_sign => VN_sign_out(5603),
        codeword => codeword(933),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN934 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5609 downto 5604),
        Din0 => VN934_in0,
        Din1 => VN934_in1,
        Din2 => VN934_in2,
        Din3 => VN934_in3,
        Din4 => VN934_in4,
        Din5 => VN934_in5,
        VN2CN0_bit => VN_data_out(5604),
        VN2CN1_bit => VN_data_out(5605),
        VN2CN2_bit => VN_data_out(5606),
        VN2CN3_bit => VN_data_out(5607),
        VN2CN4_bit => VN_data_out(5608),
        VN2CN5_bit => VN_data_out(5609),
        VN2CN0_sign => VN_sign_out(5604),
        VN2CN1_sign => VN_sign_out(5605),
        VN2CN2_sign => VN_sign_out(5606),
        VN2CN3_sign => VN_sign_out(5607),
        VN2CN4_sign => VN_sign_out(5608),
        VN2CN5_sign => VN_sign_out(5609),
        codeword => codeword(934),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN935 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5615 downto 5610),
        Din0 => VN935_in0,
        Din1 => VN935_in1,
        Din2 => VN935_in2,
        Din3 => VN935_in3,
        Din4 => VN935_in4,
        Din5 => VN935_in5,
        VN2CN0_bit => VN_data_out(5610),
        VN2CN1_bit => VN_data_out(5611),
        VN2CN2_bit => VN_data_out(5612),
        VN2CN3_bit => VN_data_out(5613),
        VN2CN4_bit => VN_data_out(5614),
        VN2CN5_bit => VN_data_out(5615),
        VN2CN0_sign => VN_sign_out(5610),
        VN2CN1_sign => VN_sign_out(5611),
        VN2CN2_sign => VN_sign_out(5612),
        VN2CN3_sign => VN_sign_out(5613),
        VN2CN4_sign => VN_sign_out(5614),
        VN2CN5_sign => VN_sign_out(5615),
        codeword => codeword(935),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN936 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5621 downto 5616),
        Din0 => VN936_in0,
        Din1 => VN936_in1,
        Din2 => VN936_in2,
        Din3 => VN936_in3,
        Din4 => VN936_in4,
        Din5 => VN936_in5,
        VN2CN0_bit => VN_data_out(5616),
        VN2CN1_bit => VN_data_out(5617),
        VN2CN2_bit => VN_data_out(5618),
        VN2CN3_bit => VN_data_out(5619),
        VN2CN4_bit => VN_data_out(5620),
        VN2CN5_bit => VN_data_out(5621),
        VN2CN0_sign => VN_sign_out(5616),
        VN2CN1_sign => VN_sign_out(5617),
        VN2CN2_sign => VN_sign_out(5618),
        VN2CN3_sign => VN_sign_out(5619),
        VN2CN4_sign => VN_sign_out(5620),
        VN2CN5_sign => VN_sign_out(5621),
        codeword => codeword(936),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN937 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5627 downto 5622),
        Din0 => VN937_in0,
        Din1 => VN937_in1,
        Din2 => VN937_in2,
        Din3 => VN937_in3,
        Din4 => VN937_in4,
        Din5 => VN937_in5,
        VN2CN0_bit => VN_data_out(5622),
        VN2CN1_bit => VN_data_out(5623),
        VN2CN2_bit => VN_data_out(5624),
        VN2CN3_bit => VN_data_out(5625),
        VN2CN4_bit => VN_data_out(5626),
        VN2CN5_bit => VN_data_out(5627),
        VN2CN0_sign => VN_sign_out(5622),
        VN2CN1_sign => VN_sign_out(5623),
        VN2CN2_sign => VN_sign_out(5624),
        VN2CN3_sign => VN_sign_out(5625),
        VN2CN4_sign => VN_sign_out(5626),
        VN2CN5_sign => VN_sign_out(5627),
        codeword => codeword(937),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN938 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5633 downto 5628),
        Din0 => VN938_in0,
        Din1 => VN938_in1,
        Din2 => VN938_in2,
        Din3 => VN938_in3,
        Din4 => VN938_in4,
        Din5 => VN938_in5,
        VN2CN0_bit => VN_data_out(5628),
        VN2CN1_bit => VN_data_out(5629),
        VN2CN2_bit => VN_data_out(5630),
        VN2CN3_bit => VN_data_out(5631),
        VN2CN4_bit => VN_data_out(5632),
        VN2CN5_bit => VN_data_out(5633),
        VN2CN0_sign => VN_sign_out(5628),
        VN2CN1_sign => VN_sign_out(5629),
        VN2CN2_sign => VN_sign_out(5630),
        VN2CN3_sign => VN_sign_out(5631),
        VN2CN4_sign => VN_sign_out(5632),
        VN2CN5_sign => VN_sign_out(5633),
        codeword => codeword(938),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN939 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5639 downto 5634),
        Din0 => VN939_in0,
        Din1 => VN939_in1,
        Din2 => VN939_in2,
        Din3 => VN939_in3,
        Din4 => VN939_in4,
        Din5 => VN939_in5,
        VN2CN0_bit => VN_data_out(5634),
        VN2CN1_bit => VN_data_out(5635),
        VN2CN2_bit => VN_data_out(5636),
        VN2CN3_bit => VN_data_out(5637),
        VN2CN4_bit => VN_data_out(5638),
        VN2CN5_bit => VN_data_out(5639),
        VN2CN0_sign => VN_sign_out(5634),
        VN2CN1_sign => VN_sign_out(5635),
        VN2CN2_sign => VN_sign_out(5636),
        VN2CN3_sign => VN_sign_out(5637),
        VN2CN4_sign => VN_sign_out(5638),
        VN2CN5_sign => VN_sign_out(5639),
        codeword => codeword(939),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN940 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5645 downto 5640),
        Din0 => VN940_in0,
        Din1 => VN940_in1,
        Din2 => VN940_in2,
        Din3 => VN940_in3,
        Din4 => VN940_in4,
        Din5 => VN940_in5,
        VN2CN0_bit => VN_data_out(5640),
        VN2CN1_bit => VN_data_out(5641),
        VN2CN2_bit => VN_data_out(5642),
        VN2CN3_bit => VN_data_out(5643),
        VN2CN4_bit => VN_data_out(5644),
        VN2CN5_bit => VN_data_out(5645),
        VN2CN0_sign => VN_sign_out(5640),
        VN2CN1_sign => VN_sign_out(5641),
        VN2CN2_sign => VN_sign_out(5642),
        VN2CN3_sign => VN_sign_out(5643),
        VN2CN4_sign => VN_sign_out(5644),
        VN2CN5_sign => VN_sign_out(5645),
        codeword => codeword(940),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN941 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5651 downto 5646),
        Din0 => VN941_in0,
        Din1 => VN941_in1,
        Din2 => VN941_in2,
        Din3 => VN941_in3,
        Din4 => VN941_in4,
        Din5 => VN941_in5,
        VN2CN0_bit => VN_data_out(5646),
        VN2CN1_bit => VN_data_out(5647),
        VN2CN2_bit => VN_data_out(5648),
        VN2CN3_bit => VN_data_out(5649),
        VN2CN4_bit => VN_data_out(5650),
        VN2CN5_bit => VN_data_out(5651),
        VN2CN0_sign => VN_sign_out(5646),
        VN2CN1_sign => VN_sign_out(5647),
        VN2CN2_sign => VN_sign_out(5648),
        VN2CN3_sign => VN_sign_out(5649),
        VN2CN4_sign => VN_sign_out(5650),
        VN2CN5_sign => VN_sign_out(5651),
        codeword => codeword(941),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN942 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5657 downto 5652),
        Din0 => VN942_in0,
        Din1 => VN942_in1,
        Din2 => VN942_in2,
        Din3 => VN942_in3,
        Din4 => VN942_in4,
        Din5 => VN942_in5,
        VN2CN0_bit => VN_data_out(5652),
        VN2CN1_bit => VN_data_out(5653),
        VN2CN2_bit => VN_data_out(5654),
        VN2CN3_bit => VN_data_out(5655),
        VN2CN4_bit => VN_data_out(5656),
        VN2CN5_bit => VN_data_out(5657),
        VN2CN0_sign => VN_sign_out(5652),
        VN2CN1_sign => VN_sign_out(5653),
        VN2CN2_sign => VN_sign_out(5654),
        VN2CN3_sign => VN_sign_out(5655),
        VN2CN4_sign => VN_sign_out(5656),
        VN2CN5_sign => VN_sign_out(5657),
        codeword => codeword(942),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN943 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5663 downto 5658),
        Din0 => VN943_in0,
        Din1 => VN943_in1,
        Din2 => VN943_in2,
        Din3 => VN943_in3,
        Din4 => VN943_in4,
        Din5 => VN943_in5,
        VN2CN0_bit => VN_data_out(5658),
        VN2CN1_bit => VN_data_out(5659),
        VN2CN2_bit => VN_data_out(5660),
        VN2CN3_bit => VN_data_out(5661),
        VN2CN4_bit => VN_data_out(5662),
        VN2CN5_bit => VN_data_out(5663),
        VN2CN0_sign => VN_sign_out(5658),
        VN2CN1_sign => VN_sign_out(5659),
        VN2CN2_sign => VN_sign_out(5660),
        VN2CN3_sign => VN_sign_out(5661),
        VN2CN4_sign => VN_sign_out(5662),
        VN2CN5_sign => VN_sign_out(5663),
        codeword => codeword(943),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN944 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5669 downto 5664),
        Din0 => VN944_in0,
        Din1 => VN944_in1,
        Din2 => VN944_in2,
        Din3 => VN944_in3,
        Din4 => VN944_in4,
        Din5 => VN944_in5,
        VN2CN0_bit => VN_data_out(5664),
        VN2CN1_bit => VN_data_out(5665),
        VN2CN2_bit => VN_data_out(5666),
        VN2CN3_bit => VN_data_out(5667),
        VN2CN4_bit => VN_data_out(5668),
        VN2CN5_bit => VN_data_out(5669),
        VN2CN0_sign => VN_sign_out(5664),
        VN2CN1_sign => VN_sign_out(5665),
        VN2CN2_sign => VN_sign_out(5666),
        VN2CN3_sign => VN_sign_out(5667),
        VN2CN4_sign => VN_sign_out(5668),
        VN2CN5_sign => VN_sign_out(5669),
        codeword => codeword(944),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN945 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5675 downto 5670),
        Din0 => VN945_in0,
        Din1 => VN945_in1,
        Din2 => VN945_in2,
        Din3 => VN945_in3,
        Din4 => VN945_in4,
        Din5 => VN945_in5,
        VN2CN0_bit => VN_data_out(5670),
        VN2CN1_bit => VN_data_out(5671),
        VN2CN2_bit => VN_data_out(5672),
        VN2CN3_bit => VN_data_out(5673),
        VN2CN4_bit => VN_data_out(5674),
        VN2CN5_bit => VN_data_out(5675),
        VN2CN0_sign => VN_sign_out(5670),
        VN2CN1_sign => VN_sign_out(5671),
        VN2CN2_sign => VN_sign_out(5672),
        VN2CN3_sign => VN_sign_out(5673),
        VN2CN4_sign => VN_sign_out(5674),
        VN2CN5_sign => VN_sign_out(5675),
        codeword => codeword(945),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN946 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5681 downto 5676),
        Din0 => VN946_in0,
        Din1 => VN946_in1,
        Din2 => VN946_in2,
        Din3 => VN946_in3,
        Din4 => VN946_in4,
        Din5 => VN946_in5,
        VN2CN0_bit => VN_data_out(5676),
        VN2CN1_bit => VN_data_out(5677),
        VN2CN2_bit => VN_data_out(5678),
        VN2CN3_bit => VN_data_out(5679),
        VN2CN4_bit => VN_data_out(5680),
        VN2CN5_bit => VN_data_out(5681),
        VN2CN0_sign => VN_sign_out(5676),
        VN2CN1_sign => VN_sign_out(5677),
        VN2CN2_sign => VN_sign_out(5678),
        VN2CN3_sign => VN_sign_out(5679),
        VN2CN4_sign => VN_sign_out(5680),
        VN2CN5_sign => VN_sign_out(5681),
        codeword => codeword(946),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN947 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5687 downto 5682),
        Din0 => VN947_in0,
        Din1 => VN947_in1,
        Din2 => VN947_in2,
        Din3 => VN947_in3,
        Din4 => VN947_in4,
        Din5 => VN947_in5,
        VN2CN0_bit => VN_data_out(5682),
        VN2CN1_bit => VN_data_out(5683),
        VN2CN2_bit => VN_data_out(5684),
        VN2CN3_bit => VN_data_out(5685),
        VN2CN4_bit => VN_data_out(5686),
        VN2CN5_bit => VN_data_out(5687),
        VN2CN0_sign => VN_sign_out(5682),
        VN2CN1_sign => VN_sign_out(5683),
        VN2CN2_sign => VN_sign_out(5684),
        VN2CN3_sign => VN_sign_out(5685),
        VN2CN4_sign => VN_sign_out(5686),
        VN2CN5_sign => VN_sign_out(5687),
        codeword => codeword(947),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN948 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5693 downto 5688),
        Din0 => VN948_in0,
        Din1 => VN948_in1,
        Din2 => VN948_in2,
        Din3 => VN948_in3,
        Din4 => VN948_in4,
        Din5 => VN948_in5,
        VN2CN0_bit => VN_data_out(5688),
        VN2CN1_bit => VN_data_out(5689),
        VN2CN2_bit => VN_data_out(5690),
        VN2CN3_bit => VN_data_out(5691),
        VN2CN4_bit => VN_data_out(5692),
        VN2CN5_bit => VN_data_out(5693),
        VN2CN0_sign => VN_sign_out(5688),
        VN2CN1_sign => VN_sign_out(5689),
        VN2CN2_sign => VN_sign_out(5690),
        VN2CN3_sign => VN_sign_out(5691),
        VN2CN4_sign => VN_sign_out(5692),
        VN2CN5_sign => VN_sign_out(5693),
        codeword => codeword(948),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN949 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5699 downto 5694),
        Din0 => VN949_in0,
        Din1 => VN949_in1,
        Din2 => VN949_in2,
        Din3 => VN949_in3,
        Din4 => VN949_in4,
        Din5 => VN949_in5,
        VN2CN0_bit => VN_data_out(5694),
        VN2CN1_bit => VN_data_out(5695),
        VN2CN2_bit => VN_data_out(5696),
        VN2CN3_bit => VN_data_out(5697),
        VN2CN4_bit => VN_data_out(5698),
        VN2CN5_bit => VN_data_out(5699),
        VN2CN0_sign => VN_sign_out(5694),
        VN2CN1_sign => VN_sign_out(5695),
        VN2CN2_sign => VN_sign_out(5696),
        VN2CN3_sign => VN_sign_out(5697),
        VN2CN4_sign => VN_sign_out(5698),
        VN2CN5_sign => VN_sign_out(5699),
        codeword => codeword(949),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN950 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5705 downto 5700),
        Din0 => VN950_in0,
        Din1 => VN950_in1,
        Din2 => VN950_in2,
        Din3 => VN950_in3,
        Din4 => VN950_in4,
        Din5 => VN950_in5,
        VN2CN0_bit => VN_data_out(5700),
        VN2CN1_bit => VN_data_out(5701),
        VN2CN2_bit => VN_data_out(5702),
        VN2CN3_bit => VN_data_out(5703),
        VN2CN4_bit => VN_data_out(5704),
        VN2CN5_bit => VN_data_out(5705),
        VN2CN0_sign => VN_sign_out(5700),
        VN2CN1_sign => VN_sign_out(5701),
        VN2CN2_sign => VN_sign_out(5702),
        VN2CN3_sign => VN_sign_out(5703),
        VN2CN4_sign => VN_sign_out(5704),
        VN2CN5_sign => VN_sign_out(5705),
        codeword => codeword(950),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN951 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5711 downto 5706),
        Din0 => VN951_in0,
        Din1 => VN951_in1,
        Din2 => VN951_in2,
        Din3 => VN951_in3,
        Din4 => VN951_in4,
        Din5 => VN951_in5,
        VN2CN0_bit => VN_data_out(5706),
        VN2CN1_bit => VN_data_out(5707),
        VN2CN2_bit => VN_data_out(5708),
        VN2CN3_bit => VN_data_out(5709),
        VN2CN4_bit => VN_data_out(5710),
        VN2CN5_bit => VN_data_out(5711),
        VN2CN0_sign => VN_sign_out(5706),
        VN2CN1_sign => VN_sign_out(5707),
        VN2CN2_sign => VN_sign_out(5708),
        VN2CN3_sign => VN_sign_out(5709),
        VN2CN4_sign => VN_sign_out(5710),
        VN2CN5_sign => VN_sign_out(5711),
        codeword => codeword(951),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN952 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5717 downto 5712),
        Din0 => VN952_in0,
        Din1 => VN952_in1,
        Din2 => VN952_in2,
        Din3 => VN952_in3,
        Din4 => VN952_in4,
        Din5 => VN952_in5,
        VN2CN0_bit => VN_data_out(5712),
        VN2CN1_bit => VN_data_out(5713),
        VN2CN2_bit => VN_data_out(5714),
        VN2CN3_bit => VN_data_out(5715),
        VN2CN4_bit => VN_data_out(5716),
        VN2CN5_bit => VN_data_out(5717),
        VN2CN0_sign => VN_sign_out(5712),
        VN2CN1_sign => VN_sign_out(5713),
        VN2CN2_sign => VN_sign_out(5714),
        VN2CN3_sign => VN_sign_out(5715),
        VN2CN4_sign => VN_sign_out(5716),
        VN2CN5_sign => VN_sign_out(5717),
        codeword => codeword(952),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN953 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5723 downto 5718),
        Din0 => VN953_in0,
        Din1 => VN953_in1,
        Din2 => VN953_in2,
        Din3 => VN953_in3,
        Din4 => VN953_in4,
        Din5 => VN953_in5,
        VN2CN0_bit => VN_data_out(5718),
        VN2CN1_bit => VN_data_out(5719),
        VN2CN2_bit => VN_data_out(5720),
        VN2CN3_bit => VN_data_out(5721),
        VN2CN4_bit => VN_data_out(5722),
        VN2CN5_bit => VN_data_out(5723),
        VN2CN0_sign => VN_sign_out(5718),
        VN2CN1_sign => VN_sign_out(5719),
        VN2CN2_sign => VN_sign_out(5720),
        VN2CN3_sign => VN_sign_out(5721),
        VN2CN4_sign => VN_sign_out(5722),
        VN2CN5_sign => VN_sign_out(5723),
        codeword => codeword(953),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN954 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5729 downto 5724),
        Din0 => VN954_in0,
        Din1 => VN954_in1,
        Din2 => VN954_in2,
        Din3 => VN954_in3,
        Din4 => VN954_in4,
        Din5 => VN954_in5,
        VN2CN0_bit => VN_data_out(5724),
        VN2CN1_bit => VN_data_out(5725),
        VN2CN2_bit => VN_data_out(5726),
        VN2CN3_bit => VN_data_out(5727),
        VN2CN4_bit => VN_data_out(5728),
        VN2CN5_bit => VN_data_out(5729),
        VN2CN0_sign => VN_sign_out(5724),
        VN2CN1_sign => VN_sign_out(5725),
        VN2CN2_sign => VN_sign_out(5726),
        VN2CN3_sign => VN_sign_out(5727),
        VN2CN4_sign => VN_sign_out(5728),
        VN2CN5_sign => VN_sign_out(5729),
        codeword => codeword(954),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN955 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5735 downto 5730),
        Din0 => VN955_in0,
        Din1 => VN955_in1,
        Din2 => VN955_in2,
        Din3 => VN955_in3,
        Din4 => VN955_in4,
        Din5 => VN955_in5,
        VN2CN0_bit => VN_data_out(5730),
        VN2CN1_bit => VN_data_out(5731),
        VN2CN2_bit => VN_data_out(5732),
        VN2CN3_bit => VN_data_out(5733),
        VN2CN4_bit => VN_data_out(5734),
        VN2CN5_bit => VN_data_out(5735),
        VN2CN0_sign => VN_sign_out(5730),
        VN2CN1_sign => VN_sign_out(5731),
        VN2CN2_sign => VN_sign_out(5732),
        VN2CN3_sign => VN_sign_out(5733),
        VN2CN4_sign => VN_sign_out(5734),
        VN2CN5_sign => VN_sign_out(5735),
        codeword => codeword(955),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN956 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5741 downto 5736),
        Din0 => VN956_in0,
        Din1 => VN956_in1,
        Din2 => VN956_in2,
        Din3 => VN956_in3,
        Din4 => VN956_in4,
        Din5 => VN956_in5,
        VN2CN0_bit => VN_data_out(5736),
        VN2CN1_bit => VN_data_out(5737),
        VN2CN2_bit => VN_data_out(5738),
        VN2CN3_bit => VN_data_out(5739),
        VN2CN4_bit => VN_data_out(5740),
        VN2CN5_bit => VN_data_out(5741),
        VN2CN0_sign => VN_sign_out(5736),
        VN2CN1_sign => VN_sign_out(5737),
        VN2CN2_sign => VN_sign_out(5738),
        VN2CN3_sign => VN_sign_out(5739),
        VN2CN4_sign => VN_sign_out(5740),
        VN2CN5_sign => VN_sign_out(5741),
        codeword => codeword(956),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN957 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5747 downto 5742),
        Din0 => VN957_in0,
        Din1 => VN957_in1,
        Din2 => VN957_in2,
        Din3 => VN957_in3,
        Din4 => VN957_in4,
        Din5 => VN957_in5,
        VN2CN0_bit => VN_data_out(5742),
        VN2CN1_bit => VN_data_out(5743),
        VN2CN2_bit => VN_data_out(5744),
        VN2CN3_bit => VN_data_out(5745),
        VN2CN4_bit => VN_data_out(5746),
        VN2CN5_bit => VN_data_out(5747),
        VN2CN0_sign => VN_sign_out(5742),
        VN2CN1_sign => VN_sign_out(5743),
        VN2CN2_sign => VN_sign_out(5744),
        VN2CN3_sign => VN_sign_out(5745),
        VN2CN4_sign => VN_sign_out(5746),
        VN2CN5_sign => VN_sign_out(5747),
        codeword => codeword(957),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN958 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5753 downto 5748),
        Din0 => VN958_in0,
        Din1 => VN958_in1,
        Din2 => VN958_in2,
        Din3 => VN958_in3,
        Din4 => VN958_in4,
        Din5 => VN958_in5,
        VN2CN0_bit => VN_data_out(5748),
        VN2CN1_bit => VN_data_out(5749),
        VN2CN2_bit => VN_data_out(5750),
        VN2CN3_bit => VN_data_out(5751),
        VN2CN4_bit => VN_data_out(5752),
        VN2CN5_bit => VN_data_out(5753),
        VN2CN0_sign => VN_sign_out(5748),
        VN2CN1_sign => VN_sign_out(5749),
        VN2CN2_sign => VN_sign_out(5750),
        VN2CN3_sign => VN_sign_out(5751),
        VN2CN4_sign => VN_sign_out(5752),
        VN2CN5_sign => VN_sign_out(5753),
        codeword => codeword(958),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN959 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5759 downto 5754),
        Din0 => VN959_in0,
        Din1 => VN959_in1,
        Din2 => VN959_in2,
        Din3 => VN959_in3,
        Din4 => VN959_in4,
        Din5 => VN959_in5,
        VN2CN0_bit => VN_data_out(5754),
        VN2CN1_bit => VN_data_out(5755),
        VN2CN2_bit => VN_data_out(5756),
        VN2CN3_bit => VN_data_out(5757),
        VN2CN4_bit => VN_data_out(5758),
        VN2CN5_bit => VN_data_out(5759),
        VN2CN0_sign => VN_sign_out(5754),
        VN2CN1_sign => VN_sign_out(5755),
        VN2CN2_sign => VN_sign_out(5756),
        VN2CN3_sign => VN_sign_out(5757),
        VN2CN4_sign => VN_sign_out(5758),
        VN2CN5_sign => VN_sign_out(5759),
        codeword => codeword(959),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN960 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5765 downto 5760),
        Din0 => VN960_in0,
        Din1 => VN960_in1,
        Din2 => VN960_in2,
        Din3 => VN960_in3,
        Din4 => VN960_in4,
        Din5 => VN960_in5,
        VN2CN0_bit => VN_data_out(5760),
        VN2CN1_bit => VN_data_out(5761),
        VN2CN2_bit => VN_data_out(5762),
        VN2CN3_bit => VN_data_out(5763),
        VN2CN4_bit => VN_data_out(5764),
        VN2CN5_bit => VN_data_out(5765),
        VN2CN0_sign => VN_sign_out(5760),
        VN2CN1_sign => VN_sign_out(5761),
        VN2CN2_sign => VN_sign_out(5762),
        VN2CN3_sign => VN_sign_out(5763),
        VN2CN4_sign => VN_sign_out(5764),
        VN2CN5_sign => VN_sign_out(5765),
        codeword => codeword(960),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN961 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5771 downto 5766),
        Din0 => VN961_in0,
        Din1 => VN961_in1,
        Din2 => VN961_in2,
        Din3 => VN961_in3,
        Din4 => VN961_in4,
        Din5 => VN961_in5,
        VN2CN0_bit => VN_data_out(5766),
        VN2CN1_bit => VN_data_out(5767),
        VN2CN2_bit => VN_data_out(5768),
        VN2CN3_bit => VN_data_out(5769),
        VN2CN4_bit => VN_data_out(5770),
        VN2CN5_bit => VN_data_out(5771),
        VN2CN0_sign => VN_sign_out(5766),
        VN2CN1_sign => VN_sign_out(5767),
        VN2CN2_sign => VN_sign_out(5768),
        VN2CN3_sign => VN_sign_out(5769),
        VN2CN4_sign => VN_sign_out(5770),
        VN2CN5_sign => VN_sign_out(5771),
        codeword => codeword(961),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN962 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5777 downto 5772),
        Din0 => VN962_in0,
        Din1 => VN962_in1,
        Din2 => VN962_in2,
        Din3 => VN962_in3,
        Din4 => VN962_in4,
        Din5 => VN962_in5,
        VN2CN0_bit => VN_data_out(5772),
        VN2CN1_bit => VN_data_out(5773),
        VN2CN2_bit => VN_data_out(5774),
        VN2CN3_bit => VN_data_out(5775),
        VN2CN4_bit => VN_data_out(5776),
        VN2CN5_bit => VN_data_out(5777),
        VN2CN0_sign => VN_sign_out(5772),
        VN2CN1_sign => VN_sign_out(5773),
        VN2CN2_sign => VN_sign_out(5774),
        VN2CN3_sign => VN_sign_out(5775),
        VN2CN4_sign => VN_sign_out(5776),
        VN2CN5_sign => VN_sign_out(5777),
        codeword => codeword(962),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN963 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5783 downto 5778),
        Din0 => VN963_in0,
        Din1 => VN963_in1,
        Din2 => VN963_in2,
        Din3 => VN963_in3,
        Din4 => VN963_in4,
        Din5 => VN963_in5,
        VN2CN0_bit => VN_data_out(5778),
        VN2CN1_bit => VN_data_out(5779),
        VN2CN2_bit => VN_data_out(5780),
        VN2CN3_bit => VN_data_out(5781),
        VN2CN4_bit => VN_data_out(5782),
        VN2CN5_bit => VN_data_out(5783),
        VN2CN0_sign => VN_sign_out(5778),
        VN2CN1_sign => VN_sign_out(5779),
        VN2CN2_sign => VN_sign_out(5780),
        VN2CN3_sign => VN_sign_out(5781),
        VN2CN4_sign => VN_sign_out(5782),
        VN2CN5_sign => VN_sign_out(5783),
        codeword => codeword(963),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN964 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5789 downto 5784),
        Din0 => VN964_in0,
        Din1 => VN964_in1,
        Din2 => VN964_in2,
        Din3 => VN964_in3,
        Din4 => VN964_in4,
        Din5 => VN964_in5,
        VN2CN0_bit => VN_data_out(5784),
        VN2CN1_bit => VN_data_out(5785),
        VN2CN2_bit => VN_data_out(5786),
        VN2CN3_bit => VN_data_out(5787),
        VN2CN4_bit => VN_data_out(5788),
        VN2CN5_bit => VN_data_out(5789),
        VN2CN0_sign => VN_sign_out(5784),
        VN2CN1_sign => VN_sign_out(5785),
        VN2CN2_sign => VN_sign_out(5786),
        VN2CN3_sign => VN_sign_out(5787),
        VN2CN4_sign => VN_sign_out(5788),
        VN2CN5_sign => VN_sign_out(5789),
        codeword => codeword(964),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN965 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5795 downto 5790),
        Din0 => VN965_in0,
        Din1 => VN965_in1,
        Din2 => VN965_in2,
        Din3 => VN965_in3,
        Din4 => VN965_in4,
        Din5 => VN965_in5,
        VN2CN0_bit => VN_data_out(5790),
        VN2CN1_bit => VN_data_out(5791),
        VN2CN2_bit => VN_data_out(5792),
        VN2CN3_bit => VN_data_out(5793),
        VN2CN4_bit => VN_data_out(5794),
        VN2CN5_bit => VN_data_out(5795),
        VN2CN0_sign => VN_sign_out(5790),
        VN2CN1_sign => VN_sign_out(5791),
        VN2CN2_sign => VN_sign_out(5792),
        VN2CN3_sign => VN_sign_out(5793),
        VN2CN4_sign => VN_sign_out(5794),
        VN2CN5_sign => VN_sign_out(5795),
        codeword => codeword(965),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN966 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5801 downto 5796),
        Din0 => VN966_in0,
        Din1 => VN966_in1,
        Din2 => VN966_in2,
        Din3 => VN966_in3,
        Din4 => VN966_in4,
        Din5 => VN966_in5,
        VN2CN0_bit => VN_data_out(5796),
        VN2CN1_bit => VN_data_out(5797),
        VN2CN2_bit => VN_data_out(5798),
        VN2CN3_bit => VN_data_out(5799),
        VN2CN4_bit => VN_data_out(5800),
        VN2CN5_bit => VN_data_out(5801),
        VN2CN0_sign => VN_sign_out(5796),
        VN2CN1_sign => VN_sign_out(5797),
        VN2CN2_sign => VN_sign_out(5798),
        VN2CN3_sign => VN_sign_out(5799),
        VN2CN4_sign => VN_sign_out(5800),
        VN2CN5_sign => VN_sign_out(5801),
        codeword => codeword(966),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN967 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5807 downto 5802),
        Din0 => VN967_in0,
        Din1 => VN967_in1,
        Din2 => VN967_in2,
        Din3 => VN967_in3,
        Din4 => VN967_in4,
        Din5 => VN967_in5,
        VN2CN0_bit => VN_data_out(5802),
        VN2CN1_bit => VN_data_out(5803),
        VN2CN2_bit => VN_data_out(5804),
        VN2CN3_bit => VN_data_out(5805),
        VN2CN4_bit => VN_data_out(5806),
        VN2CN5_bit => VN_data_out(5807),
        VN2CN0_sign => VN_sign_out(5802),
        VN2CN1_sign => VN_sign_out(5803),
        VN2CN2_sign => VN_sign_out(5804),
        VN2CN3_sign => VN_sign_out(5805),
        VN2CN4_sign => VN_sign_out(5806),
        VN2CN5_sign => VN_sign_out(5807),
        codeword => codeword(967),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN968 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5813 downto 5808),
        Din0 => VN968_in0,
        Din1 => VN968_in1,
        Din2 => VN968_in2,
        Din3 => VN968_in3,
        Din4 => VN968_in4,
        Din5 => VN968_in5,
        VN2CN0_bit => VN_data_out(5808),
        VN2CN1_bit => VN_data_out(5809),
        VN2CN2_bit => VN_data_out(5810),
        VN2CN3_bit => VN_data_out(5811),
        VN2CN4_bit => VN_data_out(5812),
        VN2CN5_bit => VN_data_out(5813),
        VN2CN0_sign => VN_sign_out(5808),
        VN2CN1_sign => VN_sign_out(5809),
        VN2CN2_sign => VN_sign_out(5810),
        VN2CN3_sign => VN_sign_out(5811),
        VN2CN4_sign => VN_sign_out(5812),
        VN2CN5_sign => VN_sign_out(5813),
        codeword => codeword(968),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN969 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5819 downto 5814),
        Din0 => VN969_in0,
        Din1 => VN969_in1,
        Din2 => VN969_in2,
        Din3 => VN969_in3,
        Din4 => VN969_in4,
        Din5 => VN969_in5,
        VN2CN0_bit => VN_data_out(5814),
        VN2CN1_bit => VN_data_out(5815),
        VN2CN2_bit => VN_data_out(5816),
        VN2CN3_bit => VN_data_out(5817),
        VN2CN4_bit => VN_data_out(5818),
        VN2CN5_bit => VN_data_out(5819),
        VN2CN0_sign => VN_sign_out(5814),
        VN2CN1_sign => VN_sign_out(5815),
        VN2CN2_sign => VN_sign_out(5816),
        VN2CN3_sign => VN_sign_out(5817),
        VN2CN4_sign => VN_sign_out(5818),
        VN2CN5_sign => VN_sign_out(5819),
        codeword => codeword(969),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN970 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5825 downto 5820),
        Din0 => VN970_in0,
        Din1 => VN970_in1,
        Din2 => VN970_in2,
        Din3 => VN970_in3,
        Din4 => VN970_in4,
        Din5 => VN970_in5,
        VN2CN0_bit => VN_data_out(5820),
        VN2CN1_bit => VN_data_out(5821),
        VN2CN2_bit => VN_data_out(5822),
        VN2CN3_bit => VN_data_out(5823),
        VN2CN4_bit => VN_data_out(5824),
        VN2CN5_bit => VN_data_out(5825),
        VN2CN0_sign => VN_sign_out(5820),
        VN2CN1_sign => VN_sign_out(5821),
        VN2CN2_sign => VN_sign_out(5822),
        VN2CN3_sign => VN_sign_out(5823),
        VN2CN4_sign => VN_sign_out(5824),
        VN2CN5_sign => VN_sign_out(5825),
        codeword => codeword(970),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN971 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5831 downto 5826),
        Din0 => VN971_in0,
        Din1 => VN971_in1,
        Din2 => VN971_in2,
        Din3 => VN971_in3,
        Din4 => VN971_in4,
        Din5 => VN971_in5,
        VN2CN0_bit => VN_data_out(5826),
        VN2CN1_bit => VN_data_out(5827),
        VN2CN2_bit => VN_data_out(5828),
        VN2CN3_bit => VN_data_out(5829),
        VN2CN4_bit => VN_data_out(5830),
        VN2CN5_bit => VN_data_out(5831),
        VN2CN0_sign => VN_sign_out(5826),
        VN2CN1_sign => VN_sign_out(5827),
        VN2CN2_sign => VN_sign_out(5828),
        VN2CN3_sign => VN_sign_out(5829),
        VN2CN4_sign => VN_sign_out(5830),
        VN2CN5_sign => VN_sign_out(5831),
        codeword => codeword(971),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN972 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5837 downto 5832),
        Din0 => VN972_in0,
        Din1 => VN972_in1,
        Din2 => VN972_in2,
        Din3 => VN972_in3,
        Din4 => VN972_in4,
        Din5 => VN972_in5,
        VN2CN0_bit => VN_data_out(5832),
        VN2CN1_bit => VN_data_out(5833),
        VN2CN2_bit => VN_data_out(5834),
        VN2CN3_bit => VN_data_out(5835),
        VN2CN4_bit => VN_data_out(5836),
        VN2CN5_bit => VN_data_out(5837),
        VN2CN0_sign => VN_sign_out(5832),
        VN2CN1_sign => VN_sign_out(5833),
        VN2CN2_sign => VN_sign_out(5834),
        VN2CN3_sign => VN_sign_out(5835),
        VN2CN4_sign => VN_sign_out(5836),
        VN2CN5_sign => VN_sign_out(5837),
        codeword => codeword(972),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN973 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5843 downto 5838),
        Din0 => VN973_in0,
        Din1 => VN973_in1,
        Din2 => VN973_in2,
        Din3 => VN973_in3,
        Din4 => VN973_in4,
        Din5 => VN973_in5,
        VN2CN0_bit => VN_data_out(5838),
        VN2CN1_bit => VN_data_out(5839),
        VN2CN2_bit => VN_data_out(5840),
        VN2CN3_bit => VN_data_out(5841),
        VN2CN4_bit => VN_data_out(5842),
        VN2CN5_bit => VN_data_out(5843),
        VN2CN0_sign => VN_sign_out(5838),
        VN2CN1_sign => VN_sign_out(5839),
        VN2CN2_sign => VN_sign_out(5840),
        VN2CN3_sign => VN_sign_out(5841),
        VN2CN4_sign => VN_sign_out(5842),
        VN2CN5_sign => VN_sign_out(5843),
        codeword => codeword(973),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN974 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5849 downto 5844),
        Din0 => VN974_in0,
        Din1 => VN974_in1,
        Din2 => VN974_in2,
        Din3 => VN974_in3,
        Din4 => VN974_in4,
        Din5 => VN974_in5,
        VN2CN0_bit => VN_data_out(5844),
        VN2CN1_bit => VN_data_out(5845),
        VN2CN2_bit => VN_data_out(5846),
        VN2CN3_bit => VN_data_out(5847),
        VN2CN4_bit => VN_data_out(5848),
        VN2CN5_bit => VN_data_out(5849),
        VN2CN0_sign => VN_sign_out(5844),
        VN2CN1_sign => VN_sign_out(5845),
        VN2CN2_sign => VN_sign_out(5846),
        VN2CN3_sign => VN_sign_out(5847),
        VN2CN4_sign => VN_sign_out(5848),
        VN2CN5_sign => VN_sign_out(5849),
        codeword => codeword(974),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN975 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5855 downto 5850),
        Din0 => VN975_in0,
        Din1 => VN975_in1,
        Din2 => VN975_in2,
        Din3 => VN975_in3,
        Din4 => VN975_in4,
        Din5 => VN975_in5,
        VN2CN0_bit => VN_data_out(5850),
        VN2CN1_bit => VN_data_out(5851),
        VN2CN2_bit => VN_data_out(5852),
        VN2CN3_bit => VN_data_out(5853),
        VN2CN4_bit => VN_data_out(5854),
        VN2CN5_bit => VN_data_out(5855),
        VN2CN0_sign => VN_sign_out(5850),
        VN2CN1_sign => VN_sign_out(5851),
        VN2CN2_sign => VN_sign_out(5852),
        VN2CN3_sign => VN_sign_out(5853),
        VN2CN4_sign => VN_sign_out(5854),
        VN2CN5_sign => VN_sign_out(5855),
        codeword => codeword(975),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN976 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5861 downto 5856),
        Din0 => VN976_in0,
        Din1 => VN976_in1,
        Din2 => VN976_in2,
        Din3 => VN976_in3,
        Din4 => VN976_in4,
        Din5 => VN976_in5,
        VN2CN0_bit => VN_data_out(5856),
        VN2CN1_bit => VN_data_out(5857),
        VN2CN2_bit => VN_data_out(5858),
        VN2CN3_bit => VN_data_out(5859),
        VN2CN4_bit => VN_data_out(5860),
        VN2CN5_bit => VN_data_out(5861),
        VN2CN0_sign => VN_sign_out(5856),
        VN2CN1_sign => VN_sign_out(5857),
        VN2CN2_sign => VN_sign_out(5858),
        VN2CN3_sign => VN_sign_out(5859),
        VN2CN4_sign => VN_sign_out(5860),
        VN2CN5_sign => VN_sign_out(5861),
        codeword => codeword(976),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN977 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5867 downto 5862),
        Din0 => VN977_in0,
        Din1 => VN977_in1,
        Din2 => VN977_in2,
        Din3 => VN977_in3,
        Din4 => VN977_in4,
        Din5 => VN977_in5,
        VN2CN0_bit => VN_data_out(5862),
        VN2CN1_bit => VN_data_out(5863),
        VN2CN2_bit => VN_data_out(5864),
        VN2CN3_bit => VN_data_out(5865),
        VN2CN4_bit => VN_data_out(5866),
        VN2CN5_bit => VN_data_out(5867),
        VN2CN0_sign => VN_sign_out(5862),
        VN2CN1_sign => VN_sign_out(5863),
        VN2CN2_sign => VN_sign_out(5864),
        VN2CN3_sign => VN_sign_out(5865),
        VN2CN4_sign => VN_sign_out(5866),
        VN2CN5_sign => VN_sign_out(5867),
        codeword => codeword(977),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN978 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5873 downto 5868),
        Din0 => VN978_in0,
        Din1 => VN978_in1,
        Din2 => VN978_in2,
        Din3 => VN978_in3,
        Din4 => VN978_in4,
        Din5 => VN978_in5,
        VN2CN0_bit => VN_data_out(5868),
        VN2CN1_bit => VN_data_out(5869),
        VN2CN2_bit => VN_data_out(5870),
        VN2CN3_bit => VN_data_out(5871),
        VN2CN4_bit => VN_data_out(5872),
        VN2CN5_bit => VN_data_out(5873),
        VN2CN0_sign => VN_sign_out(5868),
        VN2CN1_sign => VN_sign_out(5869),
        VN2CN2_sign => VN_sign_out(5870),
        VN2CN3_sign => VN_sign_out(5871),
        VN2CN4_sign => VN_sign_out(5872),
        VN2CN5_sign => VN_sign_out(5873),
        codeword => codeword(978),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN979 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5879 downto 5874),
        Din0 => VN979_in0,
        Din1 => VN979_in1,
        Din2 => VN979_in2,
        Din3 => VN979_in3,
        Din4 => VN979_in4,
        Din5 => VN979_in5,
        VN2CN0_bit => VN_data_out(5874),
        VN2CN1_bit => VN_data_out(5875),
        VN2CN2_bit => VN_data_out(5876),
        VN2CN3_bit => VN_data_out(5877),
        VN2CN4_bit => VN_data_out(5878),
        VN2CN5_bit => VN_data_out(5879),
        VN2CN0_sign => VN_sign_out(5874),
        VN2CN1_sign => VN_sign_out(5875),
        VN2CN2_sign => VN_sign_out(5876),
        VN2CN3_sign => VN_sign_out(5877),
        VN2CN4_sign => VN_sign_out(5878),
        VN2CN5_sign => VN_sign_out(5879),
        codeword => codeword(979),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN980 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5885 downto 5880),
        Din0 => VN980_in0,
        Din1 => VN980_in1,
        Din2 => VN980_in2,
        Din3 => VN980_in3,
        Din4 => VN980_in4,
        Din5 => VN980_in5,
        VN2CN0_bit => VN_data_out(5880),
        VN2CN1_bit => VN_data_out(5881),
        VN2CN2_bit => VN_data_out(5882),
        VN2CN3_bit => VN_data_out(5883),
        VN2CN4_bit => VN_data_out(5884),
        VN2CN5_bit => VN_data_out(5885),
        VN2CN0_sign => VN_sign_out(5880),
        VN2CN1_sign => VN_sign_out(5881),
        VN2CN2_sign => VN_sign_out(5882),
        VN2CN3_sign => VN_sign_out(5883),
        VN2CN4_sign => VN_sign_out(5884),
        VN2CN5_sign => VN_sign_out(5885),
        codeword => codeword(980),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN981 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5891 downto 5886),
        Din0 => VN981_in0,
        Din1 => VN981_in1,
        Din2 => VN981_in2,
        Din3 => VN981_in3,
        Din4 => VN981_in4,
        Din5 => VN981_in5,
        VN2CN0_bit => VN_data_out(5886),
        VN2CN1_bit => VN_data_out(5887),
        VN2CN2_bit => VN_data_out(5888),
        VN2CN3_bit => VN_data_out(5889),
        VN2CN4_bit => VN_data_out(5890),
        VN2CN5_bit => VN_data_out(5891),
        VN2CN0_sign => VN_sign_out(5886),
        VN2CN1_sign => VN_sign_out(5887),
        VN2CN2_sign => VN_sign_out(5888),
        VN2CN3_sign => VN_sign_out(5889),
        VN2CN4_sign => VN_sign_out(5890),
        VN2CN5_sign => VN_sign_out(5891),
        codeword => codeword(981),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN982 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5897 downto 5892),
        Din0 => VN982_in0,
        Din1 => VN982_in1,
        Din2 => VN982_in2,
        Din3 => VN982_in3,
        Din4 => VN982_in4,
        Din5 => VN982_in5,
        VN2CN0_bit => VN_data_out(5892),
        VN2CN1_bit => VN_data_out(5893),
        VN2CN2_bit => VN_data_out(5894),
        VN2CN3_bit => VN_data_out(5895),
        VN2CN4_bit => VN_data_out(5896),
        VN2CN5_bit => VN_data_out(5897),
        VN2CN0_sign => VN_sign_out(5892),
        VN2CN1_sign => VN_sign_out(5893),
        VN2CN2_sign => VN_sign_out(5894),
        VN2CN3_sign => VN_sign_out(5895),
        VN2CN4_sign => VN_sign_out(5896),
        VN2CN5_sign => VN_sign_out(5897),
        codeword => codeword(982),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN983 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5903 downto 5898),
        Din0 => VN983_in0,
        Din1 => VN983_in1,
        Din2 => VN983_in2,
        Din3 => VN983_in3,
        Din4 => VN983_in4,
        Din5 => VN983_in5,
        VN2CN0_bit => VN_data_out(5898),
        VN2CN1_bit => VN_data_out(5899),
        VN2CN2_bit => VN_data_out(5900),
        VN2CN3_bit => VN_data_out(5901),
        VN2CN4_bit => VN_data_out(5902),
        VN2CN5_bit => VN_data_out(5903),
        VN2CN0_sign => VN_sign_out(5898),
        VN2CN1_sign => VN_sign_out(5899),
        VN2CN2_sign => VN_sign_out(5900),
        VN2CN3_sign => VN_sign_out(5901),
        VN2CN4_sign => VN_sign_out(5902),
        VN2CN5_sign => VN_sign_out(5903),
        codeword => codeword(983),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN984 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5909 downto 5904),
        Din0 => VN984_in0,
        Din1 => VN984_in1,
        Din2 => VN984_in2,
        Din3 => VN984_in3,
        Din4 => VN984_in4,
        Din5 => VN984_in5,
        VN2CN0_bit => VN_data_out(5904),
        VN2CN1_bit => VN_data_out(5905),
        VN2CN2_bit => VN_data_out(5906),
        VN2CN3_bit => VN_data_out(5907),
        VN2CN4_bit => VN_data_out(5908),
        VN2CN5_bit => VN_data_out(5909),
        VN2CN0_sign => VN_sign_out(5904),
        VN2CN1_sign => VN_sign_out(5905),
        VN2CN2_sign => VN_sign_out(5906),
        VN2CN3_sign => VN_sign_out(5907),
        VN2CN4_sign => VN_sign_out(5908),
        VN2CN5_sign => VN_sign_out(5909),
        codeword => codeword(984),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN985 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5915 downto 5910),
        Din0 => VN985_in0,
        Din1 => VN985_in1,
        Din2 => VN985_in2,
        Din3 => VN985_in3,
        Din4 => VN985_in4,
        Din5 => VN985_in5,
        VN2CN0_bit => VN_data_out(5910),
        VN2CN1_bit => VN_data_out(5911),
        VN2CN2_bit => VN_data_out(5912),
        VN2CN3_bit => VN_data_out(5913),
        VN2CN4_bit => VN_data_out(5914),
        VN2CN5_bit => VN_data_out(5915),
        VN2CN0_sign => VN_sign_out(5910),
        VN2CN1_sign => VN_sign_out(5911),
        VN2CN2_sign => VN_sign_out(5912),
        VN2CN3_sign => VN_sign_out(5913),
        VN2CN4_sign => VN_sign_out(5914),
        VN2CN5_sign => VN_sign_out(5915),
        codeword => codeword(985),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN986 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5921 downto 5916),
        Din0 => VN986_in0,
        Din1 => VN986_in1,
        Din2 => VN986_in2,
        Din3 => VN986_in3,
        Din4 => VN986_in4,
        Din5 => VN986_in5,
        VN2CN0_bit => VN_data_out(5916),
        VN2CN1_bit => VN_data_out(5917),
        VN2CN2_bit => VN_data_out(5918),
        VN2CN3_bit => VN_data_out(5919),
        VN2CN4_bit => VN_data_out(5920),
        VN2CN5_bit => VN_data_out(5921),
        VN2CN0_sign => VN_sign_out(5916),
        VN2CN1_sign => VN_sign_out(5917),
        VN2CN2_sign => VN_sign_out(5918),
        VN2CN3_sign => VN_sign_out(5919),
        VN2CN4_sign => VN_sign_out(5920),
        VN2CN5_sign => VN_sign_out(5921),
        codeword => codeword(986),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN987 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5927 downto 5922),
        Din0 => VN987_in0,
        Din1 => VN987_in1,
        Din2 => VN987_in2,
        Din3 => VN987_in3,
        Din4 => VN987_in4,
        Din5 => VN987_in5,
        VN2CN0_bit => VN_data_out(5922),
        VN2CN1_bit => VN_data_out(5923),
        VN2CN2_bit => VN_data_out(5924),
        VN2CN3_bit => VN_data_out(5925),
        VN2CN4_bit => VN_data_out(5926),
        VN2CN5_bit => VN_data_out(5927),
        VN2CN0_sign => VN_sign_out(5922),
        VN2CN1_sign => VN_sign_out(5923),
        VN2CN2_sign => VN_sign_out(5924),
        VN2CN3_sign => VN_sign_out(5925),
        VN2CN4_sign => VN_sign_out(5926),
        VN2CN5_sign => VN_sign_out(5927),
        codeword => codeword(987),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN988 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5933 downto 5928),
        Din0 => VN988_in0,
        Din1 => VN988_in1,
        Din2 => VN988_in2,
        Din3 => VN988_in3,
        Din4 => VN988_in4,
        Din5 => VN988_in5,
        VN2CN0_bit => VN_data_out(5928),
        VN2CN1_bit => VN_data_out(5929),
        VN2CN2_bit => VN_data_out(5930),
        VN2CN3_bit => VN_data_out(5931),
        VN2CN4_bit => VN_data_out(5932),
        VN2CN5_bit => VN_data_out(5933),
        VN2CN0_sign => VN_sign_out(5928),
        VN2CN1_sign => VN_sign_out(5929),
        VN2CN2_sign => VN_sign_out(5930),
        VN2CN3_sign => VN_sign_out(5931),
        VN2CN4_sign => VN_sign_out(5932),
        VN2CN5_sign => VN_sign_out(5933),
        codeword => codeword(988),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN989 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5939 downto 5934),
        Din0 => VN989_in0,
        Din1 => VN989_in1,
        Din2 => VN989_in2,
        Din3 => VN989_in3,
        Din4 => VN989_in4,
        Din5 => VN989_in5,
        VN2CN0_bit => VN_data_out(5934),
        VN2CN1_bit => VN_data_out(5935),
        VN2CN2_bit => VN_data_out(5936),
        VN2CN3_bit => VN_data_out(5937),
        VN2CN4_bit => VN_data_out(5938),
        VN2CN5_bit => VN_data_out(5939),
        VN2CN0_sign => VN_sign_out(5934),
        VN2CN1_sign => VN_sign_out(5935),
        VN2CN2_sign => VN_sign_out(5936),
        VN2CN3_sign => VN_sign_out(5937),
        VN2CN4_sign => VN_sign_out(5938),
        VN2CN5_sign => VN_sign_out(5939),
        codeword => codeword(989),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN990 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5945 downto 5940),
        Din0 => VN990_in0,
        Din1 => VN990_in1,
        Din2 => VN990_in2,
        Din3 => VN990_in3,
        Din4 => VN990_in4,
        Din5 => VN990_in5,
        VN2CN0_bit => VN_data_out(5940),
        VN2CN1_bit => VN_data_out(5941),
        VN2CN2_bit => VN_data_out(5942),
        VN2CN3_bit => VN_data_out(5943),
        VN2CN4_bit => VN_data_out(5944),
        VN2CN5_bit => VN_data_out(5945),
        VN2CN0_sign => VN_sign_out(5940),
        VN2CN1_sign => VN_sign_out(5941),
        VN2CN2_sign => VN_sign_out(5942),
        VN2CN3_sign => VN_sign_out(5943),
        VN2CN4_sign => VN_sign_out(5944),
        VN2CN5_sign => VN_sign_out(5945),
        codeword => codeword(990),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN991 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5951 downto 5946),
        Din0 => VN991_in0,
        Din1 => VN991_in1,
        Din2 => VN991_in2,
        Din3 => VN991_in3,
        Din4 => VN991_in4,
        Din5 => VN991_in5,
        VN2CN0_bit => VN_data_out(5946),
        VN2CN1_bit => VN_data_out(5947),
        VN2CN2_bit => VN_data_out(5948),
        VN2CN3_bit => VN_data_out(5949),
        VN2CN4_bit => VN_data_out(5950),
        VN2CN5_bit => VN_data_out(5951),
        VN2CN0_sign => VN_sign_out(5946),
        VN2CN1_sign => VN_sign_out(5947),
        VN2CN2_sign => VN_sign_out(5948),
        VN2CN3_sign => VN_sign_out(5949),
        VN2CN4_sign => VN_sign_out(5950),
        VN2CN5_sign => VN_sign_out(5951),
        codeword => codeword(991),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN992 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5957 downto 5952),
        Din0 => VN992_in0,
        Din1 => VN992_in1,
        Din2 => VN992_in2,
        Din3 => VN992_in3,
        Din4 => VN992_in4,
        Din5 => VN992_in5,
        VN2CN0_bit => VN_data_out(5952),
        VN2CN1_bit => VN_data_out(5953),
        VN2CN2_bit => VN_data_out(5954),
        VN2CN3_bit => VN_data_out(5955),
        VN2CN4_bit => VN_data_out(5956),
        VN2CN5_bit => VN_data_out(5957),
        VN2CN0_sign => VN_sign_out(5952),
        VN2CN1_sign => VN_sign_out(5953),
        VN2CN2_sign => VN_sign_out(5954),
        VN2CN3_sign => VN_sign_out(5955),
        VN2CN4_sign => VN_sign_out(5956),
        VN2CN5_sign => VN_sign_out(5957),
        codeword => codeword(992),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN993 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5963 downto 5958),
        Din0 => VN993_in0,
        Din1 => VN993_in1,
        Din2 => VN993_in2,
        Din3 => VN993_in3,
        Din4 => VN993_in4,
        Din5 => VN993_in5,
        VN2CN0_bit => VN_data_out(5958),
        VN2CN1_bit => VN_data_out(5959),
        VN2CN2_bit => VN_data_out(5960),
        VN2CN3_bit => VN_data_out(5961),
        VN2CN4_bit => VN_data_out(5962),
        VN2CN5_bit => VN_data_out(5963),
        VN2CN0_sign => VN_sign_out(5958),
        VN2CN1_sign => VN_sign_out(5959),
        VN2CN2_sign => VN_sign_out(5960),
        VN2CN3_sign => VN_sign_out(5961),
        VN2CN4_sign => VN_sign_out(5962),
        VN2CN5_sign => VN_sign_out(5963),
        codeword => codeword(993),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN994 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5969 downto 5964),
        Din0 => VN994_in0,
        Din1 => VN994_in1,
        Din2 => VN994_in2,
        Din3 => VN994_in3,
        Din4 => VN994_in4,
        Din5 => VN994_in5,
        VN2CN0_bit => VN_data_out(5964),
        VN2CN1_bit => VN_data_out(5965),
        VN2CN2_bit => VN_data_out(5966),
        VN2CN3_bit => VN_data_out(5967),
        VN2CN4_bit => VN_data_out(5968),
        VN2CN5_bit => VN_data_out(5969),
        VN2CN0_sign => VN_sign_out(5964),
        VN2CN1_sign => VN_sign_out(5965),
        VN2CN2_sign => VN_sign_out(5966),
        VN2CN3_sign => VN_sign_out(5967),
        VN2CN4_sign => VN_sign_out(5968),
        VN2CN5_sign => VN_sign_out(5969),
        codeword => codeword(994),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN995 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5975 downto 5970),
        Din0 => VN995_in0,
        Din1 => VN995_in1,
        Din2 => VN995_in2,
        Din3 => VN995_in3,
        Din4 => VN995_in4,
        Din5 => VN995_in5,
        VN2CN0_bit => VN_data_out(5970),
        VN2CN1_bit => VN_data_out(5971),
        VN2CN2_bit => VN_data_out(5972),
        VN2CN3_bit => VN_data_out(5973),
        VN2CN4_bit => VN_data_out(5974),
        VN2CN5_bit => VN_data_out(5975),
        VN2CN0_sign => VN_sign_out(5970),
        VN2CN1_sign => VN_sign_out(5971),
        VN2CN2_sign => VN_sign_out(5972),
        VN2CN3_sign => VN_sign_out(5973),
        VN2CN4_sign => VN_sign_out(5974),
        VN2CN5_sign => VN_sign_out(5975),
        codeword => codeword(995),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN996 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5981 downto 5976),
        Din0 => VN996_in0,
        Din1 => VN996_in1,
        Din2 => VN996_in2,
        Din3 => VN996_in3,
        Din4 => VN996_in4,
        Din5 => VN996_in5,
        VN2CN0_bit => VN_data_out(5976),
        VN2CN1_bit => VN_data_out(5977),
        VN2CN2_bit => VN_data_out(5978),
        VN2CN3_bit => VN_data_out(5979),
        VN2CN4_bit => VN_data_out(5980),
        VN2CN5_bit => VN_data_out(5981),
        VN2CN0_sign => VN_sign_out(5976),
        VN2CN1_sign => VN_sign_out(5977),
        VN2CN2_sign => VN_sign_out(5978),
        VN2CN3_sign => VN_sign_out(5979),
        VN2CN4_sign => VN_sign_out(5980),
        VN2CN5_sign => VN_sign_out(5981),
        codeword => codeword(996),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN997 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5987 downto 5982),
        Din0 => VN997_in0,
        Din1 => VN997_in1,
        Din2 => VN997_in2,
        Din3 => VN997_in3,
        Din4 => VN997_in4,
        Din5 => VN997_in5,
        VN2CN0_bit => VN_data_out(5982),
        VN2CN1_bit => VN_data_out(5983),
        VN2CN2_bit => VN_data_out(5984),
        VN2CN3_bit => VN_data_out(5985),
        VN2CN4_bit => VN_data_out(5986),
        VN2CN5_bit => VN_data_out(5987),
        VN2CN0_sign => VN_sign_out(5982),
        VN2CN1_sign => VN_sign_out(5983),
        VN2CN2_sign => VN_sign_out(5984),
        VN2CN3_sign => VN_sign_out(5985),
        VN2CN4_sign => VN_sign_out(5986),
        VN2CN5_sign => VN_sign_out(5987),
        codeword => codeword(997),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN998 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5993 downto 5988),
        Din0 => VN998_in0,
        Din1 => VN998_in1,
        Din2 => VN998_in2,
        Din3 => VN998_in3,
        Din4 => VN998_in4,
        Din5 => VN998_in5,
        VN2CN0_bit => VN_data_out(5988),
        VN2CN1_bit => VN_data_out(5989),
        VN2CN2_bit => VN_data_out(5990),
        VN2CN3_bit => VN_data_out(5991),
        VN2CN4_bit => VN_data_out(5992),
        VN2CN5_bit => VN_data_out(5993),
        VN2CN0_sign => VN_sign_out(5988),
        VN2CN1_sign => VN_sign_out(5989),
        VN2CN2_sign => VN_sign_out(5990),
        VN2CN3_sign => VN_sign_out(5991),
        VN2CN4_sign => VN_sign_out(5992),
        VN2CN5_sign => VN_sign_out(5993),
        codeword => codeword(998),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN999 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(5999 downto 5994),
        Din0 => VN999_in0,
        Din1 => VN999_in1,
        Din2 => VN999_in2,
        Din3 => VN999_in3,
        Din4 => VN999_in4,
        Din5 => VN999_in5,
        VN2CN0_bit => VN_data_out(5994),
        VN2CN1_bit => VN_data_out(5995),
        VN2CN2_bit => VN_data_out(5996),
        VN2CN3_bit => VN_data_out(5997),
        VN2CN4_bit => VN_data_out(5998),
        VN2CN5_bit => VN_data_out(5999),
        VN2CN0_sign => VN_sign_out(5994),
        VN2CN1_sign => VN_sign_out(5995),
        VN2CN2_sign => VN_sign_out(5996),
        VN2CN3_sign => VN_sign_out(5997),
        VN2CN4_sign => VN_sign_out(5998),
        VN2CN5_sign => VN_sign_out(5999),
        codeword => codeword(999),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1000 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6005 downto 6000),
        Din0 => VN1000_in0,
        Din1 => VN1000_in1,
        Din2 => VN1000_in2,
        Din3 => VN1000_in3,
        Din4 => VN1000_in4,
        Din5 => VN1000_in5,
        VN2CN0_bit => VN_data_out(6000),
        VN2CN1_bit => VN_data_out(6001),
        VN2CN2_bit => VN_data_out(6002),
        VN2CN3_bit => VN_data_out(6003),
        VN2CN4_bit => VN_data_out(6004),
        VN2CN5_bit => VN_data_out(6005),
        VN2CN0_sign => VN_sign_out(6000),
        VN2CN1_sign => VN_sign_out(6001),
        VN2CN2_sign => VN_sign_out(6002),
        VN2CN3_sign => VN_sign_out(6003),
        VN2CN4_sign => VN_sign_out(6004),
        VN2CN5_sign => VN_sign_out(6005),
        codeword => codeword(1000),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1001 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6011 downto 6006),
        Din0 => VN1001_in0,
        Din1 => VN1001_in1,
        Din2 => VN1001_in2,
        Din3 => VN1001_in3,
        Din4 => VN1001_in4,
        Din5 => VN1001_in5,
        VN2CN0_bit => VN_data_out(6006),
        VN2CN1_bit => VN_data_out(6007),
        VN2CN2_bit => VN_data_out(6008),
        VN2CN3_bit => VN_data_out(6009),
        VN2CN4_bit => VN_data_out(6010),
        VN2CN5_bit => VN_data_out(6011),
        VN2CN0_sign => VN_sign_out(6006),
        VN2CN1_sign => VN_sign_out(6007),
        VN2CN2_sign => VN_sign_out(6008),
        VN2CN3_sign => VN_sign_out(6009),
        VN2CN4_sign => VN_sign_out(6010),
        VN2CN5_sign => VN_sign_out(6011),
        codeword => codeword(1001),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1002 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6017 downto 6012),
        Din0 => VN1002_in0,
        Din1 => VN1002_in1,
        Din2 => VN1002_in2,
        Din3 => VN1002_in3,
        Din4 => VN1002_in4,
        Din5 => VN1002_in5,
        VN2CN0_bit => VN_data_out(6012),
        VN2CN1_bit => VN_data_out(6013),
        VN2CN2_bit => VN_data_out(6014),
        VN2CN3_bit => VN_data_out(6015),
        VN2CN4_bit => VN_data_out(6016),
        VN2CN5_bit => VN_data_out(6017),
        VN2CN0_sign => VN_sign_out(6012),
        VN2CN1_sign => VN_sign_out(6013),
        VN2CN2_sign => VN_sign_out(6014),
        VN2CN3_sign => VN_sign_out(6015),
        VN2CN4_sign => VN_sign_out(6016),
        VN2CN5_sign => VN_sign_out(6017),
        codeword => codeword(1002),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1003 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6023 downto 6018),
        Din0 => VN1003_in0,
        Din1 => VN1003_in1,
        Din2 => VN1003_in2,
        Din3 => VN1003_in3,
        Din4 => VN1003_in4,
        Din5 => VN1003_in5,
        VN2CN0_bit => VN_data_out(6018),
        VN2CN1_bit => VN_data_out(6019),
        VN2CN2_bit => VN_data_out(6020),
        VN2CN3_bit => VN_data_out(6021),
        VN2CN4_bit => VN_data_out(6022),
        VN2CN5_bit => VN_data_out(6023),
        VN2CN0_sign => VN_sign_out(6018),
        VN2CN1_sign => VN_sign_out(6019),
        VN2CN2_sign => VN_sign_out(6020),
        VN2CN3_sign => VN_sign_out(6021),
        VN2CN4_sign => VN_sign_out(6022),
        VN2CN5_sign => VN_sign_out(6023),
        codeword => codeword(1003),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1004 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6029 downto 6024),
        Din0 => VN1004_in0,
        Din1 => VN1004_in1,
        Din2 => VN1004_in2,
        Din3 => VN1004_in3,
        Din4 => VN1004_in4,
        Din5 => VN1004_in5,
        VN2CN0_bit => VN_data_out(6024),
        VN2CN1_bit => VN_data_out(6025),
        VN2CN2_bit => VN_data_out(6026),
        VN2CN3_bit => VN_data_out(6027),
        VN2CN4_bit => VN_data_out(6028),
        VN2CN5_bit => VN_data_out(6029),
        VN2CN0_sign => VN_sign_out(6024),
        VN2CN1_sign => VN_sign_out(6025),
        VN2CN2_sign => VN_sign_out(6026),
        VN2CN3_sign => VN_sign_out(6027),
        VN2CN4_sign => VN_sign_out(6028),
        VN2CN5_sign => VN_sign_out(6029),
        codeword => codeword(1004),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1005 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6035 downto 6030),
        Din0 => VN1005_in0,
        Din1 => VN1005_in1,
        Din2 => VN1005_in2,
        Din3 => VN1005_in3,
        Din4 => VN1005_in4,
        Din5 => VN1005_in5,
        VN2CN0_bit => VN_data_out(6030),
        VN2CN1_bit => VN_data_out(6031),
        VN2CN2_bit => VN_data_out(6032),
        VN2CN3_bit => VN_data_out(6033),
        VN2CN4_bit => VN_data_out(6034),
        VN2CN5_bit => VN_data_out(6035),
        VN2CN0_sign => VN_sign_out(6030),
        VN2CN1_sign => VN_sign_out(6031),
        VN2CN2_sign => VN_sign_out(6032),
        VN2CN3_sign => VN_sign_out(6033),
        VN2CN4_sign => VN_sign_out(6034),
        VN2CN5_sign => VN_sign_out(6035),
        codeword => codeword(1005),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1006 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6041 downto 6036),
        Din0 => VN1006_in0,
        Din1 => VN1006_in1,
        Din2 => VN1006_in2,
        Din3 => VN1006_in3,
        Din4 => VN1006_in4,
        Din5 => VN1006_in5,
        VN2CN0_bit => VN_data_out(6036),
        VN2CN1_bit => VN_data_out(6037),
        VN2CN2_bit => VN_data_out(6038),
        VN2CN3_bit => VN_data_out(6039),
        VN2CN4_bit => VN_data_out(6040),
        VN2CN5_bit => VN_data_out(6041),
        VN2CN0_sign => VN_sign_out(6036),
        VN2CN1_sign => VN_sign_out(6037),
        VN2CN2_sign => VN_sign_out(6038),
        VN2CN3_sign => VN_sign_out(6039),
        VN2CN4_sign => VN_sign_out(6040),
        VN2CN5_sign => VN_sign_out(6041),
        codeword => codeword(1006),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1007 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6047 downto 6042),
        Din0 => VN1007_in0,
        Din1 => VN1007_in1,
        Din2 => VN1007_in2,
        Din3 => VN1007_in3,
        Din4 => VN1007_in4,
        Din5 => VN1007_in5,
        VN2CN0_bit => VN_data_out(6042),
        VN2CN1_bit => VN_data_out(6043),
        VN2CN2_bit => VN_data_out(6044),
        VN2CN3_bit => VN_data_out(6045),
        VN2CN4_bit => VN_data_out(6046),
        VN2CN5_bit => VN_data_out(6047),
        VN2CN0_sign => VN_sign_out(6042),
        VN2CN1_sign => VN_sign_out(6043),
        VN2CN2_sign => VN_sign_out(6044),
        VN2CN3_sign => VN_sign_out(6045),
        VN2CN4_sign => VN_sign_out(6046),
        VN2CN5_sign => VN_sign_out(6047),
        codeword => codeword(1007),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1008 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6053 downto 6048),
        Din0 => VN1008_in0,
        Din1 => VN1008_in1,
        Din2 => VN1008_in2,
        Din3 => VN1008_in3,
        Din4 => VN1008_in4,
        Din5 => VN1008_in5,
        VN2CN0_bit => VN_data_out(6048),
        VN2CN1_bit => VN_data_out(6049),
        VN2CN2_bit => VN_data_out(6050),
        VN2CN3_bit => VN_data_out(6051),
        VN2CN4_bit => VN_data_out(6052),
        VN2CN5_bit => VN_data_out(6053),
        VN2CN0_sign => VN_sign_out(6048),
        VN2CN1_sign => VN_sign_out(6049),
        VN2CN2_sign => VN_sign_out(6050),
        VN2CN3_sign => VN_sign_out(6051),
        VN2CN4_sign => VN_sign_out(6052),
        VN2CN5_sign => VN_sign_out(6053),
        codeword => codeword(1008),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1009 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6059 downto 6054),
        Din0 => VN1009_in0,
        Din1 => VN1009_in1,
        Din2 => VN1009_in2,
        Din3 => VN1009_in3,
        Din4 => VN1009_in4,
        Din5 => VN1009_in5,
        VN2CN0_bit => VN_data_out(6054),
        VN2CN1_bit => VN_data_out(6055),
        VN2CN2_bit => VN_data_out(6056),
        VN2CN3_bit => VN_data_out(6057),
        VN2CN4_bit => VN_data_out(6058),
        VN2CN5_bit => VN_data_out(6059),
        VN2CN0_sign => VN_sign_out(6054),
        VN2CN1_sign => VN_sign_out(6055),
        VN2CN2_sign => VN_sign_out(6056),
        VN2CN3_sign => VN_sign_out(6057),
        VN2CN4_sign => VN_sign_out(6058),
        VN2CN5_sign => VN_sign_out(6059),
        codeword => codeword(1009),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1010 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6065 downto 6060),
        Din0 => VN1010_in0,
        Din1 => VN1010_in1,
        Din2 => VN1010_in2,
        Din3 => VN1010_in3,
        Din4 => VN1010_in4,
        Din5 => VN1010_in5,
        VN2CN0_bit => VN_data_out(6060),
        VN2CN1_bit => VN_data_out(6061),
        VN2CN2_bit => VN_data_out(6062),
        VN2CN3_bit => VN_data_out(6063),
        VN2CN4_bit => VN_data_out(6064),
        VN2CN5_bit => VN_data_out(6065),
        VN2CN0_sign => VN_sign_out(6060),
        VN2CN1_sign => VN_sign_out(6061),
        VN2CN2_sign => VN_sign_out(6062),
        VN2CN3_sign => VN_sign_out(6063),
        VN2CN4_sign => VN_sign_out(6064),
        VN2CN5_sign => VN_sign_out(6065),
        codeword => codeword(1010),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1011 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6071 downto 6066),
        Din0 => VN1011_in0,
        Din1 => VN1011_in1,
        Din2 => VN1011_in2,
        Din3 => VN1011_in3,
        Din4 => VN1011_in4,
        Din5 => VN1011_in5,
        VN2CN0_bit => VN_data_out(6066),
        VN2CN1_bit => VN_data_out(6067),
        VN2CN2_bit => VN_data_out(6068),
        VN2CN3_bit => VN_data_out(6069),
        VN2CN4_bit => VN_data_out(6070),
        VN2CN5_bit => VN_data_out(6071),
        VN2CN0_sign => VN_sign_out(6066),
        VN2CN1_sign => VN_sign_out(6067),
        VN2CN2_sign => VN_sign_out(6068),
        VN2CN3_sign => VN_sign_out(6069),
        VN2CN4_sign => VN_sign_out(6070),
        VN2CN5_sign => VN_sign_out(6071),
        codeword => codeword(1011),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1012 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6077 downto 6072),
        Din0 => VN1012_in0,
        Din1 => VN1012_in1,
        Din2 => VN1012_in2,
        Din3 => VN1012_in3,
        Din4 => VN1012_in4,
        Din5 => VN1012_in5,
        VN2CN0_bit => VN_data_out(6072),
        VN2CN1_bit => VN_data_out(6073),
        VN2CN2_bit => VN_data_out(6074),
        VN2CN3_bit => VN_data_out(6075),
        VN2CN4_bit => VN_data_out(6076),
        VN2CN5_bit => VN_data_out(6077),
        VN2CN0_sign => VN_sign_out(6072),
        VN2CN1_sign => VN_sign_out(6073),
        VN2CN2_sign => VN_sign_out(6074),
        VN2CN3_sign => VN_sign_out(6075),
        VN2CN4_sign => VN_sign_out(6076),
        VN2CN5_sign => VN_sign_out(6077),
        codeword => codeword(1012),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1013 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6083 downto 6078),
        Din0 => VN1013_in0,
        Din1 => VN1013_in1,
        Din2 => VN1013_in2,
        Din3 => VN1013_in3,
        Din4 => VN1013_in4,
        Din5 => VN1013_in5,
        VN2CN0_bit => VN_data_out(6078),
        VN2CN1_bit => VN_data_out(6079),
        VN2CN2_bit => VN_data_out(6080),
        VN2CN3_bit => VN_data_out(6081),
        VN2CN4_bit => VN_data_out(6082),
        VN2CN5_bit => VN_data_out(6083),
        VN2CN0_sign => VN_sign_out(6078),
        VN2CN1_sign => VN_sign_out(6079),
        VN2CN2_sign => VN_sign_out(6080),
        VN2CN3_sign => VN_sign_out(6081),
        VN2CN4_sign => VN_sign_out(6082),
        VN2CN5_sign => VN_sign_out(6083),
        codeword => codeword(1013),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1014 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6089 downto 6084),
        Din0 => VN1014_in0,
        Din1 => VN1014_in1,
        Din2 => VN1014_in2,
        Din3 => VN1014_in3,
        Din4 => VN1014_in4,
        Din5 => VN1014_in5,
        VN2CN0_bit => VN_data_out(6084),
        VN2CN1_bit => VN_data_out(6085),
        VN2CN2_bit => VN_data_out(6086),
        VN2CN3_bit => VN_data_out(6087),
        VN2CN4_bit => VN_data_out(6088),
        VN2CN5_bit => VN_data_out(6089),
        VN2CN0_sign => VN_sign_out(6084),
        VN2CN1_sign => VN_sign_out(6085),
        VN2CN2_sign => VN_sign_out(6086),
        VN2CN3_sign => VN_sign_out(6087),
        VN2CN4_sign => VN_sign_out(6088),
        VN2CN5_sign => VN_sign_out(6089),
        codeword => codeword(1014),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1015 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6095 downto 6090),
        Din0 => VN1015_in0,
        Din1 => VN1015_in1,
        Din2 => VN1015_in2,
        Din3 => VN1015_in3,
        Din4 => VN1015_in4,
        Din5 => VN1015_in5,
        VN2CN0_bit => VN_data_out(6090),
        VN2CN1_bit => VN_data_out(6091),
        VN2CN2_bit => VN_data_out(6092),
        VN2CN3_bit => VN_data_out(6093),
        VN2CN4_bit => VN_data_out(6094),
        VN2CN5_bit => VN_data_out(6095),
        VN2CN0_sign => VN_sign_out(6090),
        VN2CN1_sign => VN_sign_out(6091),
        VN2CN2_sign => VN_sign_out(6092),
        VN2CN3_sign => VN_sign_out(6093),
        VN2CN4_sign => VN_sign_out(6094),
        VN2CN5_sign => VN_sign_out(6095),
        codeword => codeword(1015),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1016 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6101 downto 6096),
        Din0 => VN1016_in0,
        Din1 => VN1016_in1,
        Din2 => VN1016_in2,
        Din3 => VN1016_in3,
        Din4 => VN1016_in4,
        Din5 => VN1016_in5,
        VN2CN0_bit => VN_data_out(6096),
        VN2CN1_bit => VN_data_out(6097),
        VN2CN2_bit => VN_data_out(6098),
        VN2CN3_bit => VN_data_out(6099),
        VN2CN4_bit => VN_data_out(6100),
        VN2CN5_bit => VN_data_out(6101),
        VN2CN0_sign => VN_sign_out(6096),
        VN2CN1_sign => VN_sign_out(6097),
        VN2CN2_sign => VN_sign_out(6098),
        VN2CN3_sign => VN_sign_out(6099),
        VN2CN4_sign => VN_sign_out(6100),
        VN2CN5_sign => VN_sign_out(6101),
        codeword => codeword(1016),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1017 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6107 downto 6102),
        Din0 => VN1017_in0,
        Din1 => VN1017_in1,
        Din2 => VN1017_in2,
        Din3 => VN1017_in3,
        Din4 => VN1017_in4,
        Din5 => VN1017_in5,
        VN2CN0_bit => VN_data_out(6102),
        VN2CN1_bit => VN_data_out(6103),
        VN2CN2_bit => VN_data_out(6104),
        VN2CN3_bit => VN_data_out(6105),
        VN2CN4_bit => VN_data_out(6106),
        VN2CN5_bit => VN_data_out(6107),
        VN2CN0_sign => VN_sign_out(6102),
        VN2CN1_sign => VN_sign_out(6103),
        VN2CN2_sign => VN_sign_out(6104),
        VN2CN3_sign => VN_sign_out(6105),
        VN2CN4_sign => VN_sign_out(6106),
        VN2CN5_sign => VN_sign_out(6107),
        codeword => codeword(1017),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1018 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6113 downto 6108),
        Din0 => VN1018_in0,
        Din1 => VN1018_in1,
        Din2 => VN1018_in2,
        Din3 => VN1018_in3,
        Din4 => VN1018_in4,
        Din5 => VN1018_in5,
        VN2CN0_bit => VN_data_out(6108),
        VN2CN1_bit => VN_data_out(6109),
        VN2CN2_bit => VN_data_out(6110),
        VN2CN3_bit => VN_data_out(6111),
        VN2CN4_bit => VN_data_out(6112),
        VN2CN5_bit => VN_data_out(6113),
        VN2CN0_sign => VN_sign_out(6108),
        VN2CN1_sign => VN_sign_out(6109),
        VN2CN2_sign => VN_sign_out(6110),
        VN2CN3_sign => VN_sign_out(6111),
        VN2CN4_sign => VN_sign_out(6112),
        VN2CN5_sign => VN_sign_out(6113),
        codeword => codeword(1018),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1019 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6119 downto 6114),
        Din0 => VN1019_in0,
        Din1 => VN1019_in1,
        Din2 => VN1019_in2,
        Din3 => VN1019_in3,
        Din4 => VN1019_in4,
        Din5 => VN1019_in5,
        VN2CN0_bit => VN_data_out(6114),
        VN2CN1_bit => VN_data_out(6115),
        VN2CN2_bit => VN_data_out(6116),
        VN2CN3_bit => VN_data_out(6117),
        VN2CN4_bit => VN_data_out(6118),
        VN2CN5_bit => VN_data_out(6119),
        VN2CN0_sign => VN_sign_out(6114),
        VN2CN1_sign => VN_sign_out(6115),
        VN2CN2_sign => VN_sign_out(6116),
        VN2CN3_sign => VN_sign_out(6117),
        VN2CN4_sign => VN_sign_out(6118),
        VN2CN5_sign => VN_sign_out(6119),
        codeword => codeword(1019),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1020 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6125 downto 6120),
        Din0 => VN1020_in0,
        Din1 => VN1020_in1,
        Din2 => VN1020_in2,
        Din3 => VN1020_in3,
        Din4 => VN1020_in4,
        Din5 => VN1020_in5,
        VN2CN0_bit => VN_data_out(6120),
        VN2CN1_bit => VN_data_out(6121),
        VN2CN2_bit => VN_data_out(6122),
        VN2CN3_bit => VN_data_out(6123),
        VN2CN4_bit => VN_data_out(6124),
        VN2CN5_bit => VN_data_out(6125),
        VN2CN0_sign => VN_sign_out(6120),
        VN2CN1_sign => VN_sign_out(6121),
        VN2CN2_sign => VN_sign_out(6122),
        VN2CN3_sign => VN_sign_out(6123),
        VN2CN4_sign => VN_sign_out(6124),
        VN2CN5_sign => VN_sign_out(6125),
        codeword => codeword(1020),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1021 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6131 downto 6126),
        Din0 => VN1021_in0,
        Din1 => VN1021_in1,
        Din2 => VN1021_in2,
        Din3 => VN1021_in3,
        Din4 => VN1021_in4,
        Din5 => VN1021_in5,
        VN2CN0_bit => VN_data_out(6126),
        VN2CN1_bit => VN_data_out(6127),
        VN2CN2_bit => VN_data_out(6128),
        VN2CN3_bit => VN_data_out(6129),
        VN2CN4_bit => VN_data_out(6130),
        VN2CN5_bit => VN_data_out(6131),
        VN2CN0_sign => VN_sign_out(6126),
        VN2CN1_sign => VN_sign_out(6127),
        VN2CN2_sign => VN_sign_out(6128),
        VN2CN3_sign => VN_sign_out(6129),
        VN2CN4_sign => VN_sign_out(6130),
        VN2CN5_sign => VN_sign_out(6131),
        codeword => codeword(1021),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1022 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6137 downto 6132),
        Din0 => VN1022_in0,
        Din1 => VN1022_in1,
        Din2 => VN1022_in2,
        Din3 => VN1022_in3,
        Din4 => VN1022_in4,
        Din5 => VN1022_in5,
        VN2CN0_bit => VN_data_out(6132),
        VN2CN1_bit => VN_data_out(6133),
        VN2CN2_bit => VN_data_out(6134),
        VN2CN3_bit => VN_data_out(6135),
        VN2CN4_bit => VN_data_out(6136),
        VN2CN5_bit => VN_data_out(6137),
        VN2CN0_sign => VN_sign_out(6132),
        VN2CN1_sign => VN_sign_out(6133),
        VN2CN2_sign => VN_sign_out(6134),
        VN2CN3_sign => VN_sign_out(6135),
        VN2CN4_sign => VN_sign_out(6136),
        VN2CN5_sign => VN_sign_out(6137),
        codeword => codeword(1022),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1023 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6143 downto 6138),
        Din0 => VN1023_in0,
        Din1 => VN1023_in1,
        Din2 => VN1023_in2,
        Din3 => VN1023_in3,
        Din4 => VN1023_in4,
        Din5 => VN1023_in5,
        VN2CN0_bit => VN_data_out(6138),
        VN2CN1_bit => VN_data_out(6139),
        VN2CN2_bit => VN_data_out(6140),
        VN2CN3_bit => VN_data_out(6141),
        VN2CN4_bit => VN_data_out(6142),
        VN2CN5_bit => VN_data_out(6143),
        VN2CN0_sign => VN_sign_out(6138),
        VN2CN1_sign => VN_sign_out(6139),
        VN2CN2_sign => VN_sign_out(6140),
        VN2CN3_sign => VN_sign_out(6141),
        VN2CN4_sign => VN_sign_out(6142),
        VN2CN5_sign => VN_sign_out(6143),
        codeword => codeword(1023),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1024 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6149 downto 6144),
        Din0 => VN1024_in0,
        Din1 => VN1024_in1,
        Din2 => VN1024_in2,
        Din3 => VN1024_in3,
        Din4 => VN1024_in4,
        Din5 => VN1024_in5,
        VN2CN0_bit => VN_data_out(6144),
        VN2CN1_bit => VN_data_out(6145),
        VN2CN2_bit => VN_data_out(6146),
        VN2CN3_bit => VN_data_out(6147),
        VN2CN4_bit => VN_data_out(6148),
        VN2CN5_bit => VN_data_out(6149),
        VN2CN0_sign => VN_sign_out(6144),
        VN2CN1_sign => VN_sign_out(6145),
        VN2CN2_sign => VN_sign_out(6146),
        VN2CN3_sign => VN_sign_out(6147),
        VN2CN4_sign => VN_sign_out(6148),
        VN2CN5_sign => VN_sign_out(6149),
        codeword => codeword(1024),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1025 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6155 downto 6150),
        Din0 => VN1025_in0,
        Din1 => VN1025_in1,
        Din2 => VN1025_in2,
        Din3 => VN1025_in3,
        Din4 => VN1025_in4,
        Din5 => VN1025_in5,
        VN2CN0_bit => VN_data_out(6150),
        VN2CN1_bit => VN_data_out(6151),
        VN2CN2_bit => VN_data_out(6152),
        VN2CN3_bit => VN_data_out(6153),
        VN2CN4_bit => VN_data_out(6154),
        VN2CN5_bit => VN_data_out(6155),
        VN2CN0_sign => VN_sign_out(6150),
        VN2CN1_sign => VN_sign_out(6151),
        VN2CN2_sign => VN_sign_out(6152),
        VN2CN3_sign => VN_sign_out(6153),
        VN2CN4_sign => VN_sign_out(6154),
        VN2CN5_sign => VN_sign_out(6155),
        codeword => codeword(1025),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1026 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6161 downto 6156),
        Din0 => VN1026_in0,
        Din1 => VN1026_in1,
        Din2 => VN1026_in2,
        Din3 => VN1026_in3,
        Din4 => VN1026_in4,
        Din5 => VN1026_in5,
        VN2CN0_bit => VN_data_out(6156),
        VN2CN1_bit => VN_data_out(6157),
        VN2CN2_bit => VN_data_out(6158),
        VN2CN3_bit => VN_data_out(6159),
        VN2CN4_bit => VN_data_out(6160),
        VN2CN5_bit => VN_data_out(6161),
        VN2CN0_sign => VN_sign_out(6156),
        VN2CN1_sign => VN_sign_out(6157),
        VN2CN2_sign => VN_sign_out(6158),
        VN2CN3_sign => VN_sign_out(6159),
        VN2CN4_sign => VN_sign_out(6160),
        VN2CN5_sign => VN_sign_out(6161),
        codeword => codeword(1026),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1027 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6167 downto 6162),
        Din0 => VN1027_in0,
        Din1 => VN1027_in1,
        Din2 => VN1027_in2,
        Din3 => VN1027_in3,
        Din4 => VN1027_in4,
        Din5 => VN1027_in5,
        VN2CN0_bit => VN_data_out(6162),
        VN2CN1_bit => VN_data_out(6163),
        VN2CN2_bit => VN_data_out(6164),
        VN2CN3_bit => VN_data_out(6165),
        VN2CN4_bit => VN_data_out(6166),
        VN2CN5_bit => VN_data_out(6167),
        VN2CN0_sign => VN_sign_out(6162),
        VN2CN1_sign => VN_sign_out(6163),
        VN2CN2_sign => VN_sign_out(6164),
        VN2CN3_sign => VN_sign_out(6165),
        VN2CN4_sign => VN_sign_out(6166),
        VN2CN5_sign => VN_sign_out(6167),
        codeword => codeword(1027),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1028 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6173 downto 6168),
        Din0 => VN1028_in0,
        Din1 => VN1028_in1,
        Din2 => VN1028_in2,
        Din3 => VN1028_in3,
        Din4 => VN1028_in4,
        Din5 => VN1028_in5,
        VN2CN0_bit => VN_data_out(6168),
        VN2CN1_bit => VN_data_out(6169),
        VN2CN2_bit => VN_data_out(6170),
        VN2CN3_bit => VN_data_out(6171),
        VN2CN4_bit => VN_data_out(6172),
        VN2CN5_bit => VN_data_out(6173),
        VN2CN0_sign => VN_sign_out(6168),
        VN2CN1_sign => VN_sign_out(6169),
        VN2CN2_sign => VN_sign_out(6170),
        VN2CN3_sign => VN_sign_out(6171),
        VN2CN4_sign => VN_sign_out(6172),
        VN2CN5_sign => VN_sign_out(6173),
        codeword => codeword(1028),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1029 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6179 downto 6174),
        Din0 => VN1029_in0,
        Din1 => VN1029_in1,
        Din2 => VN1029_in2,
        Din3 => VN1029_in3,
        Din4 => VN1029_in4,
        Din5 => VN1029_in5,
        VN2CN0_bit => VN_data_out(6174),
        VN2CN1_bit => VN_data_out(6175),
        VN2CN2_bit => VN_data_out(6176),
        VN2CN3_bit => VN_data_out(6177),
        VN2CN4_bit => VN_data_out(6178),
        VN2CN5_bit => VN_data_out(6179),
        VN2CN0_sign => VN_sign_out(6174),
        VN2CN1_sign => VN_sign_out(6175),
        VN2CN2_sign => VN_sign_out(6176),
        VN2CN3_sign => VN_sign_out(6177),
        VN2CN4_sign => VN_sign_out(6178),
        VN2CN5_sign => VN_sign_out(6179),
        codeword => codeword(1029),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1030 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6185 downto 6180),
        Din0 => VN1030_in0,
        Din1 => VN1030_in1,
        Din2 => VN1030_in2,
        Din3 => VN1030_in3,
        Din4 => VN1030_in4,
        Din5 => VN1030_in5,
        VN2CN0_bit => VN_data_out(6180),
        VN2CN1_bit => VN_data_out(6181),
        VN2CN2_bit => VN_data_out(6182),
        VN2CN3_bit => VN_data_out(6183),
        VN2CN4_bit => VN_data_out(6184),
        VN2CN5_bit => VN_data_out(6185),
        VN2CN0_sign => VN_sign_out(6180),
        VN2CN1_sign => VN_sign_out(6181),
        VN2CN2_sign => VN_sign_out(6182),
        VN2CN3_sign => VN_sign_out(6183),
        VN2CN4_sign => VN_sign_out(6184),
        VN2CN5_sign => VN_sign_out(6185),
        codeword => codeword(1030),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1031 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6191 downto 6186),
        Din0 => VN1031_in0,
        Din1 => VN1031_in1,
        Din2 => VN1031_in2,
        Din3 => VN1031_in3,
        Din4 => VN1031_in4,
        Din5 => VN1031_in5,
        VN2CN0_bit => VN_data_out(6186),
        VN2CN1_bit => VN_data_out(6187),
        VN2CN2_bit => VN_data_out(6188),
        VN2CN3_bit => VN_data_out(6189),
        VN2CN4_bit => VN_data_out(6190),
        VN2CN5_bit => VN_data_out(6191),
        VN2CN0_sign => VN_sign_out(6186),
        VN2CN1_sign => VN_sign_out(6187),
        VN2CN2_sign => VN_sign_out(6188),
        VN2CN3_sign => VN_sign_out(6189),
        VN2CN4_sign => VN_sign_out(6190),
        VN2CN5_sign => VN_sign_out(6191),
        codeword => codeword(1031),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1032 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6197 downto 6192),
        Din0 => VN1032_in0,
        Din1 => VN1032_in1,
        Din2 => VN1032_in2,
        Din3 => VN1032_in3,
        Din4 => VN1032_in4,
        Din5 => VN1032_in5,
        VN2CN0_bit => VN_data_out(6192),
        VN2CN1_bit => VN_data_out(6193),
        VN2CN2_bit => VN_data_out(6194),
        VN2CN3_bit => VN_data_out(6195),
        VN2CN4_bit => VN_data_out(6196),
        VN2CN5_bit => VN_data_out(6197),
        VN2CN0_sign => VN_sign_out(6192),
        VN2CN1_sign => VN_sign_out(6193),
        VN2CN2_sign => VN_sign_out(6194),
        VN2CN3_sign => VN_sign_out(6195),
        VN2CN4_sign => VN_sign_out(6196),
        VN2CN5_sign => VN_sign_out(6197),
        codeword => codeword(1032),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1033 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6203 downto 6198),
        Din0 => VN1033_in0,
        Din1 => VN1033_in1,
        Din2 => VN1033_in2,
        Din3 => VN1033_in3,
        Din4 => VN1033_in4,
        Din5 => VN1033_in5,
        VN2CN0_bit => VN_data_out(6198),
        VN2CN1_bit => VN_data_out(6199),
        VN2CN2_bit => VN_data_out(6200),
        VN2CN3_bit => VN_data_out(6201),
        VN2CN4_bit => VN_data_out(6202),
        VN2CN5_bit => VN_data_out(6203),
        VN2CN0_sign => VN_sign_out(6198),
        VN2CN1_sign => VN_sign_out(6199),
        VN2CN2_sign => VN_sign_out(6200),
        VN2CN3_sign => VN_sign_out(6201),
        VN2CN4_sign => VN_sign_out(6202),
        VN2CN5_sign => VN_sign_out(6203),
        codeword => codeword(1033),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1034 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6209 downto 6204),
        Din0 => VN1034_in0,
        Din1 => VN1034_in1,
        Din2 => VN1034_in2,
        Din3 => VN1034_in3,
        Din4 => VN1034_in4,
        Din5 => VN1034_in5,
        VN2CN0_bit => VN_data_out(6204),
        VN2CN1_bit => VN_data_out(6205),
        VN2CN2_bit => VN_data_out(6206),
        VN2CN3_bit => VN_data_out(6207),
        VN2CN4_bit => VN_data_out(6208),
        VN2CN5_bit => VN_data_out(6209),
        VN2CN0_sign => VN_sign_out(6204),
        VN2CN1_sign => VN_sign_out(6205),
        VN2CN2_sign => VN_sign_out(6206),
        VN2CN3_sign => VN_sign_out(6207),
        VN2CN4_sign => VN_sign_out(6208),
        VN2CN5_sign => VN_sign_out(6209),
        codeword => codeword(1034),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1035 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6215 downto 6210),
        Din0 => VN1035_in0,
        Din1 => VN1035_in1,
        Din2 => VN1035_in2,
        Din3 => VN1035_in3,
        Din4 => VN1035_in4,
        Din5 => VN1035_in5,
        VN2CN0_bit => VN_data_out(6210),
        VN2CN1_bit => VN_data_out(6211),
        VN2CN2_bit => VN_data_out(6212),
        VN2CN3_bit => VN_data_out(6213),
        VN2CN4_bit => VN_data_out(6214),
        VN2CN5_bit => VN_data_out(6215),
        VN2CN0_sign => VN_sign_out(6210),
        VN2CN1_sign => VN_sign_out(6211),
        VN2CN2_sign => VN_sign_out(6212),
        VN2CN3_sign => VN_sign_out(6213),
        VN2CN4_sign => VN_sign_out(6214),
        VN2CN5_sign => VN_sign_out(6215),
        codeword => codeword(1035),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1036 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6221 downto 6216),
        Din0 => VN1036_in0,
        Din1 => VN1036_in1,
        Din2 => VN1036_in2,
        Din3 => VN1036_in3,
        Din4 => VN1036_in4,
        Din5 => VN1036_in5,
        VN2CN0_bit => VN_data_out(6216),
        VN2CN1_bit => VN_data_out(6217),
        VN2CN2_bit => VN_data_out(6218),
        VN2CN3_bit => VN_data_out(6219),
        VN2CN4_bit => VN_data_out(6220),
        VN2CN5_bit => VN_data_out(6221),
        VN2CN0_sign => VN_sign_out(6216),
        VN2CN1_sign => VN_sign_out(6217),
        VN2CN2_sign => VN_sign_out(6218),
        VN2CN3_sign => VN_sign_out(6219),
        VN2CN4_sign => VN_sign_out(6220),
        VN2CN5_sign => VN_sign_out(6221),
        codeword => codeword(1036),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1037 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6227 downto 6222),
        Din0 => VN1037_in0,
        Din1 => VN1037_in1,
        Din2 => VN1037_in2,
        Din3 => VN1037_in3,
        Din4 => VN1037_in4,
        Din5 => VN1037_in5,
        VN2CN0_bit => VN_data_out(6222),
        VN2CN1_bit => VN_data_out(6223),
        VN2CN2_bit => VN_data_out(6224),
        VN2CN3_bit => VN_data_out(6225),
        VN2CN4_bit => VN_data_out(6226),
        VN2CN5_bit => VN_data_out(6227),
        VN2CN0_sign => VN_sign_out(6222),
        VN2CN1_sign => VN_sign_out(6223),
        VN2CN2_sign => VN_sign_out(6224),
        VN2CN3_sign => VN_sign_out(6225),
        VN2CN4_sign => VN_sign_out(6226),
        VN2CN5_sign => VN_sign_out(6227),
        codeword => codeword(1037),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1038 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6233 downto 6228),
        Din0 => VN1038_in0,
        Din1 => VN1038_in1,
        Din2 => VN1038_in2,
        Din3 => VN1038_in3,
        Din4 => VN1038_in4,
        Din5 => VN1038_in5,
        VN2CN0_bit => VN_data_out(6228),
        VN2CN1_bit => VN_data_out(6229),
        VN2CN2_bit => VN_data_out(6230),
        VN2CN3_bit => VN_data_out(6231),
        VN2CN4_bit => VN_data_out(6232),
        VN2CN5_bit => VN_data_out(6233),
        VN2CN0_sign => VN_sign_out(6228),
        VN2CN1_sign => VN_sign_out(6229),
        VN2CN2_sign => VN_sign_out(6230),
        VN2CN3_sign => VN_sign_out(6231),
        VN2CN4_sign => VN_sign_out(6232),
        VN2CN5_sign => VN_sign_out(6233),
        codeword => codeword(1038),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1039 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6239 downto 6234),
        Din0 => VN1039_in0,
        Din1 => VN1039_in1,
        Din2 => VN1039_in2,
        Din3 => VN1039_in3,
        Din4 => VN1039_in4,
        Din5 => VN1039_in5,
        VN2CN0_bit => VN_data_out(6234),
        VN2CN1_bit => VN_data_out(6235),
        VN2CN2_bit => VN_data_out(6236),
        VN2CN3_bit => VN_data_out(6237),
        VN2CN4_bit => VN_data_out(6238),
        VN2CN5_bit => VN_data_out(6239),
        VN2CN0_sign => VN_sign_out(6234),
        VN2CN1_sign => VN_sign_out(6235),
        VN2CN2_sign => VN_sign_out(6236),
        VN2CN3_sign => VN_sign_out(6237),
        VN2CN4_sign => VN_sign_out(6238),
        VN2CN5_sign => VN_sign_out(6239),
        codeword => codeword(1039),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1040 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6245 downto 6240),
        Din0 => VN1040_in0,
        Din1 => VN1040_in1,
        Din2 => VN1040_in2,
        Din3 => VN1040_in3,
        Din4 => VN1040_in4,
        Din5 => VN1040_in5,
        VN2CN0_bit => VN_data_out(6240),
        VN2CN1_bit => VN_data_out(6241),
        VN2CN2_bit => VN_data_out(6242),
        VN2CN3_bit => VN_data_out(6243),
        VN2CN4_bit => VN_data_out(6244),
        VN2CN5_bit => VN_data_out(6245),
        VN2CN0_sign => VN_sign_out(6240),
        VN2CN1_sign => VN_sign_out(6241),
        VN2CN2_sign => VN_sign_out(6242),
        VN2CN3_sign => VN_sign_out(6243),
        VN2CN4_sign => VN_sign_out(6244),
        VN2CN5_sign => VN_sign_out(6245),
        codeword => codeword(1040),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1041 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6251 downto 6246),
        Din0 => VN1041_in0,
        Din1 => VN1041_in1,
        Din2 => VN1041_in2,
        Din3 => VN1041_in3,
        Din4 => VN1041_in4,
        Din5 => VN1041_in5,
        VN2CN0_bit => VN_data_out(6246),
        VN2CN1_bit => VN_data_out(6247),
        VN2CN2_bit => VN_data_out(6248),
        VN2CN3_bit => VN_data_out(6249),
        VN2CN4_bit => VN_data_out(6250),
        VN2CN5_bit => VN_data_out(6251),
        VN2CN0_sign => VN_sign_out(6246),
        VN2CN1_sign => VN_sign_out(6247),
        VN2CN2_sign => VN_sign_out(6248),
        VN2CN3_sign => VN_sign_out(6249),
        VN2CN4_sign => VN_sign_out(6250),
        VN2CN5_sign => VN_sign_out(6251),
        codeword => codeword(1041),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1042 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6257 downto 6252),
        Din0 => VN1042_in0,
        Din1 => VN1042_in1,
        Din2 => VN1042_in2,
        Din3 => VN1042_in3,
        Din4 => VN1042_in4,
        Din5 => VN1042_in5,
        VN2CN0_bit => VN_data_out(6252),
        VN2CN1_bit => VN_data_out(6253),
        VN2CN2_bit => VN_data_out(6254),
        VN2CN3_bit => VN_data_out(6255),
        VN2CN4_bit => VN_data_out(6256),
        VN2CN5_bit => VN_data_out(6257),
        VN2CN0_sign => VN_sign_out(6252),
        VN2CN1_sign => VN_sign_out(6253),
        VN2CN2_sign => VN_sign_out(6254),
        VN2CN3_sign => VN_sign_out(6255),
        VN2CN4_sign => VN_sign_out(6256),
        VN2CN5_sign => VN_sign_out(6257),
        codeword => codeword(1042),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1043 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6263 downto 6258),
        Din0 => VN1043_in0,
        Din1 => VN1043_in1,
        Din2 => VN1043_in2,
        Din3 => VN1043_in3,
        Din4 => VN1043_in4,
        Din5 => VN1043_in5,
        VN2CN0_bit => VN_data_out(6258),
        VN2CN1_bit => VN_data_out(6259),
        VN2CN2_bit => VN_data_out(6260),
        VN2CN3_bit => VN_data_out(6261),
        VN2CN4_bit => VN_data_out(6262),
        VN2CN5_bit => VN_data_out(6263),
        VN2CN0_sign => VN_sign_out(6258),
        VN2CN1_sign => VN_sign_out(6259),
        VN2CN2_sign => VN_sign_out(6260),
        VN2CN3_sign => VN_sign_out(6261),
        VN2CN4_sign => VN_sign_out(6262),
        VN2CN5_sign => VN_sign_out(6263),
        codeword => codeword(1043),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1044 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6269 downto 6264),
        Din0 => VN1044_in0,
        Din1 => VN1044_in1,
        Din2 => VN1044_in2,
        Din3 => VN1044_in3,
        Din4 => VN1044_in4,
        Din5 => VN1044_in5,
        VN2CN0_bit => VN_data_out(6264),
        VN2CN1_bit => VN_data_out(6265),
        VN2CN2_bit => VN_data_out(6266),
        VN2CN3_bit => VN_data_out(6267),
        VN2CN4_bit => VN_data_out(6268),
        VN2CN5_bit => VN_data_out(6269),
        VN2CN0_sign => VN_sign_out(6264),
        VN2CN1_sign => VN_sign_out(6265),
        VN2CN2_sign => VN_sign_out(6266),
        VN2CN3_sign => VN_sign_out(6267),
        VN2CN4_sign => VN_sign_out(6268),
        VN2CN5_sign => VN_sign_out(6269),
        codeword => codeword(1044),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1045 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6275 downto 6270),
        Din0 => VN1045_in0,
        Din1 => VN1045_in1,
        Din2 => VN1045_in2,
        Din3 => VN1045_in3,
        Din4 => VN1045_in4,
        Din5 => VN1045_in5,
        VN2CN0_bit => VN_data_out(6270),
        VN2CN1_bit => VN_data_out(6271),
        VN2CN2_bit => VN_data_out(6272),
        VN2CN3_bit => VN_data_out(6273),
        VN2CN4_bit => VN_data_out(6274),
        VN2CN5_bit => VN_data_out(6275),
        VN2CN0_sign => VN_sign_out(6270),
        VN2CN1_sign => VN_sign_out(6271),
        VN2CN2_sign => VN_sign_out(6272),
        VN2CN3_sign => VN_sign_out(6273),
        VN2CN4_sign => VN_sign_out(6274),
        VN2CN5_sign => VN_sign_out(6275),
        codeword => codeword(1045),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1046 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6281 downto 6276),
        Din0 => VN1046_in0,
        Din1 => VN1046_in1,
        Din2 => VN1046_in2,
        Din3 => VN1046_in3,
        Din4 => VN1046_in4,
        Din5 => VN1046_in5,
        VN2CN0_bit => VN_data_out(6276),
        VN2CN1_bit => VN_data_out(6277),
        VN2CN2_bit => VN_data_out(6278),
        VN2CN3_bit => VN_data_out(6279),
        VN2CN4_bit => VN_data_out(6280),
        VN2CN5_bit => VN_data_out(6281),
        VN2CN0_sign => VN_sign_out(6276),
        VN2CN1_sign => VN_sign_out(6277),
        VN2CN2_sign => VN_sign_out(6278),
        VN2CN3_sign => VN_sign_out(6279),
        VN2CN4_sign => VN_sign_out(6280),
        VN2CN5_sign => VN_sign_out(6281),
        codeword => codeword(1046),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1047 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6287 downto 6282),
        Din0 => VN1047_in0,
        Din1 => VN1047_in1,
        Din2 => VN1047_in2,
        Din3 => VN1047_in3,
        Din4 => VN1047_in4,
        Din5 => VN1047_in5,
        VN2CN0_bit => VN_data_out(6282),
        VN2CN1_bit => VN_data_out(6283),
        VN2CN2_bit => VN_data_out(6284),
        VN2CN3_bit => VN_data_out(6285),
        VN2CN4_bit => VN_data_out(6286),
        VN2CN5_bit => VN_data_out(6287),
        VN2CN0_sign => VN_sign_out(6282),
        VN2CN1_sign => VN_sign_out(6283),
        VN2CN2_sign => VN_sign_out(6284),
        VN2CN3_sign => VN_sign_out(6285),
        VN2CN4_sign => VN_sign_out(6286),
        VN2CN5_sign => VN_sign_out(6287),
        codeword => codeword(1047),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1048 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6293 downto 6288),
        Din0 => VN1048_in0,
        Din1 => VN1048_in1,
        Din2 => VN1048_in2,
        Din3 => VN1048_in3,
        Din4 => VN1048_in4,
        Din5 => VN1048_in5,
        VN2CN0_bit => VN_data_out(6288),
        VN2CN1_bit => VN_data_out(6289),
        VN2CN2_bit => VN_data_out(6290),
        VN2CN3_bit => VN_data_out(6291),
        VN2CN4_bit => VN_data_out(6292),
        VN2CN5_bit => VN_data_out(6293),
        VN2CN0_sign => VN_sign_out(6288),
        VN2CN1_sign => VN_sign_out(6289),
        VN2CN2_sign => VN_sign_out(6290),
        VN2CN3_sign => VN_sign_out(6291),
        VN2CN4_sign => VN_sign_out(6292),
        VN2CN5_sign => VN_sign_out(6293),
        codeword => codeword(1048),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1049 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6299 downto 6294),
        Din0 => VN1049_in0,
        Din1 => VN1049_in1,
        Din2 => VN1049_in2,
        Din3 => VN1049_in3,
        Din4 => VN1049_in4,
        Din5 => VN1049_in5,
        VN2CN0_bit => VN_data_out(6294),
        VN2CN1_bit => VN_data_out(6295),
        VN2CN2_bit => VN_data_out(6296),
        VN2CN3_bit => VN_data_out(6297),
        VN2CN4_bit => VN_data_out(6298),
        VN2CN5_bit => VN_data_out(6299),
        VN2CN0_sign => VN_sign_out(6294),
        VN2CN1_sign => VN_sign_out(6295),
        VN2CN2_sign => VN_sign_out(6296),
        VN2CN3_sign => VN_sign_out(6297),
        VN2CN4_sign => VN_sign_out(6298),
        VN2CN5_sign => VN_sign_out(6299),
        codeword => codeword(1049),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1050 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6305 downto 6300),
        Din0 => VN1050_in0,
        Din1 => VN1050_in1,
        Din2 => VN1050_in2,
        Din3 => VN1050_in3,
        Din4 => VN1050_in4,
        Din5 => VN1050_in5,
        VN2CN0_bit => VN_data_out(6300),
        VN2CN1_bit => VN_data_out(6301),
        VN2CN2_bit => VN_data_out(6302),
        VN2CN3_bit => VN_data_out(6303),
        VN2CN4_bit => VN_data_out(6304),
        VN2CN5_bit => VN_data_out(6305),
        VN2CN0_sign => VN_sign_out(6300),
        VN2CN1_sign => VN_sign_out(6301),
        VN2CN2_sign => VN_sign_out(6302),
        VN2CN3_sign => VN_sign_out(6303),
        VN2CN4_sign => VN_sign_out(6304),
        VN2CN5_sign => VN_sign_out(6305),
        codeword => codeword(1050),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1051 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6311 downto 6306),
        Din0 => VN1051_in0,
        Din1 => VN1051_in1,
        Din2 => VN1051_in2,
        Din3 => VN1051_in3,
        Din4 => VN1051_in4,
        Din5 => VN1051_in5,
        VN2CN0_bit => VN_data_out(6306),
        VN2CN1_bit => VN_data_out(6307),
        VN2CN2_bit => VN_data_out(6308),
        VN2CN3_bit => VN_data_out(6309),
        VN2CN4_bit => VN_data_out(6310),
        VN2CN5_bit => VN_data_out(6311),
        VN2CN0_sign => VN_sign_out(6306),
        VN2CN1_sign => VN_sign_out(6307),
        VN2CN2_sign => VN_sign_out(6308),
        VN2CN3_sign => VN_sign_out(6309),
        VN2CN4_sign => VN_sign_out(6310),
        VN2CN5_sign => VN_sign_out(6311),
        codeword => codeword(1051),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1052 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6317 downto 6312),
        Din0 => VN1052_in0,
        Din1 => VN1052_in1,
        Din2 => VN1052_in2,
        Din3 => VN1052_in3,
        Din4 => VN1052_in4,
        Din5 => VN1052_in5,
        VN2CN0_bit => VN_data_out(6312),
        VN2CN1_bit => VN_data_out(6313),
        VN2CN2_bit => VN_data_out(6314),
        VN2CN3_bit => VN_data_out(6315),
        VN2CN4_bit => VN_data_out(6316),
        VN2CN5_bit => VN_data_out(6317),
        VN2CN0_sign => VN_sign_out(6312),
        VN2CN1_sign => VN_sign_out(6313),
        VN2CN2_sign => VN_sign_out(6314),
        VN2CN3_sign => VN_sign_out(6315),
        VN2CN4_sign => VN_sign_out(6316),
        VN2CN5_sign => VN_sign_out(6317),
        codeword => codeword(1052),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1053 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6323 downto 6318),
        Din0 => VN1053_in0,
        Din1 => VN1053_in1,
        Din2 => VN1053_in2,
        Din3 => VN1053_in3,
        Din4 => VN1053_in4,
        Din5 => VN1053_in5,
        VN2CN0_bit => VN_data_out(6318),
        VN2CN1_bit => VN_data_out(6319),
        VN2CN2_bit => VN_data_out(6320),
        VN2CN3_bit => VN_data_out(6321),
        VN2CN4_bit => VN_data_out(6322),
        VN2CN5_bit => VN_data_out(6323),
        VN2CN0_sign => VN_sign_out(6318),
        VN2CN1_sign => VN_sign_out(6319),
        VN2CN2_sign => VN_sign_out(6320),
        VN2CN3_sign => VN_sign_out(6321),
        VN2CN4_sign => VN_sign_out(6322),
        VN2CN5_sign => VN_sign_out(6323),
        codeword => codeword(1053),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1054 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6329 downto 6324),
        Din0 => VN1054_in0,
        Din1 => VN1054_in1,
        Din2 => VN1054_in2,
        Din3 => VN1054_in3,
        Din4 => VN1054_in4,
        Din5 => VN1054_in5,
        VN2CN0_bit => VN_data_out(6324),
        VN2CN1_bit => VN_data_out(6325),
        VN2CN2_bit => VN_data_out(6326),
        VN2CN3_bit => VN_data_out(6327),
        VN2CN4_bit => VN_data_out(6328),
        VN2CN5_bit => VN_data_out(6329),
        VN2CN0_sign => VN_sign_out(6324),
        VN2CN1_sign => VN_sign_out(6325),
        VN2CN2_sign => VN_sign_out(6326),
        VN2CN3_sign => VN_sign_out(6327),
        VN2CN4_sign => VN_sign_out(6328),
        VN2CN5_sign => VN_sign_out(6329),
        codeword => codeword(1054),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1055 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6335 downto 6330),
        Din0 => VN1055_in0,
        Din1 => VN1055_in1,
        Din2 => VN1055_in2,
        Din3 => VN1055_in3,
        Din4 => VN1055_in4,
        Din5 => VN1055_in5,
        VN2CN0_bit => VN_data_out(6330),
        VN2CN1_bit => VN_data_out(6331),
        VN2CN2_bit => VN_data_out(6332),
        VN2CN3_bit => VN_data_out(6333),
        VN2CN4_bit => VN_data_out(6334),
        VN2CN5_bit => VN_data_out(6335),
        VN2CN0_sign => VN_sign_out(6330),
        VN2CN1_sign => VN_sign_out(6331),
        VN2CN2_sign => VN_sign_out(6332),
        VN2CN3_sign => VN_sign_out(6333),
        VN2CN4_sign => VN_sign_out(6334),
        VN2CN5_sign => VN_sign_out(6335),
        codeword => codeword(1055),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1056 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6341 downto 6336),
        Din0 => VN1056_in0,
        Din1 => VN1056_in1,
        Din2 => VN1056_in2,
        Din3 => VN1056_in3,
        Din4 => VN1056_in4,
        Din5 => VN1056_in5,
        VN2CN0_bit => VN_data_out(6336),
        VN2CN1_bit => VN_data_out(6337),
        VN2CN2_bit => VN_data_out(6338),
        VN2CN3_bit => VN_data_out(6339),
        VN2CN4_bit => VN_data_out(6340),
        VN2CN5_bit => VN_data_out(6341),
        VN2CN0_sign => VN_sign_out(6336),
        VN2CN1_sign => VN_sign_out(6337),
        VN2CN2_sign => VN_sign_out(6338),
        VN2CN3_sign => VN_sign_out(6339),
        VN2CN4_sign => VN_sign_out(6340),
        VN2CN5_sign => VN_sign_out(6341),
        codeword => codeword(1056),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1057 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6347 downto 6342),
        Din0 => VN1057_in0,
        Din1 => VN1057_in1,
        Din2 => VN1057_in2,
        Din3 => VN1057_in3,
        Din4 => VN1057_in4,
        Din5 => VN1057_in5,
        VN2CN0_bit => VN_data_out(6342),
        VN2CN1_bit => VN_data_out(6343),
        VN2CN2_bit => VN_data_out(6344),
        VN2CN3_bit => VN_data_out(6345),
        VN2CN4_bit => VN_data_out(6346),
        VN2CN5_bit => VN_data_out(6347),
        VN2CN0_sign => VN_sign_out(6342),
        VN2CN1_sign => VN_sign_out(6343),
        VN2CN2_sign => VN_sign_out(6344),
        VN2CN3_sign => VN_sign_out(6345),
        VN2CN4_sign => VN_sign_out(6346),
        VN2CN5_sign => VN_sign_out(6347),
        codeword => codeword(1057),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1058 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6353 downto 6348),
        Din0 => VN1058_in0,
        Din1 => VN1058_in1,
        Din2 => VN1058_in2,
        Din3 => VN1058_in3,
        Din4 => VN1058_in4,
        Din5 => VN1058_in5,
        VN2CN0_bit => VN_data_out(6348),
        VN2CN1_bit => VN_data_out(6349),
        VN2CN2_bit => VN_data_out(6350),
        VN2CN3_bit => VN_data_out(6351),
        VN2CN4_bit => VN_data_out(6352),
        VN2CN5_bit => VN_data_out(6353),
        VN2CN0_sign => VN_sign_out(6348),
        VN2CN1_sign => VN_sign_out(6349),
        VN2CN2_sign => VN_sign_out(6350),
        VN2CN3_sign => VN_sign_out(6351),
        VN2CN4_sign => VN_sign_out(6352),
        VN2CN5_sign => VN_sign_out(6353),
        codeword => codeword(1058),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1059 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6359 downto 6354),
        Din0 => VN1059_in0,
        Din1 => VN1059_in1,
        Din2 => VN1059_in2,
        Din3 => VN1059_in3,
        Din4 => VN1059_in4,
        Din5 => VN1059_in5,
        VN2CN0_bit => VN_data_out(6354),
        VN2CN1_bit => VN_data_out(6355),
        VN2CN2_bit => VN_data_out(6356),
        VN2CN3_bit => VN_data_out(6357),
        VN2CN4_bit => VN_data_out(6358),
        VN2CN5_bit => VN_data_out(6359),
        VN2CN0_sign => VN_sign_out(6354),
        VN2CN1_sign => VN_sign_out(6355),
        VN2CN2_sign => VN_sign_out(6356),
        VN2CN3_sign => VN_sign_out(6357),
        VN2CN4_sign => VN_sign_out(6358),
        VN2CN5_sign => VN_sign_out(6359),
        codeword => codeword(1059),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1060 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6365 downto 6360),
        Din0 => VN1060_in0,
        Din1 => VN1060_in1,
        Din2 => VN1060_in2,
        Din3 => VN1060_in3,
        Din4 => VN1060_in4,
        Din5 => VN1060_in5,
        VN2CN0_bit => VN_data_out(6360),
        VN2CN1_bit => VN_data_out(6361),
        VN2CN2_bit => VN_data_out(6362),
        VN2CN3_bit => VN_data_out(6363),
        VN2CN4_bit => VN_data_out(6364),
        VN2CN5_bit => VN_data_out(6365),
        VN2CN0_sign => VN_sign_out(6360),
        VN2CN1_sign => VN_sign_out(6361),
        VN2CN2_sign => VN_sign_out(6362),
        VN2CN3_sign => VN_sign_out(6363),
        VN2CN4_sign => VN_sign_out(6364),
        VN2CN5_sign => VN_sign_out(6365),
        codeword => codeword(1060),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1061 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6371 downto 6366),
        Din0 => VN1061_in0,
        Din1 => VN1061_in1,
        Din2 => VN1061_in2,
        Din3 => VN1061_in3,
        Din4 => VN1061_in4,
        Din5 => VN1061_in5,
        VN2CN0_bit => VN_data_out(6366),
        VN2CN1_bit => VN_data_out(6367),
        VN2CN2_bit => VN_data_out(6368),
        VN2CN3_bit => VN_data_out(6369),
        VN2CN4_bit => VN_data_out(6370),
        VN2CN5_bit => VN_data_out(6371),
        VN2CN0_sign => VN_sign_out(6366),
        VN2CN1_sign => VN_sign_out(6367),
        VN2CN2_sign => VN_sign_out(6368),
        VN2CN3_sign => VN_sign_out(6369),
        VN2CN4_sign => VN_sign_out(6370),
        VN2CN5_sign => VN_sign_out(6371),
        codeword => codeword(1061),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1062 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6377 downto 6372),
        Din0 => VN1062_in0,
        Din1 => VN1062_in1,
        Din2 => VN1062_in2,
        Din3 => VN1062_in3,
        Din4 => VN1062_in4,
        Din5 => VN1062_in5,
        VN2CN0_bit => VN_data_out(6372),
        VN2CN1_bit => VN_data_out(6373),
        VN2CN2_bit => VN_data_out(6374),
        VN2CN3_bit => VN_data_out(6375),
        VN2CN4_bit => VN_data_out(6376),
        VN2CN5_bit => VN_data_out(6377),
        VN2CN0_sign => VN_sign_out(6372),
        VN2CN1_sign => VN_sign_out(6373),
        VN2CN2_sign => VN_sign_out(6374),
        VN2CN3_sign => VN_sign_out(6375),
        VN2CN4_sign => VN_sign_out(6376),
        VN2CN5_sign => VN_sign_out(6377),
        codeword => codeword(1062),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1063 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6383 downto 6378),
        Din0 => VN1063_in0,
        Din1 => VN1063_in1,
        Din2 => VN1063_in2,
        Din3 => VN1063_in3,
        Din4 => VN1063_in4,
        Din5 => VN1063_in5,
        VN2CN0_bit => VN_data_out(6378),
        VN2CN1_bit => VN_data_out(6379),
        VN2CN2_bit => VN_data_out(6380),
        VN2CN3_bit => VN_data_out(6381),
        VN2CN4_bit => VN_data_out(6382),
        VN2CN5_bit => VN_data_out(6383),
        VN2CN0_sign => VN_sign_out(6378),
        VN2CN1_sign => VN_sign_out(6379),
        VN2CN2_sign => VN_sign_out(6380),
        VN2CN3_sign => VN_sign_out(6381),
        VN2CN4_sign => VN_sign_out(6382),
        VN2CN5_sign => VN_sign_out(6383),
        codeword => codeword(1063),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1064 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6389 downto 6384),
        Din0 => VN1064_in0,
        Din1 => VN1064_in1,
        Din2 => VN1064_in2,
        Din3 => VN1064_in3,
        Din4 => VN1064_in4,
        Din5 => VN1064_in5,
        VN2CN0_bit => VN_data_out(6384),
        VN2CN1_bit => VN_data_out(6385),
        VN2CN2_bit => VN_data_out(6386),
        VN2CN3_bit => VN_data_out(6387),
        VN2CN4_bit => VN_data_out(6388),
        VN2CN5_bit => VN_data_out(6389),
        VN2CN0_sign => VN_sign_out(6384),
        VN2CN1_sign => VN_sign_out(6385),
        VN2CN2_sign => VN_sign_out(6386),
        VN2CN3_sign => VN_sign_out(6387),
        VN2CN4_sign => VN_sign_out(6388),
        VN2CN5_sign => VN_sign_out(6389),
        codeword => codeword(1064),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1065 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6395 downto 6390),
        Din0 => VN1065_in0,
        Din1 => VN1065_in1,
        Din2 => VN1065_in2,
        Din3 => VN1065_in3,
        Din4 => VN1065_in4,
        Din5 => VN1065_in5,
        VN2CN0_bit => VN_data_out(6390),
        VN2CN1_bit => VN_data_out(6391),
        VN2CN2_bit => VN_data_out(6392),
        VN2CN3_bit => VN_data_out(6393),
        VN2CN4_bit => VN_data_out(6394),
        VN2CN5_bit => VN_data_out(6395),
        VN2CN0_sign => VN_sign_out(6390),
        VN2CN1_sign => VN_sign_out(6391),
        VN2CN2_sign => VN_sign_out(6392),
        VN2CN3_sign => VN_sign_out(6393),
        VN2CN4_sign => VN_sign_out(6394),
        VN2CN5_sign => VN_sign_out(6395),
        codeword => codeword(1065),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1066 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6401 downto 6396),
        Din0 => VN1066_in0,
        Din1 => VN1066_in1,
        Din2 => VN1066_in2,
        Din3 => VN1066_in3,
        Din4 => VN1066_in4,
        Din5 => VN1066_in5,
        VN2CN0_bit => VN_data_out(6396),
        VN2CN1_bit => VN_data_out(6397),
        VN2CN2_bit => VN_data_out(6398),
        VN2CN3_bit => VN_data_out(6399),
        VN2CN4_bit => VN_data_out(6400),
        VN2CN5_bit => VN_data_out(6401),
        VN2CN0_sign => VN_sign_out(6396),
        VN2CN1_sign => VN_sign_out(6397),
        VN2CN2_sign => VN_sign_out(6398),
        VN2CN3_sign => VN_sign_out(6399),
        VN2CN4_sign => VN_sign_out(6400),
        VN2CN5_sign => VN_sign_out(6401),
        codeword => codeword(1066),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1067 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6407 downto 6402),
        Din0 => VN1067_in0,
        Din1 => VN1067_in1,
        Din2 => VN1067_in2,
        Din3 => VN1067_in3,
        Din4 => VN1067_in4,
        Din5 => VN1067_in5,
        VN2CN0_bit => VN_data_out(6402),
        VN2CN1_bit => VN_data_out(6403),
        VN2CN2_bit => VN_data_out(6404),
        VN2CN3_bit => VN_data_out(6405),
        VN2CN4_bit => VN_data_out(6406),
        VN2CN5_bit => VN_data_out(6407),
        VN2CN0_sign => VN_sign_out(6402),
        VN2CN1_sign => VN_sign_out(6403),
        VN2CN2_sign => VN_sign_out(6404),
        VN2CN3_sign => VN_sign_out(6405),
        VN2CN4_sign => VN_sign_out(6406),
        VN2CN5_sign => VN_sign_out(6407),
        codeword => codeword(1067),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1068 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6413 downto 6408),
        Din0 => VN1068_in0,
        Din1 => VN1068_in1,
        Din2 => VN1068_in2,
        Din3 => VN1068_in3,
        Din4 => VN1068_in4,
        Din5 => VN1068_in5,
        VN2CN0_bit => VN_data_out(6408),
        VN2CN1_bit => VN_data_out(6409),
        VN2CN2_bit => VN_data_out(6410),
        VN2CN3_bit => VN_data_out(6411),
        VN2CN4_bit => VN_data_out(6412),
        VN2CN5_bit => VN_data_out(6413),
        VN2CN0_sign => VN_sign_out(6408),
        VN2CN1_sign => VN_sign_out(6409),
        VN2CN2_sign => VN_sign_out(6410),
        VN2CN3_sign => VN_sign_out(6411),
        VN2CN4_sign => VN_sign_out(6412),
        VN2CN5_sign => VN_sign_out(6413),
        codeword => codeword(1068),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1069 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6419 downto 6414),
        Din0 => VN1069_in0,
        Din1 => VN1069_in1,
        Din2 => VN1069_in2,
        Din3 => VN1069_in3,
        Din4 => VN1069_in4,
        Din5 => VN1069_in5,
        VN2CN0_bit => VN_data_out(6414),
        VN2CN1_bit => VN_data_out(6415),
        VN2CN2_bit => VN_data_out(6416),
        VN2CN3_bit => VN_data_out(6417),
        VN2CN4_bit => VN_data_out(6418),
        VN2CN5_bit => VN_data_out(6419),
        VN2CN0_sign => VN_sign_out(6414),
        VN2CN1_sign => VN_sign_out(6415),
        VN2CN2_sign => VN_sign_out(6416),
        VN2CN3_sign => VN_sign_out(6417),
        VN2CN4_sign => VN_sign_out(6418),
        VN2CN5_sign => VN_sign_out(6419),
        codeword => codeword(1069),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1070 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6425 downto 6420),
        Din0 => VN1070_in0,
        Din1 => VN1070_in1,
        Din2 => VN1070_in2,
        Din3 => VN1070_in3,
        Din4 => VN1070_in4,
        Din5 => VN1070_in5,
        VN2CN0_bit => VN_data_out(6420),
        VN2CN1_bit => VN_data_out(6421),
        VN2CN2_bit => VN_data_out(6422),
        VN2CN3_bit => VN_data_out(6423),
        VN2CN4_bit => VN_data_out(6424),
        VN2CN5_bit => VN_data_out(6425),
        VN2CN0_sign => VN_sign_out(6420),
        VN2CN1_sign => VN_sign_out(6421),
        VN2CN2_sign => VN_sign_out(6422),
        VN2CN3_sign => VN_sign_out(6423),
        VN2CN4_sign => VN_sign_out(6424),
        VN2CN5_sign => VN_sign_out(6425),
        codeword => codeword(1070),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1071 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6431 downto 6426),
        Din0 => VN1071_in0,
        Din1 => VN1071_in1,
        Din2 => VN1071_in2,
        Din3 => VN1071_in3,
        Din4 => VN1071_in4,
        Din5 => VN1071_in5,
        VN2CN0_bit => VN_data_out(6426),
        VN2CN1_bit => VN_data_out(6427),
        VN2CN2_bit => VN_data_out(6428),
        VN2CN3_bit => VN_data_out(6429),
        VN2CN4_bit => VN_data_out(6430),
        VN2CN5_bit => VN_data_out(6431),
        VN2CN0_sign => VN_sign_out(6426),
        VN2CN1_sign => VN_sign_out(6427),
        VN2CN2_sign => VN_sign_out(6428),
        VN2CN3_sign => VN_sign_out(6429),
        VN2CN4_sign => VN_sign_out(6430),
        VN2CN5_sign => VN_sign_out(6431),
        codeword => codeword(1071),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1072 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6437 downto 6432),
        Din0 => VN1072_in0,
        Din1 => VN1072_in1,
        Din2 => VN1072_in2,
        Din3 => VN1072_in3,
        Din4 => VN1072_in4,
        Din5 => VN1072_in5,
        VN2CN0_bit => VN_data_out(6432),
        VN2CN1_bit => VN_data_out(6433),
        VN2CN2_bit => VN_data_out(6434),
        VN2CN3_bit => VN_data_out(6435),
        VN2CN4_bit => VN_data_out(6436),
        VN2CN5_bit => VN_data_out(6437),
        VN2CN0_sign => VN_sign_out(6432),
        VN2CN1_sign => VN_sign_out(6433),
        VN2CN2_sign => VN_sign_out(6434),
        VN2CN3_sign => VN_sign_out(6435),
        VN2CN4_sign => VN_sign_out(6436),
        VN2CN5_sign => VN_sign_out(6437),
        codeword => codeword(1072),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1073 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6443 downto 6438),
        Din0 => VN1073_in0,
        Din1 => VN1073_in1,
        Din2 => VN1073_in2,
        Din3 => VN1073_in3,
        Din4 => VN1073_in4,
        Din5 => VN1073_in5,
        VN2CN0_bit => VN_data_out(6438),
        VN2CN1_bit => VN_data_out(6439),
        VN2CN2_bit => VN_data_out(6440),
        VN2CN3_bit => VN_data_out(6441),
        VN2CN4_bit => VN_data_out(6442),
        VN2CN5_bit => VN_data_out(6443),
        VN2CN0_sign => VN_sign_out(6438),
        VN2CN1_sign => VN_sign_out(6439),
        VN2CN2_sign => VN_sign_out(6440),
        VN2CN3_sign => VN_sign_out(6441),
        VN2CN4_sign => VN_sign_out(6442),
        VN2CN5_sign => VN_sign_out(6443),
        codeword => codeword(1073),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1074 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6449 downto 6444),
        Din0 => VN1074_in0,
        Din1 => VN1074_in1,
        Din2 => VN1074_in2,
        Din3 => VN1074_in3,
        Din4 => VN1074_in4,
        Din5 => VN1074_in5,
        VN2CN0_bit => VN_data_out(6444),
        VN2CN1_bit => VN_data_out(6445),
        VN2CN2_bit => VN_data_out(6446),
        VN2CN3_bit => VN_data_out(6447),
        VN2CN4_bit => VN_data_out(6448),
        VN2CN5_bit => VN_data_out(6449),
        VN2CN0_sign => VN_sign_out(6444),
        VN2CN1_sign => VN_sign_out(6445),
        VN2CN2_sign => VN_sign_out(6446),
        VN2CN3_sign => VN_sign_out(6447),
        VN2CN4_sign => VN_sign_out(6448),
        VN2CN5_sign => VN_sign_out(6449),
        codeword => codeword(1074),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1075 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6455 downto 6450),
        Din0 => VN1075_in0,
        Din1 => VN1075_in1,
        Din2 => VN1075_in2,
        Din3 => VN1075_in3,
        Din4 => VN1075_in4,
        Din5 => VN1075_in5,
        VN2CN0_bit => VN_data_out(6450),
        VN2CN1_bit => VN_data_out(6451),
        VN2CN2_bit => VN_data_out(6452),
        VN2CN3_bit => VN_data_out(6453),
        VN2CN4_bit => VN_data_out(6454),
        VN2CN5_bit => VN_data_out(6455),
        VN2CN0_sign => VN_sign_out(6450),
        VN2CN1_sign => VN_sign_out(6451),
        VN2CN2_sign => VN_sign_out(6452),
        VN2CN3_sign => VN_sign_out(6453),
        VN2CN4_sign => VN_sign_out(6454),
        VN2CN5_sign => VN_sign_out(6455),
        codeword => codeword(1075),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1076 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6461 downto 6456),
        Din0 => VN1076_in0,
        Din1 => VN1076_in1,
        Din2 => VN1076_in2,
        Din3 => VN1076_in3,
        Din4 => VN1076_in4,
        Din5 => VN1076_in5,
        VN2CN0_bit => VN_data_out(6456),
        VN2CN1_bit => VN_data_out(6457),
        VN2CN2_bit => VN_data_out(6458),
        VN2CN3_bit => VN_data_out(6459),
        VN2CN4_bit => VN_data_out(6460),
        VN2CN5_bit => VN_data_out(6461),
        VN2CN0_sign => VN_sign_out(6456),
        VN2CN1_sign => VN_sign_out(6457),
        VN2CN2_sign => VN_sign_out(6458),
        VN2CN3_sign => VN_sign_out(6459),
        VN2CN4_sign => VN_sign_out(6460),
        VN2CN5_sign => VN_sign_out(6461),
        codeword => codeword(1076),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1077 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6467 downto 6462),
        Din0 => VN1077_in0,
        Din1 => VN1077_in1,
        Din2 => VN1077_in2,
        Din3 => VN1077_in3,
        Din4 => VN1077_in4,
        Din5 => VN1077_in5,
        VN2CN0_bit => VN_data_out(6462),
        VN2CN1_bit => VN_data_out(6463),
        VN2CN2_bit => VN_data_out(6464),
        VN2CN3_bit => VN_data_out(6465),
        VN2CN4_bit => VN_data_out(6466),
        VN2CN5_bit => VN_data_out(6467),
        VN2CN0_sign => VN_sign_out(6462),
        VN2CN1_sign => VN_sign_out(6463),
        VN2CN2_sign => VN_sign_out(6464),
        VN2CN3_sign => VN_sign_out(6465),
        VN2CN4_sign => VN_sign_out(6466),
        VN2CN5_sign => VN_sign_out(6467),
        codeword => codeword(1077),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1078 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6473 downto 6468),
        Din0 => VN1078_in0,
        Din1 => VN1078_in1,
        Din2 => VN1078_in2,
        Din3 => VN1078_in3,
        Din4 => VN1078_in4,
        Din5 => VN1078_in5,
        VN2CN0_bit => VN_data_out(6468),
        VN2CN1_bit => VN_data_out(6469),
        VN2CN2_bit => VN_data_out(6470),
        VN2CN3_bit => VN_data_out(6471),
        VN2CN4_bit => VN_data_out(6472),
        VN2CN5_bit => VN_data_out(6473),
        VN2CN0_sign => VN_sign_out(6468),
        VN2CN1_sign => VN_sign_out(6469),
        VN2CN2_sign => VN_sign_out(6470),
        VN2CN3_sign => VN_sign_out(6471),
        VN2CN4_sign => VN_sign_out(6472),
        VN2CN5_sign => VN_sign_out(6473),
        codeword => codeword(1078),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1079 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6479 downto 6474),
        Din0 => VN1079_in0,
        Din1 => VN1079_in1,
        Din2 => VN1079_in2,
        Din3 => VN1079_in3,
        Din4 => VN1079_in4,
        Din5 => VN1079_in5,
        VN2CN0_bit => VN_data_out(6474),
        VN2CN1_bit => VN_data_out(6475),
        VN2CN2_bit => VN_data_out(6476),
        VN2CN3_bit => VN_data_out(6477),
        VN2CN4_bit => VN_data_out(6478),
        VN2CN5_bit => VN_data_out(6479),
        VN2CN0_sign => VN_sign_out(6474),
        VN2CN1_sign => VN_sign_out(6475),
        VN2CN2_sign => VN_sign_out(6476),
        VN2CN3_sign => VN_sign_out(6477),
        VN2CN4_sign => VN_sign_out(6478),
        VN2CN5_sign => VN_sign_out(6479),
        codeword => codeword(1079),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1080 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6485 downto 6480),
        Din0 => VN1080_in0,
        Din1 => VN1080_in1,
        Din2 => VN1080_in2,
        Din3 => VN1080_in3,
        Din4 => VN1080_in4,
        Din5 => VN1080_in5,
        VN2CN0_bit => VN_data_out(6480),
        VN2CN1_bit => VN_data_out(6481),
        VN2CN2_bit => VN_data_out(6482),
        VN2CN3_bit => VN_data_out(6483),
        VN2CN4_bit => VN_data_out(6484),
        VN2CN5_bit => VN_data_out(6485),
        VN2CN0_sign => VN_sign_out(6480),
        VN2CN1_sign => VN_sign_out(6481),
        VN2CN2_sign => VN_sign_out(6482),
        VN2CN3_sign => VN_sign_out(6483),
        VN2CN4_sign => VN_sign_out(6484),
        VN2CN5_sign => VN_sign_out(6485),
        codeword => codeword(1080),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1081 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6491 downto 6486),
        Din0 => VN1081_in0,
        Din1 => VN1081_in1,
        Din2 => VN1081_in2,
        Din3 => VN1081_in3,
        Din4 => VN1081_in4,
        Din5 => VN1081_in5,
        VN2CN0_bit => VN_data_out(6486),
        VN2CN1_bit => VN_data_out(6487),
        VN2CN2_bit => VN_data_out(6488),
        VN2CN3_bit => VN_data_out(6489),
        VN2CN4_bit => VN_data_out(6490),
        VN2CN5_bit => VN_data_out(6491),
        VN2CN0_sign => VN_sign_out(6486),
        VN2CN1_sign => VN_sign_out(6487),
        VN2CN2_sign => VN_sign_out(6488),
        VN2CN3_sign => VN_sign_out(6489),
        VN2CN4_sign => VN_sign_out(6490),
        VN2CN5_sign => VN_sign_out(6491),
        codeword => codeword(1081),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1082 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6497 downto 6492),
        Din0 => VN1082_in0,
        Din1 => VN1082_in1,
        Din2 => VN1082_in2,
        Din3 => VN1082_in3,
        Din4 => VN1082_in4,
        Din5 => VN1082_in5,
        VN2CN0_bit => VN_data_out(6492),
        VN2CN1_bit => VN_data_out(6493),
        VN2CN2_bit => VN_data_out(6494),
        VN2CN3_bit => VN_data_out(6495),
        VN2CN4_bit => VN_data_out(6496),
        VN2CN5_bit => VN_data_out(6497),
        VN2CN0_sign => VN_sign_out(6492),
        VN2CN1_sign => VN_sign_out(6493),
        VN2CN2_sign => VN_sign_out(6494),
        VN2CN3_sign => VN_sign_out(6495),
        VN2CN4_sign => VN_sign_out(6496),
        VN2CN5_sign => VN_sign_out(6497),
        codeword => codeword(1082),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1083 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6503 downto 6498),
        Din0 => VN1083_in0,
        Din1 => VN1083_in1,
        Din2 => VN1083_in2,
        Din3 => VN1083_in3,
        Din4 => VN1083_in4,
        Din5 => VN1083_in5,
        VN2CN0_bit => VN_data_out(6498),
        VN2CN1_bit => VN_data_out(6499),
        VN2CN2_bit => VN_data_out(6500),
        VN2CN3_bit => VN_data_out(6501),
        VN2CN4_bit => VN_data_out(6502),
        VN2CN5_bit => VN_data_out(6503),
        VN2CN0_sign => VN_sign_out(6498),
        VN2CN1_sign => VN_sign_out(6499),
        VN2CN2_sign => VN_sign_out(6500),
        VN2CN3_sign => VN_sign_out(6501),
        VN2CN4_sign => VN_sign_out(6502),
        VN2CN5_sign => VN_sign_out(6503),
        codeword => codeword(1083),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1084 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6509 downto 6504),
        Din0 => VN1084_in0,
        Din1 => VN1084_in1,
        Din2 => VN1084_in2,
        Din3 => VN1084_in3,
        Din4 => VN1084_in4,
        Din5 => VN1084_in5,
        VN2CN0_bit => VN_data_out(6504),
        VN2CN1_bit => VN_data_out(6505),
        VN2CN2_bit => VN_data_out(6506),
        VN2CN3_bit => VN_data_out(6507),
        VN2CN4_bit => VN_data_out(6508),
        VN2CN5_bit => VN_data_out(6509),
        VN2CN0_sign => VN_sign_out(6504),
        VN2CN1_sign => VN_sign_out(6505),
        VN2CN2_sign => VN_sign_out(6506),
        VN2CN3_sign => VN_sign_out(6507),
        VN2CN4_sign => VN_sign_out(6508),
        VN2CN5_sign => VN_sign_out(6509),
        codeword => codeword(1084),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1085 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6515 downto 6510),
        Din0 => VN1085_in0,
        Din1 => VN1085_in1,
        Din2 => VN1085_in2,
        Din3 => VN1085_in3,
        Din4 => VN1085_in4,
        Din5 => VN1085_in5,
        VN2CN0_bit => VN_data_out(6510),
        VN2CN1_bit => VN_data_out(6511),
        VN2CN2_bit => VN_data_out(6512),
        VN2CN3_bit => VN_data_out(6513),
        VN2CN4_bit => VN_data_out(6514),
        VN2CN5_bit => VN_data_out(6515),
        VN2CN0_sign => VN_sign_out(6510),
        VN2CN1_sign => VN_sign_out(6511),
        VN2CN2_sign => VN_sign_out(6512),
        VN2CN3_sign => VN_sign_out(6513),
        VN2CN4_sign => VN_sign_out(6514),
        VN2CN5_sign => VN_sign_out(6515),
        codeword => codeword(1085),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1086 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6521 downto 6516),
        Din0 => VN1086_in0,
        Din1 => VN1086_in1,
        Din2 => VN1086_in2,
        Din3 => VN1086_in3,
        Din4 => VN1086_in4,
        Din5 => VN1086_in5,
        VN2CN0_bit => VN_data_out(6516),
        VN2CN1_bit => VN_data_out(6517),
        VN2CN2_bit => VN_data_out(6518),
        VN2CN3_bit => VN_data_out(6519),
        VN2CN4_bit => VN_data_out(6520),
        VN2CN5_bit => VN_data_out(6521),
        VN2CN0_sign => VN_sign_out(6516),
        VN2CN1_sign => VN_sign_out(6517),
        VN2CN2_sign => VN_sign_out(6518),
        VN2CN3_sign => VN_sign_out(6519),
        VN2CN4_sign => VN_sign_out(6520),
        VN2CN5_sign => VN_sign_out(6521),
        codeword => codeword(1086),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1087 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6527 downto 6522),
        Din0 => VN1087_in0,
        Din1 => VN1087_in1,
        Din2 => VN1087_in2,
        Din3 => VN1087_in3,
        Din4 => VN1087_in4,
        Din5 => VN1087_in5,
        VN2CN0_bit => VN_data_out(6522),
        VN2CN1_bit => VN_data_out(6523),
        VN2CN2_bit => VN_data_out(6524),
        VN2CN3_bit => VN_data_out(6525),
        VN2CN4_bit => VN_data_out(6526),
        VN2CN5_bit => VN_data_out(6527),
        VN2CN0_sign => VN_sign_out(6522),
        VN2CN1_sign => VN_sign_out(6523),
        VN2CN2_sign => VN_sign_out(6524),
        VN2CN3_sign => VN_sign_out(6525),
        VN2CN4_sign => VN_sign_out(6526),
        VN2CN5_sign => VN_sign_out(6527),
        codeword => codeword(1087),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1088 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6533 downto 6528),
        Din0 => VN1088_in0,
        Din1 => VN1088_in1,
        Din2 => VN1088_in2,
        Din3 => VN1088_in3,
        Din4 => VN1088_in4,
        Din5 => VN1088_in5,
        VN2CN0_bit => VN_data_out(6528),
        VN2CN1_bit => VN_data_out(6529),
        VN2CN2_bit => VN_data_out(6530),
        VN2CN3_bit => VN_data_out(6531),
        VN2CN4_bit => VN_data_out(6532),
        VN2CN5_bit => VN_data_out(6533),
        VN2CN0_sign => VN_sign_out(6528),
        VN2CN1_sign => VN_sign_out(6529),
        VN2CN2_sign => VN_sign_out(6530),
        VN2CN3_sign => VN_sign_out(6531),
        VN2CN4_sign => VN_sign_out(6532),
        VN2CN5_sign => VN_sign_out(6533),
        codeword => codeword(1088),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1089 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6539 downto 6534),
        Din0 => VN1089_in0,
        Din1 => VN1089_in1,
        Din2 => VN1089_in2,
        Din3 => VN1089_in3,
        Din4 => VN1089_in4,
        Din5 => VN1089_in5,
        VN2CN0_bit => VN_data_out(6534),
        VN2CN1_bit => VN_data_out(6535),
        VN2CN2_bit => VN_data_out(6536),
        VN2CN3_bit => VN_data_out(6537),
        VN2CN4_bit => VN_data_out(6538),
        VN2CN5_bit => VN_data_out(6539),
        VN2CN0_sign => VN_sign_out(6534),
        VN2CN1_sign => VN_sign_out(6535),
        VN2CN2_sign => VN_sign_out(6536),
        VN2CN3_sign => VN_sign_out(6537),
        VN2CN4_sign => VN_sign_out(6538),
        VN2CN5_sign => VN_sign_out(6539),
        codeword => codeword(1089),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1090 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6545 downto 6540),
        Din0 => VN1090_in0,
        Din1 => VN1090_in1,
        Din2 => VN1090_in2,
        Din3 => VN1090_in3,
        Din4 => VN1090_in4,
        Din5 => VN1090_in5,
        VN2CN0_bit => VN_data_out(6540),
        VN2CN1_bit => VN_data_out(6541),
        VN2CN2_bit => VN_data_out(6542),
        VN2CN3_bit => VN_data_out(6543),
        VN2CN4_bit => VN_data_out(6544),
        VN2CN5_bit => VN_data_out(6545),
        VN2CN0_sign => VN_sign_out(6540),
        VN2CN1_sign => VN_sign_out(6541),
        VN2CN2_sign => VN_sign_out(6542),
        VN2CN3_sign => VN_sign_out(6543),
        VN2CN4_sign => VN_sign_out(6544),
        VN2CN5_sign => VN_sign_out(6545),
        codeword => codeword(1090),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1091 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6551 downto 6546),
        Din0 => VN1091_in0,
        Din1 => VN1091_in1,
        Din2 => VN1091_in2,
        Din3 => VN1091_in3,
        Din4 => VN1091_in4,
        Din5 => VN1091_in5,
        VN2CN0_bit => VN_data_out(6546),
        VN2CN1_bit => VN_data_out(6547),
        VN2CN2_bit => VN_data_out(6548),
        VN2CN3_bit => VN_data_out(6549),
        VN2CN4_bit => VN_data_out(6550),
        VN2CN5_bit => VN_data_out(6551),
        VN2CN0_sign => VN_sign_out(6546),
        VN2CN1_sign => VN_sign_out(6547),
        VN2CN2_sign => VN_sign_out(6548),
        VN2CN3_sign => VN_sign_out(6549),
        VN2CN4_sign => VN_sign_out(6550),
        VN2CN5_sign => VN_sign_out(6551),
        codeword => codeword(1091),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1092 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6557 downto 6552),
        Din0 => VN1092_in0,
        Din1 => VN1092_in1,
        Din2 => VN1092_in2,
        Din3 => VN1092_in3,
        Din4 => VN1092_in4,
        Din5 => VN1092_in5,
        VN2CN0_bit => VN_data_out(6552),
        VN2CN1_bit => VN_data_out(6553),
        VN2CN2_bit => VN_data_out(6554),
        VN2CN3_bit => VN_data_out(6555),
        VN2CN4_bit => VN_data_out(6556),
        VN2CN5_bit => VN_data_out(6557),
        VN2CN0_sign => VN_sign_out(6552),
        VN2CN1_sign => VN_sign_out(6553),
        VN2CN2_sign => VN_sign_out(6554),
        VN2CN3_sign => VN_sign_out(6555),
        VN2CN4_sign => VN_sign_out(6556),
        VN2CN5_sign => VN_sign_out(6557),
        codeword => codeword(1092),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1093 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6563 downto 6558),
        Din0 => VN1093_in0,
        Din1 => VN1093_in1,
        Din2 => VN1093_in2,
        Din3 => VN1093_in3,
        Din4 => VN1093_in4,
        Din5 => VN1093_in5,
        VN2CN0_bit => VN_data_out(6558),
        VN2CN1_bit => VN_data_out(6559),
        VN2CN2_bit => VN_data_out(6560),
        VN2CN3_bit => VN_data_out(6561),
        VN2CN4_bit => VN_data_out(6562),
        VN2CN5_bit => VN_data_out(6563),
        VN2CN0_sign => VN_sign_out(6558),
        VN2CN1_sign => VN_sign_out(6559),
        VN2CN2_sign => VN_sign_out(6560),
        VN2CN3_sign => VN_sign_out(6561),
        VN2CN4_sign => VN_sign_out(6562),
        VN2CN5_sign => VN_sign_out(6563),
        codeword => codeword(1093),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1094 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6569 downto 6564),
        Din0 => VN1094_in0,
        Din1 => VN1094_in1,
        Din2 => VN1094_in2,
        Din3 => VN1094_in3,
        Din4 => VN1094_in4,
        Din5 => VN1094_in5,
        VN2CN0_bit => VN_data_out(6564),
        VN2CN1_bit => VN_data_out(6565),
        VN2CN2_bit => VN_data_out(6566),
        VN2CN3_bit => VN_data_out(6567),
        VN2CN4_bit => VN_data_out(6568),
        VN2CN5_bit => VN_data_out(6569),
        VN2CN0_sign => VN_sign_out(6564),
        VN2CN1_sign => VN_sign_out(6565),
        VN2CN2_sign => VN_sign_out(6566),
        VN2CN3_sign => VN_sign_out(6567),
        VN2CN4_sign => VN_sign_out(6568),
        VN2CN5_sign => VN_sign_out(6569),
        codeword => codeword(1094),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1095 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6575 downto 6570),
        Din0 => VN1095_in0,
        Din1 => VN1095_in1,
        Din2 => VN1095_in2,
        Din3 => VN1095_in3,
        Din4 => VN1095_in4,
        Din5 => VN1095_in5,
        VN2CN0_bit => VN_data_out(6570),
        VN2CN1_bit => VN_data_out(6571),
        VN2CN2_bit => VN_data_out(6572),
        VN2CN3_bit => VN_data_out(6573),
        VN2CN4_bit => VN_data_out(6574),
        VN2CN5_bit => VN_data_out(6575),
        VN2CN0_sign => VN_sign_out(6570),
        VN2CN1_sign => VN_sign_out(6571),
        VN2CN2_sign => VN_sign_out(6572),
        VN2CN3_sign => VN_sign_out(6573),
        VN2CN4_sign => VN_sign_out(6574),
        VN2CN5_sign => VN_sign_out(6575),
        codeword => codeword(1095),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1096 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6581 downto 6576),
        Din0 => VN1096_in0,
        Din1 => VN1096_in1,
        Din2 => VN1096_in2,
        Din3 => VN1096_in3,
        Din4 => VN1096_in4,
        Din5 => VN1096_in5,
        VN2CN0_bit => VN_data_out(6576),
        VN2CN1_bit => VN_data_out(6577),
        VN2CN2_bit => VN_data_out(6578),
        VN2CN3_bit => VN_data_out(6579),
        VN2CN4_bit => VN_data_out(6580),
        VN2CN5_bit => VN_data_out(6581),
        VN2CN0_sign => VN_sign_out(6576),
        VN2CN1_sign => VN_sign_out(6577),
        VN2CN2_sign => VN_sign_out(6578),
        VN2CN3_sign => VN_sign_out(6579),
        VN2CN4_sign => VN_sign_out(6580),
        VN2CN5_sign => VN_sign_out(6581),
        codeword => codeword(1096),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1097 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6587 downto 6582),
        Din0 => VN1097_in0,
        Din1 => VN1097_in1,
        Din2 => VN1097_in2,
        Din3 => VN1097_in3,
        Din4 => VN1097_in4,
        Din5 => VN1097_in5,
        VN2CN0_bit => VN_data_out(6582),
        VN2CN1_bit => VN_data_out(6583),
        VN2CN2_bit => VN_data_out(6584),
        VN2CN3_bit => VN_data_out(6585),
        VN2CN4_bit => VN_data_out(6586),
        VN2CN5_bit => VN_data_out(6587),
        VN2CN0_sign => VN_sign_out(6582),
        VN2CN1_sign => VN_sign_out(6583),
        VN2CN2_sign => VN_sign_out(6584),
        VN2CN3_sign => VN_sign_out(6585),
        VN2CN4_sign => VN_sign_out(6586),
        VN2CN5_sign => VN_sign_out(6587),
        codeword => codeword(1097),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1098 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6593 downto 6588),
        Din0 => VN1098_in0,
        Din1 => VN1098_in1,
        Din2 => VN1098_in2,
        Din3 => VN1098_in3,
        Din4 => VN1098_in4,
        Din5 => VN1098_in5,
        VN2CN0_bit => VN_data_out(6588),
        VN2CN1_bit => VN_data_out(6589),
        VN2CN2_bit => VN_data_out(6590),
        VN2CN3_bit => VN_data_out(6591),
        VN2CN4_bit => VN_data_out(6592),
        VN2CN5_bit => VN_data_out(6593),
        VN2CN0_sign => VN_sign_out(6588),
        VN2CN1_sign => VN_sign_out(6589),
        VN2CN2_sign => VN_sign_out(6590),
        VN2CN3_sign => VN_sign_out(6591),
        VN2CN4_sign => VN_sign_out(6592),
        VN2CN5_sign => VN_sign_out(6593),
        codeword => codeword(1098),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1099 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6599 downto 6594),
        Din0 => VN1099_in0,
        Din1 => VN1099_in1,
        Din2 => VN1099_in2,
        Din3 => VN1099_in3,
        Din4 => VN1099_in4,
        Din5 => VN1099_in5,
        VN2CN0_bit => VN_data_out(6594),
        VN2CN1_bit => VN_data_out(6595),
        VN2CN2_bit => VN_data_out(6596),
        VN2CN3_bit => VN_data_out(6597),
        VN2CN4_bit => VN_data_out(6598),
        VN2CN5_bit => VN_data_out(6599),
        VN2CN0_sign => VN_sign_out(6594),
        VN2CN1_sign => VN_sign_out(6595),
        VN2CN2_sign => VN_sign_out(6596),
        VN2CN3_sign => VN_sign_out(6597),
        VN2CN4_sign => VN_sign_out(6598),
        VN2CN5_sign => VN_sign_out(6599),
        codeword => codeword(1099),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1100 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6605 downto 6600),
        Din0 => VN1100_in0,
        Din1 => VN1100_in1,
        Din2 => VN1100_in2,
        Din3 => VN1100_in3,
        Din4 => VN1100_in4,
        Din5 => VN1100_in5,
        VN2CN0_bit => VN_data_out(6600),
        VN2CN1_bit => VN_data_out(6601),
        VN2CN2_bit => VN_data_out(6602),
        VN2CN3_bit => VN_data_out(6603),
        VN2CN4_bit => VN_data_out(6604),
        VN2CN5_bit => VN_data_out(6605),
        VN2CN0_sign => VN_sign_out(6600),
        VN2CN1_sign => VN_sign_out(6601),
        VN2CN2_sign => VN_sign_out(6602),
        VN2CN3_sign => VN_sign_out(6603),
        VN2CN4_sign => VN_sign_out(6604),
        VN2CN5_sign => VN_sign_out(6605),
        codeword => codeword(1100),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1101 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6611 downto 6606),
        Din0 => VN1101_in0,
        Din1 => VN1101_in1,
        Din2 => VN1101_in2,
        Din3 => VN1101_in3,
        Din4 => VN1101_in4,
        Din5 => VN1101_in5,
        VN2CN0_bit => VN_data_out(6606),
        VN2CN1_bit => VN_data_out(6607),
        VN2CN2_bit => VN_data_out(6608),
        VN2CN3_bit => VN_data_out(6609),
        VN2CN4_bit => VN_data_out(6610),
        VN2CN5_bit => VN_data_out(6611),
        VN2CN0_sign => VN_sign_out(6606),
        VN2CN1_sign => VN_sign_out(6607),
        VN2CN2_sign => VN_sign_out(6608),
        VN2CN3_sign => VN_sign_out(6609),
        VN2CN4_sign => VN_sign_out(6610),
        VN2CN5_sign => VN_sign_out(6611),
        codeword => codeword(1101),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1102 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6617 downto 6612),
        Din0 => VN1102_in0,
        Din1 => VN1102_in1,
        Din2 => VN1102_in2,
        Din3 => VN1102_in3,
        Din4 => VN1102_in4,
        Din5 => VN1102_in5,
        VN2CN0_bit => VN_data_out(6612),
        VN2CN1_bit => VN_data_out(6613),
        VN2CN2_bit => VN_data_out(6614),
        VN2CN3_bit => VN_data_out(6615),
        VN2CN4_bit => VN_data_out(6616),
        VN2CN5_bit => VN_data_out(6617),
        VN2CN0_sign => VN_sign_out(6612),
        VN2CN1_sign => VN_sign_out(6613),
        VN2CN2_sign => VN_sign_out(6614),
        VN2CN3_sign => VN_sign_out(6615),
        VN2CN4_sign => VN_sign_out(6616),
        VN2CN5_sign => VN_sign_out(6617),
        codeword => codeword(1102),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1103 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6623 downto 6618),
        Din0 => VN1103_in0,
        Din1 => VN1103_in1,
        Din2 => VN1103_in2,
        Din3 => VN1103_in3,
        Din4 => VN1103_in4,
        Din5 => VN1103_in5,
        VN2CN0_bit => VN_data_out(6618),
        VN2CN1_bit => VN_data_out(6619),
        VN2CN2_bit => VN_data_out(6620),
        VN2CN3_bit => VN_data_out(6621),
        VN2CN4_bit => VN_data_out(6622),
        VN2CN5_bit => VN_data_out(6623),
        VN2CN0_sign => VN_sign_out(6618),
        VN2CN1_sign => VN_sign_out(6619),
        VN2CN2_sign => VN_sign_out(6620),
        VN2CN3_sign => VN_sign_out(6621),
        VN2CN4_sign => VN_sign_out(6622),
        VN2CN5_sign => VN_sign_out(6623),
        codeword => codeword(1103),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1104 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6629 downto 6624),
        Din0 => VN1104_in0,
        Din1 => VN1104_in1,
        Din2 => VN1104_in2,
        Din3 => VN1104_in3,
        Din4 => VN1104_in4,
        Din5 => VN1104_in5,
        VN2CN0_bit => VN_data_out(6624),
        VN2CN1_bit => VN_data_out(6625),
        VN2CN2_bit => VN_data_out(6626),
        VN2CN3_bit => VN_data_out(6627),
        VN2CN4_bit => VN_data_out(6628),
        VN2CN5_bit => VN_data_out(6629),
        VN2CN0_sign => VN_sign_out(6624),
        VN2CN1_sign => VN_sign_out(6625),
        VN2CN2_sign => VN_sign_out(6626),
        VN2CN3_sign => VN_sign_out(6627),
        VN2CN4_sign => VN_sign_out(6628),
        VN2CN5_sign => VN_sign_out(6629),
        codeword => codeword(1104),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1105 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6635 downto 6630),
        Din0 => VN1105_in0,
        Din1 => VN1105_in1,
        Din2 => VN1105_in2,
        Din3 => VN1105_in3,
        Din4 => VN1105_in4,
        Din5 => VN1105_in5,
        VN2CN0_bit => VN_data_out(6630),
        VN2CN1_bit => VN_data_out(6631),
        VN2CN2_bit => VN_data_out(6632),
        VN2CN3_bit => VN_data_out(6633),
        VN2CN4_bit => VN_data_out(6634),
        VN2CN5_bit => VN_data_out(6635),
        VN2CN0_sign => VN_sign_out(6630),
        VN2CN1_sign => VN_sign_out(6631),
        VN2CN2_sign => VN_sign_out(6632),
        VN2CN3_sign => VN_sign_out(6633),
        VN2CN4_sign => VN_sign_out(6634),
        VN2CN5_sign => VN_sign_out(6635),
        codeword => codeword(1105),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1106 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6641 downto 6636),
        Din0 => VN1106_in0,
        Din1 => VN1106_in1,
        Din2 => VN1106_in2,
        Din3 => VN1106_in3,
        Din4 => VN1106_in4,
        Din5 => VN1106_in5,
        VN2CN0_bit => VN_data_out(6636),
        VN2CN1_bit => VN_data_out(6637),
        VN2CN2_bit => VN_data_out(6638),
        VN2CN3_bit => VN_data_out(6639),
        VN2CN4_bit => VN_data_out(6640),
        VN2CN5_bit => VN_data_out(6641),
        VN2CN0_sign => VN_sign_out(6636),
        VN2CN1_sign => VN_sign_out(6637),
        VN2CN2_sign => VN_sign_out(6638),
        VN2CN3_sign => VN_sign_out(6639),
        VN2CN4_sign => VN_sign_out(6640),
        VN2CN5_sign => VN_sign_out(6641),
        codeword => codeword(1106),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1107 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6647 downto 6642),
        Din0 => VN1107_in0,
        Din1 => VN1107_in1,
        Din2 => VN1107_in2,
        Din3 => VN1107_in3,
        Din4 => VN1107_in4,
        Din5 => VN1107_in5,
        VN2CN0_bit => VN_data_out(6642),
        VN2CN1_bit => VN_data_out(6643),
        VN2CN2_bit => VN_data_out(6644),
        VN2CN3_bit => VN_data_out(6645),
        VN2CN4_bit => VN_data_out(6646),
        VN2CN5_bit => VN_data_out(6647),
        VN2CN0_sign => VN_sign_out(6642),
        VN2CN1_sign => VN_sign_out(6643),
        VN2CN2_sign => VN_sign_out(6644),
        VN2CN3_sign => VN_sign_out(6645),
        VN2CN4_sign => VN_sign_out(6646),
        VN2CN5_sign => VN_sign_out(6647),
        codeword => codeword(1107),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1108 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6653 downto 6648),
        Din0 => VN1108_in0,
        Din1 => VN1108_in1,
        Din2 => VN1108_in2,
        Din3 => VN1108_in3,
        Din4 => VN1108_in4,
        Din5 => VN1108_in5,
        VN2CN0_bit => VN_data_out(6648),
        VN2CN1_bit => VN_data_out(6649),
        VN2CN2_bit => VN_data_out(6650),
        VN2CN3_bit => VN_data_out(6651),
        VN2CN4_bit => VN_data_out(6652),
        VN2CN5_bit => VN_data_out(6653),
        VN2CN0_sign => VN_sign_out(6648),
        VN2CN1_sign => VN_sign_out(6649),
        VN2CN2_sign => VN_sign_out(6650),
        VN2CN3_sign => VN_sign_out(6651),
        VN2CN4_sign => VN_sign_out(6652),
        VN2CN5_sign => VN_sign_out(6653),
        codeword => codeword(1108),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1109 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6659 downto 6654),
        Din0 => VN1109_in0,
        Din1 => VN1109_in1,
        Din2 => VN1109_in2,
        Din3 => VN1109_in3,
        Din4 => VN1109_in4,
        Din5 => VN1109_in5,
        VN2CN0_bit => VN_data_out(6654),
        VN2CN1_bit => VN_data_out(6655),
        VN2CN2_bit => VN_data_out(6656),
        VN2CN3_bit => VN_data_out(6657),
        VN2CN4_bit => VN_data_out(6658),
        VN2CN5_bit => VN_data_out(6659),
        VN2CN0_sign => VN_sign_out(6654),
        VN2CN1_sign => VN_sign_out(6655),
        VN2CN2_sign => VN_sign_out(6656),
        VN2CN3_sign => VN_sign_out(6657),
        VN2CN4_sign => VN_sign_out(6658),
        VN2CN5_sign => VN_sign_out(6659),
        codeword => codeword(1109),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1110 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6665 downto 6660),
        Din0 => VN1110_in0,
        Din1 => VN1110_in1,
        Din2 => VN1110_in2,
        Din3 => VN1110_in3,
        Din4 => VN1110_in4,
        Din5 => VN1110_in5,
        VN2CN0_bit => VN_data_out(6660),
        VN2CN1_bit => VN_data_out(6661),
        VN2CN2_bit => VN_data_out(6662),
        VN2CN3_bit => VN_data_out(6663),
        VN2CN4_bit => VN_data_out(6664),
        VN2CN5_bit => VN_data_out(6665),
        VN2CN0_sign => VN_sign_out(6660),
        VN2CN1_sign => VN_sign_out(6661),
        VN2CN2_sign => VN_sign_out(6662),
        VN2CN3_sign => VN_sign_out(6663),
        VN2CN4_sign => VN_sign_out(6664),
        VN2CN5_sign => VN_sign_out(6665),
        codeword => codeword(1110),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1111 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6671 downto 6666),
        Din0 => VN1111_in0,
        Din1 => VN1111_in1,
        Din2 => VN1111_in2,
        Din3 => VN1111_in3,
        Din4 => VN1111_in4,
        Din5 => VN1111_in5,
        VN2CN0_bit => VN_data_out(6666),
        VN2CN1_bit => VN_data_out(6667),
        VN2CN2_bit => VN_data_out(6668),
        VN2CN3_bit => VN_data_out(6669),
        VN2CN4_bit => VN_data_out(6670),
        VN2CN5_bit => VN_data_out(6671),
        VN2CN0_sign => VN_sign_out(6666),
        VN2CN1_sign => VN_sign_out(6667),
        VN2CN2_sign => VN_sign_out(6668),
        VN2CN3_sign => VN_sign_out(6669),
        VN2CN4_sign => VN_sign_out(6670),
        VN2CN5_sign => VN_sign_out(6671),
        codeword => codeword(1111),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1112 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6677 downto 6672),
        Din0 => VN1112_in0,
        Din1 => VN1112_in1,
        Din2 => VN1112_in2,
        Din3 => VN1112_in3,
        Din4 => VN1112_in4,
        Din5 => VN1112_in5,
        VN2CN0_bit => VN_data_out(6672),
        VN2CN1_bit => VN_data_out(6673),
        VN2CN2_bit => VN_data_out(6674),
        VN2CN3_bit => VN_data_out(6675),
        VN2CN4_bit => VN_data_out(6676),
        VN2CN5_bit => VN_data_out(6677),
        VN2CN0_sign => VN_sign_out(6672),
        VN2CN1_sign => VN_sign_out(6673),
        VN2CN2_sign => VN_sign_out(6674),
        VN2CN3_sign => VN_sign_out(6675),
        VN2CN4_sign => VN_sign_out(6676),
        VN2CN5_sign => VN_sign_out(6677),
        codeword => codeword(1112),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1113 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6683 downto 6678),
        Din0 => VN1113_in0,
        Din1 => VN1113_in1,
        Din2 => VN1113_in2,
        Din3 => VN1113_in3,
        Din4 => VN1113_in4,
        Din5 => VN1113_in5,
        VN2CN0_bit => VN_data_out(6678),
        VN2CN1_bit => VN_data_out(6679),
        VN2CN2_bit => VN_data_out(6680),
        VN2CN3_bit => VN_data_out(6681),
        VN2CN4_bit => VN_data_out(6682),
        VN2CN5_bit => VN_data_out(6683),
        VN2CN0_sign => VN_sign_out(6678),
        VN2CN1_sign => VN_sign_out(6679),
        VN2CN2_sign => VN_sign_out(6680),
        VN2CN3_sign => VN_sign_out(6681),
        VN2CN4_sign => VN_sign_out(6682),
        VN2CN5_sign => VN_sign_out(6683),
        codeword => codeword(1113),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1114 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6689 downto 6684),
        Din0 => VN1114_in0,
        Din1 => VN1114_in1,
        Din2 => VN1114_in2,
        Din3 => VN1114_in3,
        Din4 => VN1114_in4,
        Din5 => VN1114_in5,
        VN2CN0_bit => VN_data_out(6684),
        VN2CN1_bit => VN_data_out(6685),
        VN2CN2_bit => VN_data_out(6686),
        VN2CN3_bit => VN_data_out(6687),
        VN2CN4_bit => VN_data_out(6688),
        VN2CN5_bit => VN_data_out(6689),
        VN2CN0_sign => VN_sign_out(6684),
        VN2CN1_sign => VN_sign_out(6685),
        VN2CN2_sign => VN_sign_out(6686),
        VN2CN3_sign => VN_sign_out(6687),
        VN2CN4_sign => VN_sign_out(6688),
        VN2CN5_sign => VN_sign_out(6689),
        codeword => codeword(1114),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1115 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6695 downto 6690),
        Din0 => VN1115_in0,
        Din1 => VN1115_in1,
        Din2 => VN1115_in2,
        Din3 => VN1115_in3,
        Din4 => VN1115_in4,
        Din5 => VN1115_in5,
        VN2CN0_bit => VN_data_out(6690),
        VN2CN1_bit => VN_data_out(6691),
        VN2CN2_bit => VN_data_out(6692),
        VN2CN3_bit => VN_data_out(6693),
        VN2CN4_bit => VN_data_out(6694),
        VN2CN5_bit => VN_data_out(6695),
        VN2CN0_sign => VN_sign_out(6690),
        VN2CN1_sign => VN_sign_out(6691),
        VN2CN2_sign => VN_sign_out(6692),
        VN2CN3_sign => VN_sign_out(6693),
        VN2CN4_sign => VN_sign_out(6694),
        VN2CN5_sign => VN_sign_out(6695),
        codeword => codeword(1115),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1116 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6701 downto 6696),
        Din0 => VN1116_in0,
        Din1 => VN1116_in1,
        Din2 => VN1116_in2,
        Din3 => VN1116_in3,
        Din4 => VN1116_in4,
        Din5 => VN1116_in5,
        VN2CN0_bit => VN_data_out(6696),
        VN2CN1_bit => VN_data_out(6697),
        VN2CN2_bit => VN_data_out(6698),
        VN2CN3_bit => VN_data_out(6699),
        VN2CN4_bit => VN_data_out(6700),
        VN2CN5_bit => VN_data_out(6701),
        VN2CN0_sign => VN_sign_out(6696),
        VN2CN1_sign => VN_sign_out(6697),
        VN2CN2_sign => VN_sign_out(6698),
        VN2CN3_sign => VN_sign_out(6699),
        VN2CN4_sign => VN_sign_out(6700),
        VN2CN5_sign => VN_sign_out(6701),
        codeword => codeword(1116),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1117 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6707 downto 6702),
        Din0 => VN1117_in0,
        Din1 => VN1117_in1,
        Din2 => VN1117_in2,
        Din3 => VN1117_in3,
        Din4 => VN1117_in4,
        Din5 => VN1117_in5,
        VN2CN0_bit => VN_data_out(6702),
        VN2CN1_bit => VN_data_out(6703),
        VN2CN2_bit => VN_data_out(6704),
        VN2CN3_bit => VN_data_out(6705),
        VN2CN4_bit => VN_data_out(6706),
        VN2CN5_bit => VN_data_out(6707),
        VN2CN0_sign => VN_sign_out(6702),
        VN2CN1_sign => VN_sign_out(6703),
        VN2CN2_sign => VN_sign_out(6704),
        VN2CN3_sign => VN_sign_out(6705),
        VN2CN4_sign => VN_sign_out(6706),
        VN2CN5_sign => VN_sign_out(6707),
        codeword => codeword(1117),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1118 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6713 downto 6708),
        Din0 => VN1118_in0,
        Din1 => VN1118_in1,
        Din2 => VN1118_in2,
        Din3 => VN1118_in3,
        Din4 => VN1118_in4,
        Din5 => VN1118_in5,
        VN2CN0_bit => VN_data_out(6708),
        VN2CN1_bit => VN_data_out(6709),
        VN2CN2_bit => VN_data_out(6710),
        VN2CN3_bit => VN_data_out(6711),
        VN2CN4_bit => VN_data_out(6712),
        VN2CN5_bit => VN_data_out(6713),
        VN2CN0_sign => VN_sign_out(6708),
        VN2CN1_sign => VN_sign_out(6709),
        VN2CN2_sign => VN_sign_out(6710),
        VN2CN3_sign => VN_sign_out(6711),
        VN2CN4_sign => VN_sign_out(6712),
        VN2CN5_sign => VN_sign_out(6713),
        codeword => codeword(1118),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1119 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6719 downto 6714),
        Din0 => VN1119_in0,
        Din1 => VN1119_in1,
        Din2 => VN1119_in2,
        Din3 => VN1119_in3,
        Din4 => VN1119_in4,
        Din5 => VN1119_in5,
        VN2CN0_bit => VN_data_out(6714),
        VN2CN1_bit => VN_data_out(6715),
        VN2CN2_bit => VN_data_out(6716),
        VN2CN3_bit => VN_data_out(6717),
        VN2CN4_bit => VN_data_out(6718),
        VN2CN5_bit => VN_data_out(6719),
        VN2CN0_sign => VN_sign_out(6714),
        VN2CN1_sign => VN_sign_out(6715),
        VN2CN2_sign => VN_sign_out(6716),
        VN2CN3_sign => VN_sign_out(6717),
        VN2CN4_sign => VN_sign_out(6718),
        VN2CN5_sign => VN_sign_out(6719),
        codeword => codeword(1119),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1120 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6725 downto 6720),
        Din0 => VN1120_in0,
        Din1 => VN1120_in1,
        Din2 => VN1120_in2,
        Din3 => VN1120_in3,
        Din4 => VN1120_in4,
        Din5 => VN1120_in5,
        VN2CN0_bit => VN_data_out(6720),
        VN2CN1_bit => VN_data_out(6721),
        VN2CN2_bit => VN_data_out(6722),
        VN2CN3_bit => VN_data_out(6723),
        VN2CN4_bit => VN_data_out(6724),
        VN2CN5_bit => VN_data_out(6725),
        VN2CN0_sign => VN_sign_out(6720),
        VN2CN1_sign => VN_sign_out(6721),
        VN2CN2_sign => VN_sign_out(6722),
        VN2CN3_sign => VN_sign_out(6723),
        VN2CN4_sign => VN_sign_out(6724),
        VN2CN5_sign => VN_sign_out(6725),
        codeword => codeword(1120),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1121 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6731 downto 6726),
        Din0 => VN1121_in0,
        Din1 => VN1121_in1,
        Din2 => VN1121_in2,
        Din3 => VN1121_in3,
        Din4 => VN1121_in4,
        Din5 => VN1121_in5,
        VN2CN0_bit => VN_data_out(6726),
        VN2CN1_bit => VN_data_out(6727),
        VN2CN2_bit => VN_data_out(6728),
        VN2CN3_bit => VN_data_out(6729),
        VN2CN4_bit => VN_data_out(6730),
        VN2CN5_bit => VN_data_out(6731),
        VN2CN0_sign => VN_sign_out(6726),
        VN2CN1_sign => VN_sign_out(6727),
        VN2CN2_sign => VN_sign_out(6728),
        VN2CN3_sign => VN_sign_out(6729),
        VN2CN4_sign => VN_sign_out(6730),
        VN2CN5_sign => VN_sign_out(6731),
        codeword => codeword(1121),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1122 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6737 downto 6732),
        Din0 => VN1122_in0,
        Din1 => VN1122_in1,
        Din2 => VN1122_in2,
        Din3 => VN1122_in3,
        Din4 => VN1122_in4,
        Din5 => VN1122_in5,
        VN2CN0_bit => VN_data_out(6732),
        VN2CN1_bit => VN_data_out(6733),
        VN2CN2_bit => VN_data_out(6734),
        VN2CN3_bit => VN_data_out(6735),
        VN2CN4_bit => VN_data_out(6736),
        VN2CN5_bit => VN_data_out(6737),
        VN2CN0_sign => VN_sign_out(6732),
        VN2CN1_sign => VN_sign_out(6733),
        VN2CN2_sign => VN_sign_out(6734),
        VN2CN3_sign => VN_sign_out(6735),
        VN2CN4_sign => VN_sign_out(6736),
        VN2CN5_sign => VN_sign_out(6737),
        codeword => codeword(1122),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1123 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6743 downto 6738),
        Din0 => VN1123_in0,
        Din1 => VN1123_in1,
        Din2 => VN1123_in2,
        Din3 => VN1123_in3,
        Din4 => VN1123_in4,
        Din5 => VN1123_in5,
        VN2CN0_bit => VN_data_out(6738),
        VN2CN1_bit => VN_data_out(6739),
        VN2CN2_bit => VN_data_out(6740),
        VN2CN3_bit => VN_data_out(6741),
        VN2CN4_bit => VN_data_out(6742),
        VN2CN5_bit => VN_data_out(6743),
        VN2CN0_sign => VN_sign_out(6738),
        VN2CN1_sign => VN_sign_out(6739),
        VN2CN2_sign => VN_sign_out(6740),
        VN2CN3_sign => VN_sign_out(6741),
        VN2CN4_sign => VN_sign_out(6742),
        VN2CN5_sign => VN_sign_out(6743),
        codeword => codeword(1123),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1124 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6749 downto 6744),
        Din0 => VN1124_in0,
        Din1 => VN1124_in1,
        Din2 => VN1124_in2,
        Din3 => VN1124_in3,
        Din4 => VN1124_in4,
        Din5 => VN1124_in5,
        VN2CN0_bit => VN_data_out(6744),
        VN2CN1_bit => VN_data_out(6745),
        VN2CN2_bit => VN_data_out(6746),
        VN2CN3_bit => VN_data_out(6747),
        VN2CN4_bit => VN_data_out(6748),
        VN2CN5_bit => VN_data_out(6749),
        VN2CN0_sign => VN_sign_out(6744),
        VN2CN1_sign => VN_sign_out(6745),
        VN2CN2_sign => VN_sign_out(6746),
        VN2CN3_sign => VN_sign_out(6747),
        VN2CN4_sign => VN_sign_out(6748),
        VN2CN5_sign => VN_sign_out(6749),
        codeword => codeword(1124),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1125 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6755 downto 6750),
        Din0 => VN1125_in0,
        Din1 => VN1125_in1,
        Din2 => VN1125_in2,
        Din3 => VN1125_in3,
        Din4 => VN1125_in4,
        Din5 => VN1125_in5,
        VN2CN0_bit => VN_data_out(6750),
        VN2CN1_bit => VN_data_out(6751),
        VN2CN2_bit => VN_data_out(6752),
        VN2CN3_bit => VN_data_out(6753),
        VN2CN4_bit => VN_data_out(6754),
        VN2CN5_bit => VN_data_out(6755),
        VN2CN0_sign => VN_sign_out(6750),
        VN2CN1_sign => VN_sign_out(6751),
        VN2CN2_sign => VN_sign_out(6752),
        VN2CN3_sign => VN_sign_out(6753),
        VN2CN4_sign => VN_sign_out(6754),
        VN2CN5_sign => VN_sign_out(6755),
        codeword => codeword(1125),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1126 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6761 downto 6756),
        Din0 => VN1126_in0,
        Din1 => VN1126_in1,
        Din2 => VN1126_in2,
        Din3 => VN1126_in3,
        Din4 => VN1126_in4,
        Din5 => VN1126_in5,
        VN2CN0_bit => VN_data_out(6756),
        VN2CN1_bit => VN_data_out(6757),
        VN2CN2_bit => VN_data_out(6758),
        VN2CN3_bit => VN_data_out(6759),
        VN2CN4_bit => VN_data_out(6760),
        VN2CN5_bit => VN_data_out(6761),
        VN2CN0_sign => VN_sign_out(6756),
        VN2CN1_sign => VN_sign_out(6757),
        VN2CN2_sign => VN_sign_out(6758),
        VN2CN3_sign => VN_sign_out(6759),
        VN2CN4_sign => VN_sign_out(6760),
        VN2CN5_sign => VN_sign_out(6761),
        codeword => codeword(1126),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1127 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6767 downto 6762),
        Din0 => VN1127_in0,
        Din1 => VN1127_in1,
        Din2 => VN1127_in2,
        Din3 => VN1127_in3,
        Din4 => VN1127_in4,
        Din5 => VN1127_in5,
        VN2CN0_bit => VN_data_out(6762),
        VN2CN1_bit => VN_data_out(6763),
        VN2CN2_bit => VN_data_out(6764),
        VN2CN3_bit => VN_data_out(6765),
        VN2CN4_bit => VN_data_out(6766),
        VN2CN5_bit => VN_data_out(6767),
        VN2CN0_sign => VN_sign_out(6762),
        VN2CN1_sign => VN_sign_out(6763),
        VN2CN2_sign => VN_sign_out(6764),
        VN2CN3_sign => VN_sign_out(6765),
        VN2CN4_sign => VN_sign_out(6766),
        VN2CN5_sign => VN_sign_out(6767),
        codeword => codeword(1127),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1128 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6773 downto 6768),
        Din0 => VN1128_in0,
        Din1 => VN1128_in1,
        Din2 => VN1128_in2,
        Din3 => VN1128_in3,
        Din4 => VN1128_in4,
        Din5 => VN1128_in5,
        VN2CN0_bit => VN_data_out(6768),
        VN2CN1_bit => VN_data_out(6769),
        VN2CN2_bit => VN_data_out(6770),
        VN2CN3_bit => VN_data_out(6771),
        VN2CN4_bit => VN_data_out(6772),
        VN2CN5_bit => VN_data_out(6773),
        VN2CN0_sign => VN_sign_out(6768),
        VN2CN1_sign => VN_sign_out(6769),
        VN2CN2_sign => VN_sign_out(6770),
        VN2CN3_sign => VN_sign_out(6771),
        VN2CN4_sign => VN_sign_out(6772),
        VN2CN5_sign => VN_sign_out(6773),
        codeword => codeword(1128),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1129 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6779 downto 6774),
        Din0 => VN1129_in0,
        Din1 => VN1129_in1,
        Din2 => VN1129_in2,
        Din3 => VN1129_in3,
        Din4 => VN1129_in4,
        Din5 => VN1129_in5,
        VN2CN0_bit => VN_data_out(6774),
        VN2CN1_bit => VN_data_out(6775),
        VN2CN2_bit => VN_data_out(6776),
        VN2CN3_bit => VN_data_out(6777),
        VN2CN4_bit => VN_data_out(6778),
        VN2CN5_bit => VN_data_out(6779),
        VN2CN0_sign => VN_sign_out(6774),
        VN2CN1_sign => VN_sign_out(6775),
        VN2CN2_sign => VN_sign_out(6776),
        VN2CN3_sign => VN_sign_out(6777),
        VN2CN4_sign => VN_sign_out(6778),
        VN2CN5_sign => VN_sign_out(6779),
        codeword => codeword(1129),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1130 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6785 downto 6780),
        Din0 => VN1130_in0,
        Din1 => VN1130_in1,
        Din2 => VN1130_in2,
        Din3 => VN1130_in3,
        Din4 => VN1130_in4,
        Din5 => VN1130_in5,
        VN2CN0_bit => VN_data_out(6780),
        VN2CN1_bit => VN_data_out(6781),
        VN2CN2_bit => VN_data_out(6782),
        VN2CN3_bit => VN_data_out(6783),
        VN2CN4_bit => VN_data_out(6784),
        VN2CN5_bit => VN_data_out(6785),
        VN2CN0_sign => VN_sign_out(6780),
        VN2CN1_sign => VN_sign_out(6781),
        VN2CN2_sign => VN_sign_out(6782),
        VN2CN3_sign => VN_sign_out(6783),
        VN2CN4_sign => VN_sign_out(6784),
        VN2CN5_sign => VN_sign_out(6785),
        codeword => codeword(1130),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1131 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6791 downto 6786),
        Din0 => VN1131_in0,
        Din1 => VN1131_in1,
        Din2 => VN1131_in2,
        Din3 => VN1131_in3,
        Din4 => VN1131_in4,
        Din5 => VN1131_in5,
        VN2CN0_bit => VN_data_out(6786),
        VN2CN1_bit => VN_data_out(6787),
        VN2CN2_bit => VN_data_out(6788),
        VN2CN3_bit => VN_data_out(6789),
        VN2CN4_bit => VN_data_out(6790),
        VN2CN5_bit => VN_data_out(6791),
        VN2CN0_sign => VN_sign_out(6786),
        VN2CN1_sign => VN_sign_out(6787),
        VN2CN2_sign => VN_sign_out(6788),
        VN2CN3_sign => VN_sign_out(6789),
        VN2CN4_sign => VN_sign_out(6790),
        VN2CN5_sign => VN_sign_out(6791),
        codeword => codeword(1131),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1132 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6797 downto 6792),
        Din0 => VN1132_in0,
        Din1 => VN1132_in1,
        Din2 => VN1132_in2,
        Din3 => VN1132_in3,
        Din4 => VN1132_in4,
        Din5 => VN1132_in5,
        VN2CN0_bit => VN_data_out(6792),
        VN2CN1_bit => VN_data_out(6793),
        VN2CN2_bit => VN_data_out(6794),
        VN2CN3_bit => VN_data_out(6795),
        VN2CN4_bit => VN_data_out(6796),
        VN2CN5_bit => VN_data_out(6797),
        VN2CN0_sign => VN_sign_out(6792),
        VN2CN1_sign => VN_sign_out(6793),
        VN2CN2_sign => VN_sign_out(6794),
        VN2CN3_sign => VN_sign_out(6795),
        VN2CN4_sign => VN_sign_out(6796),
        VN2CN5_sign => VN_sign_out(6797),
        codeword => codeword(1132),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1133 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6803 downto 6798),
        Din0 => VN1133_in0,
        Din1 => VN1133_in1,
        Din2 => VN1133_in2,
        Din3 => VN1133_in3,
        Din4 => VN1133_in4,
        Din5 => VN1133_in5,
        VN2CN0_bit => VN_data_out(6798),
        VN2CN1_bit => VN_data_out(6799),
        VN2CN2_bit => VN_data_out(6800),
        VN2CN3_bit => VN_data_out(6801),
        VN2CN4_bit => VN_data_out(6802),
        VN2CN5_bit => VN_data_out(6803),
        VN2CN0_sign => VN_sign_out(6798),
        VN2CN1_sign => VN_sign_out(6799),
        VN2CN2_sign => VN_sign_out(6800),
        VN2CN3_sign => VN_sign_out(6801),
        VN2CN4_sign => VN_sign_out(6802),
        VN2CN5_sign => VN_sign_out(6803),
        codeword => codeword(1133),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1134 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6809 downto 6804),
        Din0 => VN1134_in0,
        Din1 => VN1134_in1,
        Din2 => VN1134_in2,
        Din3 => VN1134_in3,
        Din4 => VN1134_in4,
        Din5 => VN1134_in5,
        VN2CN0_bit => VN_data_out(6804),
        VN2CN1_bit => VN_data_out(6805),
        VN2CN2_bit => VN_data_out(6806),
        VN2CN3_bit => VN_data_out(6807),
        VN2CN4_bit => VN_data_out(6808),
        VN2CN5_bit => VN_data_out(6809),
        VN2CN0_sign => VN_sign_out(6804),
        VN2CN1_sign => VN_sign_out(6805),
        VN2CN2_sign => VN_sign_out(6806),
        VN2CN3_sign => VN_sign_out(6807),
        VN2CN4_sign => VN_sign_out(6808),
        VN2CN5_sign => VN_sign_out(6809),
        codeword => codeword(1134),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1135 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6815 downto 6810),
        Din0 => VN1135_in0,
        Din1 => VN1135_in1,
        Din2 => VN1135_in2,
        Din3 => VN1135_in3,
        Din4 => VN1135_in4,
        Din5 => VN1135_in5,
        VN2CN0_bit => VN_data_out(6810),
        VN2CN1_bit => VN_data_out(6811),
        VN2CN2_bit => VN_data_out(6812),
        VN2CN3_bit => VN_data_out(6813),
        VN2CN4_bit => VN_data_out(6814),
        VN2CN5_bit => VN_data_out(6815),
        VN2CN0_sign => VN_sign_out(6810),
        VN2CN1_sign => VN_sign_out(6811),
        VN2CN2_sign => VN_sign_out(6812),
        VN2CN3_sign => VN_sign_out(6813),
        VN2CN4_sign => VN_sign_out(6814),
        VN2CN5_sign => VN_sign_out(6815),
        codeword => codeword(1135),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1136 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6821 downto 6816),
        Din0 => VN1136_in0,
        Din1 => VN1136_in1,
        Din2 => VN1136_in2,
        Din3 => VN1136_in3,
        Din4 => VN1136_in4,
        Din5 => VN1136_in5,
        VN2CN0_bit => VN_data_out(6816),
        VN2CN1_bit => VN_data_out(6817),
        VN2CN2_bit => VN_data_out(6818),
        VN2CN3_bit => VN_data_out(6819),
        VN2CN4_bit => VN_data_out(6820),
        VN2CN5_bit => VN_data_out(6821),
        VN2CN0_sign => VN_sign_out(6816),
        VN2CN1_sign => VN_sign_out(6817),
        VN2CN2_sign => VN_sign_out(6818),
        VN2CN3_sign => VN_sign_out(6819),
        VN2CN4_sign => VN_sign_out(6820),
        VN2CN5_sign => VN_sign_out(6821),
        codeword => codeword(1136),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1137 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6827 downto 6822),
        Din0 => VN1137_in0,
        Din1 => VN1137_in1,
        Din2 => VN1137_in2,
        Din3 => VN1137_in3,
        Din4 => VN1137_in4,
        Din5 => VN1137_in5,
        VN2CN0_bit => VN_data_out(6822),
        VN2CN1_bit => VN_data_out(6823),
        VN2CN2_bit => VN_data_out(6824),
        VN2CN3_bit => VN_data_out(6825),
        VN2CN4_bit => VN_data_out(6826),
        VN2CN5_bit => VN_data_out(6827),
        VN2CN0_sign => VN_sign_out(6822),
        VN2CN1_sign => VN_sign_out(6823),
        VN2CN2_sign => VN_sign_out(6824),
        VN2CN3_sign => VN_sign_out(6825),
        VN2CN4_sign => VN_sign_out(6826),
        VN2CN5_sign => VN_sign_out(6827),
        codeword => codeword(1137),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1138 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6833 downto 6828),
        Din0 => VN1138_in0,
        Din1 => VN1138_in1,
        Din2 => VN1138_in2,
        Din3 => VN1138_in3,
        Din4 => VN1138_in4,
        Din5 => VN1138_in5,
        VN2CN0_bit => VN_data_out(6828),
        VN2CN1_bit => VN_data_out(6829),
        VN2CN2_bit => VN_data_out(6830),
        VN2CN3_bit => VN_data_out(6831),
        VN2CN4_bit => VN_data_out(6832),
        VN2CN5_bit => VN_data_out(6833),
        VN2CN0_sign => VN_sign_out(6828),
        VN2CN1_sign => VN_sign_out(6829),
        VN2CN2_sign => VN_sign_out(6830),
        VN2CN3_sign => VN_sign_out(6831),
        VN2CN4_sign => VN_sign_out(6832),
        VN2CN5_sign => VN_sign_out(6833),
        codeword => codeword(1138),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1139 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6839 downto 6834),
        Din0 => VN1139_in0,
        Din1 => VN1139_in1,
        Din2 => VN1139_in2,
        Din3 => VN1139_in3,
        Din4 => VN1139_in4,
        Din5 => VN1139_in5,
        VN2CN0_bit => VN_data_out(6834),
        VN2CN1_bit => VN_data_out(6835),
        VN2CN2_bit => VN_data_out(6836),
        VN2CN3_bit => VN_data_out(6837),
        VN2CN4_bit => VN_data_out(6838),
        VN2CN5_bit => VN_data_out(6839),
        VN2CN0_sign => VN_sign_out(6834),
        VN2CN1_sign => VN_sign_out(6835),
        VN2CN2_sign => VN_sign_out(6836),
        VN2CN3_sign => VN_sign_out(6837),
        VN2CN4_sign => VN_sign_out(6838),
        VN2CN5_sign => VN_sign_out(6839),
        codeword => codeword(1139),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1140 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6845 downto 6840),
        Din0 => VN1140_in0,
        Din1 => VN1140_in1,
        Din2 => VN1140_in2,
        Din3 => VN1140_in3,
        Din4 => VN1140_in4,
        Din5 => VN1140_in5,
        VN2CN0_bit => VN_data_out(6840),
        VN2CN1_bit => VN_data_out(6841),
        VN2CN2_bit => VN_data_out(6842),
        VN2CN3_bit => VN_data_out(6843),
        VN2CN4_bit => VN_data_out(6844),
        VN2CN5_bit => VN_data_out(6845),
        VN2CN0_sign => VN_sign_out(6840),
        VN2CN1_sign => VN_sign_out(6841),
        VN2CN2_sign => VN_sign_out(6842),
        VN2CN3_sign => VN_sign_out(6843),
        VN2CN4_sign => VN_sign_out(6844),
        VN2CN5_sign => VN_sign_out(6845),
        codeword => codeword(1140),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1141 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6851 downto 6846),
        Din0 => VN1141_in0,
        Din1 => VN1141_in1,
        Din2 => VN1141_in2,
        Din3 => VN1141_in3,
        Din4 => VN1141_in4,
        Din5 => VN1141_in5,
        VN2CN0_bit => VN_data_out(6846),
        VN2CN1_bit => VN_data_out(6847),
        VN2CN2_bit => VN_data_out(6848),
        VN2CN3_bit => VN_data_out(6849),
        VN2CN4_bit => VN_data_out(6850),
        VN2CN5_bit => VN_data_out(6851),
        VN2CN0_sign => VN_sign_out(6846),
        VN2CN1_sign => VN_sign_out(6847),
        VN2CN2_sign => VN_sign_out(6848),
        VN2CN3_sign => VN_sign_out(6849),
        VN2CN4_sign => VN_sign_out(6850),
        VN2CN5_sign => VN_sign_out(6851),
        codeword => codeword(1141),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1142 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6857 downto 6852),
        Din0 => VN1142_in0,
        Din1 => VN1142_in1,
        Din2 => VN1142_in2,
        Din3 => VN1142_in3,
        Din4 => VN1142_in4,
        Din5 => VN1142_in5,
        VN2CN0_bit => VN_data_out(6852),
        VN2CN1_bit => VN_data_out(6853),
        VN2CN2_bit => VN_data_out(6854),
        VN2CN3_bit => VN_data_out(6855),
        VN2CN4_bit => VN_data_out(6856),
        VN2CN5_bit => VN_data_out(6857),
        VN2CN0_sign => VN_sign_out(6852),
        VN2CN1_sign => VN_sign_out(6853),
        VN2CN2_sign => VN_sign_out(6854),
        VN2CN3_sign => VN_sign_out(6855),
        VN2CN4_sign => VN_sign_out(6856),
        VN2CN5_sign => VN_sign_out(6857),
        codeword => codeword(1142),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1143 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6863 downto 6858),
        Din0 => VN1143_in0,
        Din1 => VN1143_in1,
        Din2 => VN1143_in2,
        Din3 => VN1143_in3,
        Din4 => VN1143_in4,
        Din5 => VN1143_in5,
        VN2CN0_bit => VN_data_out(6858),
        VN2CN1_bit => VN_data_out(6859),
        VN2CN2_bit => VN_data_out(6860),
        VN2CN3_bit => VN_data_out(6861),
        VN2CN4_bit => VN_data_out(6862),
        VN2CN5_bit => VN_data_out(6863),
        VN2CN0_sign => VN_sign_out(6858),
        VN2CN1_sign => VN_sign_out(6859),
        VN2CN2_sign => VN_sign_out(6860),
        VN2CN3_sign => VN_sign_out(6861),
        VN2CN4_sign => VN_sign_out(6862),
        VN2CN5_sign => VN_sign_out(6863),
        codeword => codeword(1143),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1144 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6869 downto 6864),
        Din0 => VN1144_in0,
        Din1 => VN1144_in1,
        Din2 => VN1144_in2,
        Din3 => VN1144_in3,
        Din4 => VN1144_in4,
        Din5 => VN1144_in5,
        VN2CN0_bit => VN_data_out(6864),
        VN2CN1_bit => VN_data_out(6865),
        VN2CN2_bit => VN_data_out(6866),
        VN2CN3_bit => VN_data_out(6867),
        VN2CN4_bit => VN_data_out(6868),
        VN2CN5_bit => VN_data_out(6869),
        VN2CN0_sign => VN_sign_out(6864),
        VN2CN1_sign => VN_sign_out(6865),
        VN2CN2_sign => VN_sign_out(6866),
        VN2CN3_sign => VN_sign_out(6867),
        VN2CN4_sign => VN_sign_out(6868),
        VN2CN5_sign => VN_sign_out(6869),
        codeword => codeword(1144),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1145 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6875 downto 6870),
        Din0 => VN1145_in0,
        Din1 => VN1145_in1,
        Din2 => VN1145_in2,
        Din3 => VN1145_in3,
        Din4 => VN1145_in4,
        Din5 => VN1145_in5,
        VN2CN0_bit => VN_data_out(6870),
        VN2CN1_bit => VN_data_out(6871),
        VN2CN2_bit => VN_data_out(6872),
        VN2CN3_bit => VN_data_out(6873),
        VN2CN4_bit => VN_data_out(6874),
        VN2CN5_bit => VN_data_out(6875),
        VN2CN0_sign => VN_sign_out(6870),
        VN2CN1_sign => VN_sign_out(6871),
        VN2CN2_sign => VN_sign_out(6872),
        VN2CN3_sign => VN_sign_out(6873),
        VN2CN4_sign => VN_sign_out(6874),
        VN2CN5_sign => VN_sign_out(6875),
        codeword => codeword(1145),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1146 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6881 downto 6876),
        Din0 => VN1146_in0,
        Din1 => VN1146_in1,
        Din2 => VN1146_in2,
        Din3 => VN1146_in3,
        Din4 => VN1146_in4,
        Din5 => VN1146_in5,
        VN2CN0_bit => VN_data_out(6876),
        VN2CN1_bit => VN_data_out(6877),
        VN2CN2_bit => VN_data_out(6878),
        VN2CN3_bit => VN_data_out(6879),
        VN2CN4_bit => VN_data_out(6880),
        VN2CN5_bit => VN_data_out(6881),
        VN2CN0_sign => VN_sign_out(6876),
        VN2CN1_sign => VN_sign_out(6877),
        VN2CN2_sign => VN_sign_out(6878),
        VN2CN3_sign => VN_sign_out(6879),
        VN2CN4_sign => VN_sign_out(6880),
        VN2CN5_sign => VN_sign_out(6881),
        codeword => codeword(1146),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1147 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6887 downto 6882),
        Din0 => VN1147_in0,
        Din1 => VN1147_in1,
        Din2 => VN1147_in2,
        Din3 => VN1147_in3,
        Din4 => VN1147_in4,
        Din5 => VN1147_in5,
        VN2CN0_bit => VN_data_out(6882),
        VN2CN1_bit => VN_data_out(6883),
        VN2CN2_bit => VN_data_out(6884),
        VN2CN3_bit => VN_data_out(6885),
        VN2CN4_bit => VN_data_out(6886),
        VN2CN5_bit => VN_data_out(6887),
        VN2CN0_sign => VN_sign_out(6882),
        VN2CN1_sign => VN_sign_out(6883),
        VN2CN2_sign => VN_sign_out(6884),
        VN2CN3_sign => VN_sign_out(6885),
        VN2CN4_sign => VN_sign_out(6886),
        VN2CN5_sign => VN_sign_out(6887),
        codeword => codeword(1147),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1148 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6893 downto 6888),
        Din0 => VN1148_in0,
        Din1 => VN1148_in1,
        Din2 => VN1148_in2,
        Din3 => VN1148_in3,
        Din4 => VN1148_in4,
        Din5 => VN1148_in5,
        VN2CN0_bit => VN_data_out(6888),
        VN2CN1_bit => VN_data_out(6889),
        VN2CN2_bit => VN_data_out(6890),
        VN2CN3_bit => VN_data_out(6891),
        VN2CN4_bit => VN_data_out(6892),
        VN2CN5_bit => VN_data_out(6893),
        VN2CN0_sign => VN_sign_out(6888),
        VN2CN1_sign => VN_sign_out(6889),
        VN2CN2_sign => VN_sign_out(6890),
        VN2CN3_sign => VN_sign_out(6891),
        VN2CN4_sign => VN_sign_out(6892),
        VN2CN5_sign => VN_sign_out(6893),
        codeword => codeword(1148),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1149 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6899 downto 6894),
        Din0 => VN1149_in0,
        Din1 => VN1149_in1,
        Din2 => VN1149_in2,
        Din3 => VN1149_in3,
        Din4 => VN1149_in4,
        Din5 => VN1149_in5,
        VN2CN0_bit => VN_data_out(6894),
        VN2CN1_bit => VN_data_out(6895),
        VN2CN2_bit => VN_data_out(6896),
        VN2CN3_bit => VN_data_out(6897),
        VN2CN4_bit => VN_data_out(6898),
        VN2CN5_bit => VN_data_out(6899),
        VN2CN0_sign => VN_sign_out(6894),
        VN2CN1_sign => VN_sign_out(6895),
        VN2CN2_sign => VN_sign_out(6896),
        VN2CN3_sign => VN_sign_out(6897),
        VN2CN4_sign => VN_sign_out(6898),
        VN2CN5_sign => VN_sign_out(6899),
        codeword => codeword(1149),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1150 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6905 downto 6900),
        Din0 => VN1150_in0,
        Din1 => VN1150_in1,
        Din2 => VN1150_in2,
        Din3 => VN1150_in3,
        Din4 => VN1150_in4,
        Din5 => VN1150_in5,
        VN2CN0_bit => VN_data_out(6900),
        VN2CN1_bit => VN_data_out(6901),
        VN2CN2_bit => VN_data_out(6902),
        VN2CN3_bit => VN_data_out(6903),
        VN2CN4_bit => VN_data_out(6904),
        VN2CN5_bit => VN_data_out(6905),
        VN2CN0_sign => VN_sign_out(6900),
        VN2CN1_sign => VN_sign_out(6901),
        VN2CN2_sign => VN_sign_out(6902),
        VN2CN3_sign => VN_sign_out(6903),
        VN2CN4_sign => VN_sign_out(6904),
        VN2CN5_sign => VN_sign_out(6905),
        codeword => codeword(1150),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1151 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6911 downto 6906),
        Din0 => VN1151_in0,
        Din1 => VN1151_in1,
        Din2 => VN1151_in2,
        Din3 => VN1151_in3,
        Din4 => VN1151_in4,
        Din5 => VN1151_in5,
        VN2CN0_bit => VN_data_out(6906),
        VN2CN1_bit => VN_data_out(6907),
        VN2CN2_bit => VN_data_out(6908),
        VN2CN3_bit => VN_data_out(6909),
        VN2CN4_bit => VN_data_out(6910),
        VN2CN5_bit => VN_data_out(6911),
        VN2CN0_sign => VN_sign_out(6906),
        VN2CN1_sign => VN_sign_out(6907),
        VN2CN2_sign => VN_sign_out(6908),
        VN2CN3_sign => VN_sign_out(6909),
        VN2CN4_sign => VN_sign_out(6910),
        VN2CN5_sign => VN_sign_out(6911),
        codeword => codeword(1151),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1152 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6917 downto 6912),
        Din0 => VN1152_in0,
        Din1 => VN1152_in1,
        Din2 => VN1152_in2,
        Din3 => VN1152_in3,
        Din4 => VN1152_in4,
        Din5 => VN1152_in5,
        VN2CN0_bit => VN_data_out(6912),
        VN2CN1_bit => VN_data_out(6913),
        VN2CN2_bit => VN_data_out(6914),
        VN2CN3_bit => VN_data_out(6915),
        VN2CN4_bit => VN_data_out(6916),
        VN2CN5_bit => VN_data_out(6917),
        VN2CN0_sign => VN_sign_out(6912),
        VN2CN1_sign => VN_sign_out(6913),
        VN2CN2_sign => VN_sign_out(6914),
        VN2CN3_sign => VN_sign_out(6915),
        VN2CN4_sign => VN_sign_out(6916),
        VN2CN5_sign => VN_sign_out(6917),
        codeword => codeword(1152),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1153 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6923 downto 6918),
        Din0 => VN1153_in0,
        Din1 => VN1153_in1,
        Din2 => VN1153_in2,
        Din3 => VN1153_in3,
        Din4 => VN1153_in4,
        Din5 => VN1153_in5,
        VN2CN0_bit => VN_data_out(6918),
        VN2CN1_bit => VN_data_out(6919),
        VN2CN2_bit => VN_data_out(6920),
        VN2CN3_bit => VN_data_out(6921),
        VN2CN4_bit => VN_data_out(6922),
        VN2CN5_bit => VN_data_out(6923),
        VN2CN0_sign => VN_sign_out(6918),
        VN2CN1_sign => VN_sign_out(6919),
        VN2CN2_sign => VN_sign_out(6920),
        VN2CN3_sign => VN_sign_out(6921),
        VN2CN4_sign => VN_sign_out(6922),
        VN2CN5_sign => VN_sign_out(6923),
        codeword => codeword(1153),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1154 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6929 downto 6924),
        Din0 => VN1154_in0,
        Din1 => VN1154_in1,
        Din2 => VN1154_in2,
        Din3 => VN1154_in3,
        Din4 => VN1154_in4,
        Din5 => VN1154_in5,
        VN2CN0_bit => VN_data_out(6924),
        VN2CN1_bit => VN_data_out(6925),
        VN2CN2_bit => VN_data_out(6926),
        VN2CN3_bit => VN_data_out(6927),
        VN2CN4_bit => VN_data_out(6928),
        VN2CN5_bit => VN_data_out(6929),
        VN2CN0_sign => VN_sign_out(6924),
        VN2CN1_sign => VN_sign_out(6925),
        VN2CN2_sign => VN_sign_out(6926),
        VN2CN3_sign => VN_sign_out(6927),
        VN2CN4_sign => VN_sign_out(6928),
        VN2CN5_sign => VN_sign_out(6929),
        codeword => codeword(1154),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1155 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6935 downto 6930),
        Din0 => VN1155_in0,
        Din1 => VN1155_in1,
        Din2 => VN1155_in2,
        Din3 => VN1155_in3,
        Din4 => VN1155_in4,
        Din5 => VN1155_in5,
        VN2CN0_bit => VN_data_out(6930),
        VN2CN1_bit => VN_data_out(6931),
        VN2CN2_bit => VN_data_out(6932),
        VN2CN3_bit => VN_data_out(6933),
        VN2CN4_bit => VN_data_out(6934),
        VN2CN5_bit => VN_data_out(6935),
        VN2CN0_sign => VN_sign_out(6930),
        VN2CN1_sign => VN_sign_out(6931),
        VN2CN2_sign => VN_sign_out(6932),
        VN2CN3_sign => VN_sign_out(6933),
        VN2CN4_sign => VN_sign_out(6934),
        VN2CN5_sign => VN_sign_out(6935),
        codeword => codeword(1155),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1156 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6941 downto 6936),
        Din0 => VN1156_in0,
        Din1 => VN1156_in1,
        Din2 => VN1156_in2,
        Din3 => VN1156_in3,
        Din4 => VN1156_in4,
        Din5 => VN1156_in5,
        VN2CN0_bit => VN_data_out(6936),
        VN2CN1_bit => VN_data_out(6937),
        VN2CN2_bit => VN_data_out(6938),
        VN2CN3_bit => VN_data_out(6939),
        VN2CN4_bit => VN_data_out(6940),
        VN2CN5_bit => VN_data_out(6941),
        VN2CN0_sign => VN_sign_out(6936),
        VN2CN1_sign => VN_sign_out(6937),
        VN2CN2_sign => VN_sign_out(6938),
        VN2CN3_sign => VN_sign_out(6939),
        VN2CN4_sign => VN_sign_out(6940),
        VN2CN5_sign => VN_sign_out(6941),
        codeword => codeword(1156),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1157 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6947 downto 6942),
        Din0 => VN1157_in0,
        Din1 => VN1157_in1,
        Din2 => VN1157_in2,
        Din3 => VN1157_in3,
        Din4 => VN1157_in4,
        Din5 => VN1157_in5,
        VN2CN0_bit => VN_data_out(6942),
        VN2CN1_bit => VN_data_out(6943),
        VN2CN2_bit => VN_data_out(6944),
        VN2CN3_bit => VN_data_out(6945),
        VN2CN4_bit => VN_data_out(6946),
        VN2CN5_bit => VN_data_out(6947),
        VN2CN0_sign => VN_sign_out(6942),
        VN2CN1_sign => VN_sign_out(6943),
        VN2CN2_sign => VN_sign_out(6944),
        VN2CN3_sign => VN_sign_out(6945),
        VN2CN4_sign => VN_sign_out(6946),
        VN2CN5_sign => VN_sign_out(6947),
        codeword => codeword(1157),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1158 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6953 downto 6948),
        Din0 => VN1158_in0,
        Din1 => VN1158_in1,
        Din2 => VN1158_in2,
        Din3 => VN1158_in3,
        Din4 => VN1158_in4,
        Din5 => VN1158_in5,
        VN2CN0_bit => VN_data_out(6948),
        VN2CN1_bit => VN_data_out(6949),
        VN2CN2_bit => VN_data_out(6950),
        VN2CN3_bit => VN_data_out(6951),
        VN2CN4_bit => VN_data_out(6952),
        VN2CN5_bit => VN_data_out(6953),
        VN2CN0_sign => VN_sign_out(6948),
        VN2CN1_sign => VN_sign_out(6949),
        VN2CN2_sign => VN_sign_out(6950),
        VN2CN3_sign => VN_sign_out(6951),
        VN2CN4_sign => VN_sign_out(6952),
        VN2CN5_sign => VN_sign_out(6953),
        codeword => codeword(1158),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1159 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6959 downto 6954),
        Din0 => VN1159_in0,
        Din1 => VN1159_in1,
        Din2 => VN1159_in2,
        Din3 => VN1159_in3,
        Din4 => VN1159_in4,
        Din5 => VN1159_in5,
        VN2CN0_bit => VN_data_out(6954),
        VN2CN1_bit => VN_data_out(6955),
        VN2CN2_bit => VN_data_out(6956),
        VN2CN3_bit => VN_data_out(6957),
        VN2CN4_bit => VN_data_out(6958),
        VN2CN5_bit => VN_data_out(6959),
        VN2CN0_sign => VN_sign_out(6954),
        VN2CN1_sign => VN_sign_out(6955),
        VN2CN2_sign => VN_sign_out(6956),
        VN2CN3_sign => VN_sign_out(6957),
        VN2CN4_sign => VN_sign_out(6958),
        VN2CN5_sign => VN_sign_out(6959),
        codeword => codeword(1159),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1160 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6965 downto 6960),
        Din0 => VN1160_in0,
        Din1 => VN1160_in1,
        Din2 => VN1160_in2,
        Din3 => VN1160_in3,
        Din4 => VN1160_in4,
        Din5 => VN1160_in5,
        VN2CN0_bit => VN_data_out(6960),
        VN2CN1_bit => VN_data_out(6961),
        VN2CN2_bit => VN_data_out(6962),
        VN2CN3_bit => VN_data_out(6963),
        VN2CN4_bit => VN_data_out(6964),
        VN2CN5_bit => VN_data_out(6965),
        VN2CN0_sign => VN_sign_out(6960),
        VN2CN1_sign => VN_sign_out(6961),
        VN2CN2_sign => VN_sign_out(6962),
        VN2CN3_sign => VN_sign_out(6963),
        VN2CN4_sign => VN_sign_out(6964),
        VN2CN5_sign => VN_sign_out(6965),
        codeword => codeword(1160),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1161 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6971 downto 6966),
        Din0 => VN1161_in0,
        Din1 => VN1161_in1,
        Din2 => VN1161_in2,
        Din3 => VN1161_in3,
        Din4 => VN1161_in4,
        Din5 => VN1161_in5,
        VN2CN0_bit => VN_data_out(6966),
        VN2CN1_bit => VN_data_out(6967),
        VN2CN2_bit => VN_data_out(6968),
        VN2CN3_bit => VN_data_out(6969),
        VN2CN4_bit => VN_data_out(6970),
        VN2CN5_bit => VN_data_out(6971),
        VN2CN0_sign => VN_sign_out(6966),
        VN2CN1_sign => VN_sign_out(6967),
        VN2CN2_sign => VN_sign_out(6968),
        VN2CN3_sign => VN_sign_out(6969),
        VN2CN4_sign => VN_sign_out(6970),
        VN2CN5_sign => VN_sign_out(6971),
        codeword => codeword(1161),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1162 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6977 downto 6972),
        Din0 => VN1162_in0,
        Din1 => VN1162_in1,
        Din2 => VN1162_in2,
        Din3 => VN1162_in3,
        Din4 => VN1162_in4,
        Din5 => VN1162_in5,
        VN2CN0_bit => VN_data_out(6972),
        VN2CN1_bit => VN_data_out(6973),
        VN2CN2_bit => VN_data_out(6974),
        VN2CN3_bit => VN_data_out(6975),
        VN2CN4_bit => VN_data_out(6976),
        VN2CN5_bit => VN_data_out(6977),
        VN2CN0_sign => VN_sign_out(6972),
        VN2CN1_sign => VN_sign_out(6973),
        VN2CN2_sign => VN_sign_out(6974),
        VN2CN3_sign => VN_sign_out(6975),
        VN2CN4_sign => VN_sign_out(6976),
        VN2CN5_sign => VN_sign_out(6977),
        codeword => codeword(1162),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1163 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6983 downto 6978),
        Din0 => VN1163_in0,
        Din1 => VN1163_in1,
        Din2 => VN1163_in2,
        Din3 => VN1163_in3,
        Din4 => VN1163_in4,
        Din5 => VN1163_in5,
        VN2CN0_bit => VN_data_out(6978),
        VN2CN1_bit => VN_data_out(6979),
        VN2CN2_bit => VN_data_out(6980),
        VN2CN3_bit => VN_data_out(6981),
        VN2CN4_bit => VN_data_out(6982),
        VN2CN5_bit => VN_data_out(6983),
        VN2CN0_sign => VN_sign_out(6978),
        VN2CN1_sign => VN_sign_out(6979),
        VN2CN2_sign => VN_sign_out(6980),
        VN2CN3_sign => VN_sign_out(6981),
        VN2CN4_sign => VN_sign_out(6982),
        VN2CN5_sign => VN_sign_out(6983),
        codeword => codeword(1163),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1164 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6989 downto 6984),
        Din0 => VN1164_in0,
        Din1 => VN1164_in1,
        Din2 => VN1164_in2,
        Din3 => VN1164_in3,
        Din4 => VN1164_in4,
        Din5 => VN1164_in5,
        VN2CN0_bit => VN_data_out(6984),
        VN2CN1_bit => VN_data_out(6985),
        VN2CN2_bit => VN_data_out(6986),
        VN2CN3_bit => VN_data_out(6987),
        VN2CN4_bit => VN_data_out(6988),
        VN2CN5_bit => VN_data_out(6989),
        VN2CN0_sign => VN_sign_out(6984),
        VN2CN1_sign => VN_sign_out(6985),
        VN2CN2_sign => VN_sign_out(6986),
        VN2CN3_sign => VN_sign_out(6987),
        VN2CN4_sign => VN_sign_out(6988),
        VN2CN5_sign => VN_sign_out(6989),
        codeword => codeword(1164),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1165 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(6995 downto 6990),
        Din0 => VN1165_in0,
        Din1 => VN1165_in1,
        Din2 => VN1165_in2,
        Din3 => VN1165_in3,
        Din4 => VN1165_in4,
        Din5 => VN1165_in5,
        VN2CN0_bit => VN_data_out(6990),
        VN2CN1_bit => VN_data_out(6991),
        VN2CN2_bit => VN_data_out(6992),
        VN2CN3_bit => VN_data_out(6993),
        VN2CN4_bit => VN_data_out(6994),
        VN2CN5_bit => VN_data_out(6995),
        VN2CN0_sign => VN_sign_out(6990),
        VN2CN1_sign => VN_sign_out(6991),
        VN2CN2_sign => VN_sign_out(6992),
        VN2CN3_sign => VN_sign_out(6993),
        VN2CN4_sign => VN_sign_out(6994),
        VN2CN5_sign => VN_sign_out(6995),
        codeword => codeword(1165),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1166 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7001 downto 6996),
        Din0 => VN1166_in0,
        Din1 => VN1166_in1,
        Din2 => VN1166_in2,
        Din3 => VN1166_in3,
        Din4 => VN1166_in4,
        Din5 => VN1166_in5,
        VN2CN0_bit => VN_data_out(6996),
        VN2CN1_bit => VN_data_out(6997),
        VN2CN2_bit => VN_data_out(6998),
        VN2CN3_bit => VN_data_out(6999),
        VN2CN4_bit => VN_data_out(7000),
        VN2CN5_bit => VN_data_out(7001),
        VN2CN0_sign => VN_sign_out(6996),
        VN2CN1_sign => VN_sign_out(6997),
        VN2CN2_sign => VN_sign_out(6998),
        VN2CN3_sign => VN_sign_out(6999),
        VN2CN4_sign => VN_sign_out(7000),
        VN2CN5_sign => VN_sign_out(7001),
        codeword => codeword(1166),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1167 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7007 downto 7002),
        Din0 => VN1167_in0,
        Din1 => VN1167_in1,
        Din2 => VN1167_in2,
        Din3 => VN1167_in3,
        Din4 => VN1167_in4,
        Din5 => VN1167_in5,
        VN2CN0_bit => VN_data_out(7002),
        VN2CN1_bit => VN_data_out(7003),
        VN2CN2_bit => VN_data_out(7004),
        VN2CN3_bit => VN_data_out(7005),
        VN2CN4_bit => VN_data_out(7006),
        VN2CN5_bit => VN_data_out(7007),
        VN2CN0_sign => VN_sign_out(7002),
        VN2CN1_sign => VN_sign_out(7003),
        VN2CN2_sign => VN_sign_out(7004),
        VN2CN3_sign => VN_sign_out(7005),
        VN2CN4_sign => VN_sign_out(7006),
        VN2CN5_sign => VN_sign_out(7007),
        codeword => codeword(1167),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1168 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7013 downto 7008),
        Din0 => VN1168_in0,
        Din1 => VN1168_in1,
        Din2 => VN1168_in2,
        Din3 => VN1168_in3,
        Din4 => VN1168_in4,
        Din5 => VN1168_in5,
        VN2CN0_bit => VN_data_out(7008),
        VN2CN1_bit => VN_data_out(7009),
        VN2CN2_bit => VN_data_out(7010),
        VN2CN3_bit => VN_data_out(7011),
        VN2CN4_bit => VN_data_out(7012),
        VN2CN5_bit => VN_data_out(7013),
        VN2CN0_sign => VN_sign_out(7008),
        VN2CN1_sign => VN_sign_out(7009),
        VN2CN2_sign => VN_sign_out(7010),
        VN2CN3_sign => VN_sign_out(7011),
        VN2CN4_sign => VN_sign_out(7012),
        VN2CN5_sign => VN_sign_out(7013),
        codeword => codeword(1168),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1169 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7019 downto 7014),
        Din0 => VN1169_in0,
        Din1 => VN1169_in1,
        Din2 => VN1169_in2,
        Din3 => VN1169_in3,
        Din4 => VN1169_in4,
        Din5 => VN1169_in5,
        VN2CN0_bit => VN_data_out(7014),
        VN2CN1_bit => VN_data_out(7015),
        VN2CN2_bit => VN_data_out(7016),
        VN2CN3_bit => VN_data_out(7017),
        VN2CN4_bit => VN_data_out(7018),
        VN2CN5_bit => VN_data_out(7019),
        VN2CN0_sign => VN_sign_out(7014),
        VN2CN1_sign => VN_sign_out(7015),
        VN2CN2_sign => VN_sign_out(7016),
        VN2CN3_sign => VN_sign_out(7017),
        VN2CN4_sign => VN_sign_out(7018),
        VN2CN5_sign => VN_sign_out(7019),
        codeword => codeword(1169),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1170 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7025 downto 7020),
        Din0 => VN1170_in0,
        Din1 => VN1170_in1,
        Din2 => VN1170_in2,
        Din3 => VN1170_in3,
        Din4 => VN1170_in4,
        Din5 => VN1170_in5,
        VN2CN0_bit => VN_data_out(7020),
        VN2CN1_bit => VN_data_out(7021),
        VN2CN2_bit => VN_data_out(7022),
        VN2CN3_bit => VN_data_out(7023),
        VN2CN4_bit => VN_data_out(7024),
        VN2CN5_bit => VN_data_out(7025),
        VN2CN0_sign => VN_sign_out(7020),
        VN2CN1_sign => VN_sign_out(7021),
        VN2CN2_sign => VN_sign_out(7022),
        VN2CN3_sign => VN_sign_out(7023),
        VN2CN4_sign => VN_sign_out(7024),
        VN2CN5_sign => VN_sign_out(7025),
        codeword => codeword(1170),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1171 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7031 downto 7026),
        Din0 => VN1171_in0,
        Din1 => VN1171_in1,
        Din2 => VN1171_in2,
        Din3 => VN1171_in3,
        Din4 => VN1171_in4,
        Din5 => VN1171_in5,
        VN2CN0_bit => VN_data_out(7026),
        VN2CN1_bit => VN_data_out(7027),
        VN2CN2_bit => VN_data_out(7028),
        VN2CN3_bit => VN_data_out(7029),
        VN2CN4_bit => VN_data_out(7030),
        VN2CN5_bit => VN_data_out(7031),
        VN2CN0_sign => VN_sign_out(7026),
        VN2CN1_sign => VN_sign_out(7027),
        VN2CN2_sign => VN_sign_out(7028),
        VN2CN3_sign => VN_sign_out(7029),
        VN2CN4_sign => VN_sign_out(7030),
        VN2CN5_sign => VN_sign_out(7031),
        codeword => codeword(1171),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1172 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7037 downto 7032),
        Din0 => VN1172_in0,
        Din1 => VN1172_in1,
        Din2 => VN1172_in2,
        Din3 => VN1172_in3,
        Din4 => VN1172_in4,
        Din5 => VN1172_in5,
        VN2CN0_bit => VN_data_out(7032),
        VN2CN1_bit => VN_data_out(7033),
        VN2CN2_bit => VN_data_out(7034),
        VN2CN3_bit => VN_data_out(7035),
        VN2CN4_bit => VN_data_out(7036),
        VN2CN5_bit => VN_data_out(7037),
        VN2CN0_sign => VN_sign_out(7032),
        VN2CN1_sign => VN_sign_out(7033),
        VN2CN2_sign => VN_sign_out(7034),
        VN2CN3_sign => VN_sign_out(7035),
        VN2CN4_sign => VN_sign_out(7036),
        VN2CN5_sign => VN_sign_out(7037),
        codeword => codeword(1172),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1173 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7043 downto 7038),
        Din0 => VN1173_in0,
        Din1 => VN1173_in1,
        Din2 => VN1173_in2,
        Din3 => VN1173_in3,
        Din4 => VN1173_in4,
        Din5 => VN1173_in5,
        VN2CN0_bit => VN_data_out(7038),
        VN2CN1_bit => VN_data_out(7039),
        VN2CN2_bit => VN_data_out(7040),
        VN2CN3_bit => VN_data_out(7041),
        VN2CN4_bit => VN_data_out(7042),
        VN2CN5_bit => VN_data_out(7043),
        VN2CN0_sign => VN_sign_out(7038),
        VN2CN1_sign => VN_sign_out(7039),
        VN2CN2_sign => VN_sign_out(7040),
        VN2CN3_sign => VN_sign_out(7041),
        VN2CN4_sign => VN_sign_out(7042),
        VN2CN5_sign => VN_sign_out(7043),
        codeword => codeword(1173),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1174 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7049 downto 7044),
        Din0 => VN1174_in0,
        Din1 => VN1174_in1,
        Din2 => VN1174_in2,
        Din3 => VN1174_in3,
        Din4 => VN1174_in4,
        Din5 => VN1174_in5,
        VN2CN0_bit => VN_data_out(7044),
        VN2CN1_bit => VN_data_out(7045),
        VN2CN2_bit => VN_data_out(7046),
        VN2CN3_bit => VN_data_out(7047),
        VN2CN4_bit => VN_data_out(7048),
        VN2CN5_bit => VN_data_out(7049),
        VN2CN0_sign => VN_sign_out(7044),
        VN2CN1_sign => VN_sign_out(7045),
        VN2CN2_sign => VN_sign_out(7046),
        VN2CN3_sign => VN_sign_out(7047),
        VN2CN4_sign => VN_sign_out(7048),
        VN2CN5_sign => VN_sign_out(7049),
        codeword => codeword(1174),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1175 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7055 downto 7050),
        Din0 => VN1175_in0,
        Din1 => VN1175_in1,
        Din2 => VN1175_in2,
        Din3 => VN1175_in3,
        Din4 => VN1175_in4,
        Din5 => VN1175_in5,
        VN2CN0_bit => VN_data_out(7050),
        VN2CN1_bit => VN_data_out(7051),
        VN2CN2_bit => VN_data_out(7052),
        VN2CN3_bit => VN_data_out(7053),
        VN2CN4_bit => VN_data_out(7054),
        VN2CN5_bit => VN_data_out(7055),
        VN2CN0_sign => VN_sign_out(7050),
        VN2CN1_sign => VN_sign_out(7051),
        VN2CN2_sign => VN_sign_out(7052),
        VN2CN3_sign => VN_sign_out(7053),
        VN2CN4_sign => VN_sign_out(7054),
        VN2CN5_sign => VN_sign_out(7055),
        codeword => codeword(1175),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1176 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7061 downto 7056),
        Din0 => VN1176_in0,
        Din1 => VN1176_in1,
        Din2 => VN1176_in2,
        Din3 => VN1176_in3,
        Din4 => VN1176_in4,
        Din5 => VN1176_in5,
        VN2CN0_bit => VN_data_out(7056),
        VN2CN1_bit => VN_data_out(7057),
        VN2CN2_bit => VN_data_out(7058),
        VN2CN3_bit => VN_data_out(7059),
        VN2CN4_bit => VN_data_out(7060),
        VN2CN5_bit => VN_data_out(7061),
        VN2CN0_sign => VN_sign_out(7056),
        VN2CN1_sign => VN_sign_out(7057),
        VN2CN2_sign => VN_sign_out(7058),
        VN2CN3_sign => VN_sign_out(7059),
        VN2CN4_sign => VN_sign_out(7060),
        VN2CN5_sign => VN_sign_out(7061),
        codeword => codeword(1176),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1177 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7067 downto 7062),
        Din0 => VN1177_in0,
        Din1 => VN1177_in1,
        Din2 => VN1177_in2,
        Din3 => VN1177_in3,
        Din4 => VN1177_in4,
        Din5 => VN1177_in5,
        VN2CN0_bit => VN_data_out(7062),
        VN2CN1_bit => VN_data_out(7063),
        VN2CN2_bit => VN_data_out(7064),
        VN2CN3_bit => VN_data_out(7065),
        VN2CN4_bit => VN_data_out(7066),
        VN2CN5_bit => VN_data_out(7067),
        VN2CN0_sign => VN_sign_out(7062),
        VN2CN1_sign => VN_sign_out(7063),
        VN2CN2_sign => VN_sign_out(7064),
        VN2CN3_sign => VN_sign_out(7065),
        VN2CN4_sign => VN_sign_out(7066),
        VN2CN5_sign => VN_sign_out(7067),
        codeword => codeword(1177),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1178 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7073 downto 7068),
        Din0 => VN1178_in0,
        Din1 => VN1178_in1,
        Din2 => VN1178_in2,
        Din3 => VN1178_in3,
        Din4 => VN1178_in4,
        Din5 => VN1178_in5,
        VN2CN0_bit => VN_data_out(7068),
        VN2CN1_bit => VN_data_out(7069),
        VN2CN2_bit => VN_data_out(7070),
        VN2CN3_bit => VN_data_out(7071),
        VN2CN4_bit => VN_data_out(7072),
        VN2CN5_bit => VN_data_out(7073),
        VN2CN0_sign => VN_sign_out(7068),
        VN2CN1_sign => VN_sign_out(7069),
        VN2CN2_sign => VN_sign_out(7070),
        VN2CN3_sign => VN_sign_out(7071),
        VN2CN4_sign => VN_sign_out(7072),
        VN2CN5_sign => VN_sign_out(7073),
        codeword => codeword(1178),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1179 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7079 downto 7074),
        Din0 => VN1179_in0,
        Din1 => VN1179_in1,
        Din2 => VN1179_in2,
        Din3 => VN1179_in3,
        Din4 => VN1179_in4,
        Din5 => VN1179_in5,
        VN2CN0_bit => VN_data_out(7074),
        VN2CN1_bit => VN_data_out(7075),
        VN2CN2_bit => VN_data_out(7076),
        VN2CN3_bit => VN_data_out(7077),
        VN2CN4_bit => VN_data_out(7078),
        VN2CN5_bit => VN_data_out(7079),
        VN2CN0_sign => VN_sign_out(7074),
        VN2CN1_sign => VN_sign_out(7075),
        VN2CN2_sign => VN_sign_out(7076),
        VN2CN3_sign => VN_sign_out(7077),
        VN2CN4_sign => VN_sign_out(7078),
        VN2CN5_sign => VN_sign_out(7079),
        codeword => codeword(1179),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1180 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7085 downto 7080),
        Din0 => VN1180_in0,
        Din1 => VN1180_in1,
        Din2 => VN1180_in2,
        Din3 => VN1180_in3,
        Din4 => VN1180_in4,
        Din5 => VN1180_in5,
        VN2CN0_bit => VN_data_out(7080),
        VN2CN1_bit => VN_data_out(7081),
        VN2CN2_bit => VN_data_out(7082),
        VN2CN3_bit => VN_data_out(7083),
        VN2CN4_bit => VN_data_out(7084),
        VN2CN5_bit => VN_data_out(7085),
        VN2CN0_sign => VN_sign_out(7080),
        VN2CN1_sign => VN_sign_out(7081),
        VN2CN2_sign => VN_sign_out(7082),
        VN2CN3_sign => VN_sign_out(7083),
        VN2CN4_sign => VN_sign_out(7084),
        VN2CN5_sign => VN_sign_out(7085),
        codeword => codeword(1180),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1181 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7091 downto 7086),
        Din0 => VN1181_in0,
        Din1 => VN1181_in1,
        Din2 => VN1181_in2,
        Din3 => VN1181_in3,
        Din4 => VN1181_in4,
        Din5 => VN1181_in5,
        VN2CN0_bit => VN_data_out(7086),
        VN2CN1_bit => VN_data_out(7087),
        VN2CN2_bit => VN_data_out(7088),
        VN2CN3_bit => VN_data_out(7089),
        VN2CN4_bit => VN_data_out(7090),
        VN2CN5_bit => VN_data_out(7091),
        VN2CN0_sign => VN_sign_out(7086),
        VN2CN1_sign => VN_sign_out(7087),
        VN2CN2_sign => VN_sign_out(7088),
        VN2CN3_sign => VN_sign_out(7089),
        VN2CN4_sign => VN_sign_out(7090),
        VN2CN5_sign => VN_sign_out(7091),
        codeword => codeword(1181),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1182 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7097 downto 7092),
        Din0 => VN1182_in0,
        Din1 => VN1182_in1,
        Din2 => VN1182_in2,
        Din3 => VN1182_in3,
        Din4 => VN1182_in4,
        Din5 => VN1182_in5,
        VN2CN0_bit => VN_data_out(7092),
        VN2CN1_bit => VN_data_out(7093),
        VN2CN2_bit => VN_data_out(7094),
        VN2CN3_bit => VN_data_out(7095),
        VN2CN4_bit => VN_data_out(7096),
        VN2CN5_bit => VN_data_out(7097),
        VN2CN0_sign => VN_sign_out(7092),
        VN2CN1_sign => VN_sign_out(7093),
        VN2CN2_sign => VN_sign_out(7094),
        VN2CN3_sign => VN_sign_out(7095),
        VN2CN4_sign => VN_sign_out(7096),
        VN2CN5_sign => VN_sign_out(7097),
        codeword => codeword(1182),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1183 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7103 downto 7098),
        Din0 => VN1183_in0,
        Din1 => VN1183_in1,
        Din2 => VN1183_in2,
        Din3 => VN1183_in3,
        Din4 => VN1183_in4,
        Din5 => VN1183_in5,
        VN2CN0_bit => VN_data_out(7098),
        VN2CN1_bit => VN_data_out(7099),
        VN2CN2_bit => VN_data_out(7100),
        VN2CN3_bit => VN_data_out(7101),
        VN2CN4_bit => VN_data_out(7102),
        VN2CN5_bit => VN_data_out(7103),
        VN2CN0_sign => VN_sign_out(7098),
        VN2CN1_sign => VN_sign_out(7099),
        VN2CN2_sign => VN_sign_out(7100),
        VN2CN3_sign => VN_sign_out(7101),
        VN2CN4_sign => VN_sign_out(7102),
        VN2CN5_sign => VN_sign_out(7103),
        codeword => codeword(1183),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1184 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7109 downto 7104),
        Din0 => VN1184_in0,
        Din1 => VN1184_in1,
        Din2 => VN1184_in2,
        Din3 => VN1184_in3,
        Din4 => VN1184_in4,
        Din5 => VN1184_in5,
        VN2CN0_bit => VN_data_out(7104),
        VN2CN1_bit => VN_data_out(7105),
        VN2CN2_bit => VN_data_out(7106),
        VN2CN3_bit => VN_data_out(7107),
        VN2CN4_bit => VN_data_out(7108),
        VN2CN5_bit => VN_data_out(7109),
        VN2CN0_sign => VN_sign_out(7104),
        VN2CN1_sign => VN_sign_out(7105),
        VN2CN2_sign => VN_sign_out(7106),
        VN2CN3_sign => VN_sign_out(7107),
        VN2CN4_sign => VN_sign_out(7108),
        VN2CN5_sign => VN_sign_out(7109),
        codeword => codeword(1184),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1185 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7115 downto 7110),
        Din0 => VN1185_in0,
        Din1 => VN1185_in1,
        Din2 => VN1185_in2,
        Din3 => VN1185_in3,
        Din4 => VN1185_in4,
        Din5 => VN1185_in5,
        VN2CN0_bit => VN_data_out(7110),
        VN2CN1_bit => VN_data_out(7111),
        VN2CN2_bit => VN_data_out(7112),
        VN2CN3_bit => VN_data_out(7113),
        VN2CN4_bit => VN_data_out(7114),
        VN2CN5_bit => VN_data_out(7115),
        VN2CN0_sign => VN_sign_out(7110),
        VN2CN1_sign => VN_sign_out(7111),
        VN2CN2_sign => VN_sign_out(7112),
        VN2CN3_sign => VN_sign_out(7113),
        VN2CN4_sign => VN_sign_out(7114),
        VN2CN5_sign => VN_sign_out(7115),
        codeword => codeword(1185),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1186 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7121 downto 7116),
        Din0 => VN1186_in0,
        Din1 => VN1186_in1,
        Din2 => VN1186_in2,
        Din3 => VN1186_in3,
        Din4 => VN1186_in4,
        Din5 => VN1186_in5,
        VN2CN0_bit => VN_data_out(7116),
        VN2CN1_bit => VN_data_out(7117),
        VN2CN2_bit => VN_data_out(7118),
        VN2CN3_bit => VN_data_out(7119),
        VN2CN4_bit => VN_data_out(7120),
        VN2CN5_bit => VN_data_out(7121),
        VN2CN0_sign => VN_sign_out(7116),
        VN2CN1_sign => VN_sign_out(7117),
        VN2CN2_sign => VN_sign_out(7118),
        VN2CN3_sign => VN_sign_out(7119),
        VN2CN4_sign => VN_sign_out(7120),
        VN2CN5_sign => VN_sign_out(7121),
        codeword => codeword(1186),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1187 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7127 downto 7122),
        Din0 => VN1187_in0,
        Din1 => VN1187_in1,
        Din2 => VN1187_in2,
        Din3 => VN1187_in3,
        Din4 => VN1187_in4,
        Din5 => VN1187_in5,
        VN2CN0_bit => VN_data_out(7122),
        VN2CN1_bit => VN_data_out(7123),
        VN2CN2_bit => VN_data_out(7124),
        VN2CN3_bit => VN_data_out(7125),
        VN2CN4_bit => VN_data_out(7126),
        VN2CN5_bit => VN_data_out(7127),
        VN2CN0_sign => VN_sign_out(7122),
        VN2CN1_sign => VN_sign_out(7123),
        VN2CN2_sign => VN_sign_out(7124),
        VN2CN3_sign => VN_sign_out(7125),
        VN2CN4_sign => VN_sign_out(7126),
        VN2CN5_sign => VN_sign_out(7127),
        codeword => codeword(1187),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1188 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7133 downto 7128),
        Din0 => VN1188_in0,
        Din1 => VN1188_in1,
        Din2 => VN1188_in2,
        Din3 => VN1188_in3,
        Din4 => VN1188_in4,
        Din5 => VN1188_in5,
        VN2CN0_bit => VN_data_out(7128),
        VN2CN1_bit => VN_data_out(7129),
        VN2CN2_bit => VN_data_out(7130),
        VN2CN3_bit => VN_data_out(7131),
        VN2CN4_bit => VN_data_out(7132),
        VN2CN5_bit => VN_data_out(7133),
        VN2CN0_sign => VN_sign_out(7128),
        VN2CN1_sign => VN_sign_out(7129),
        VN2CN2_sign => VN_sign_out(7130),
        VN2CN3_sign => VN_sign_out(7131),
        VN2CN4_sign => VN_sign_out(7132),
        VN2CN5_sign => VN_sign_out(7133),
        codeword => codeword(1188),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1189 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7139 downto 7134),
        Din0 => VN1189_in0,
        Din1 => VN1189_in1,
        Din2 => VN1189_in2,
        Din3 => VN1189_in3,
        Din4 => VN1189_in4,
        Din5 => VN1189_in5,
        VN2CN0_bit => VN_data_out(7134),
        VN2CN1_bit => VN_data_out(7135),
        VN2CN2_bit => VN_data_out(7136),
        VN2CN3_bit => VN_data_out(7137),
        VN2CN4_bit => VN_data_out(7138),
        VN2CN5_bit => VN_data_out(7139),
        VN2CN0_sign => VN_sign_out(7134),
        VN2CN1_sign => VN_sign_out(7135),
        VN2CN2_sign => VN_sign_out(7136),
        VN2CN3_sign => VN_sign_out(7137),
        VN2CN4_sign => VN_sign_out(7138),
        VN2CN5_sign => VN_sign_out(7139),
        codeword => codeword(1189),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1190 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7145 downto 7140),
        Din0 => VN1190_in0,
        Din1 => VN1190_in1,
        Din2 => VN1190_in2,
        Din3 => VN1190_in3,
        Din4 => VN1190_in4,
        Din5 => VN1190_in5,
        VN2CN0_bit => VN_data_out(7140),
        VN2CN1_bit => VN_data_out(7141),
        VN2CN2_bit => VN_data_out(7142),
        VN2CN3_bit => VN_data_out(7143),
        VN2CN4_bit => VN_data_out(7144),
        VN2CN5_bit => VN_data_out(7145),
        VN2CN0_sign => VN_sign_out(7140),
        VN2CN1_sign => VN_sign_out(7141),
        VN2CN2_sign => VN_sign_out(7142),
        VN2CN3_sign => VN_sign_out(7143),
        VN2CN4_sign => VN_sign_out(7144),
        VN2CN5_sign => VN_sign_out(7145),
        codeword => codeword(1190),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1191 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7151 downto 7146),
        Din0 => VN1191_in0,
        Din1 => VN1191_in1,
        Din2 => VN1191_in2,
        Din3 => VN1191_in3,
        Din4 => VN1191_in4,
        Din5 => VN1191_in5,
        VN2CN0_bit => VN_data_out(7146),
        VN2CN1_bit => VN_data_out(7147),
        VN2CN2_bit => VN_data_out(7148),
        VN2CN3_bit => VN_data_out(7149),
        VN2CN4_bit => VN_data_out(7150),
        VN2CN5_bit => VN_data_out(7151),
        VN2CN0_sign => VN_sign_out(7146),
        VN2CN1_sign => VN_sign_out(7147),
        VN2CN2_sign => VN_sign_out(7148),
        VN2CN3_sign => VN_sign_out(7149),
        VN2CN4_sign => VN_sign_out(7150),
        VN2CN5_sign => VN_sign_out(7151),
        codeword => codeword(1191),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1192 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7157 downto 7152),
        Din0 => VN1192_in0,
        Din1 => VN1192_in1,
        Din2 => VN1192_in2,
        Din3 => VN1192_in3,
        Din4 => VN1192_in4,
        Din5 => VN1192_in5,
        VN2CN0_bit => VN_data_out(7152),
        VN2CN1_bit => VN_data_out(7153),
        VN2CN2_bit => VN_data_out(7154),
        VN2CN3_bit => VN_data_out(7155),
        VN2CN4_bit => VN_data_out(7156),
        VN2CN5_bit => VN_data_out(7157),
        VN2CN0_sign => VN_sign_out(7152),
        VN2CN1_sign => VN_sign_out(7153),
        VN2CN2_sign => VN_sign_out(7154),
        VN2CN3_sign => VN_sign_out(7155),
        VN2CN4_sign => VN_sign_out(7156),
        VN2CN5_sign => VN_sign_out(7157),
        codeword => codeword(1192),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1193 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7163 downto 7158),
        Din0 => VN1193_in0,
        Din1 => VN1193_in1,
        Din2 => VN1193_in2,
        Din3 => VN1193_in3,
        Din4 => VN1193_in4,
        Din5 => VN1193_in5,
        VN2CN0_bit => VN_data_out(7158),
        VN2CN1_bit => VN_data_out(7159),
        VN2CN2_bit => VN_data_out(7160),
        VN2CN3_bit => VN_data_out(7161),
        VN2CN4_bit => VN_data_out(7162),
        VN2CN5_bit => VN_data_out(7163),
        VN2CN0_sign => VN_sign_out(7158),
        VN2CN1_sign => VN_sign_out(7159),
        VN2CN2_sign => VN_sign_out(7160),
        VN2CN3_sign => VN_sign_out(7161),
        VN2CN4_sign => VN_sign_out(7162),
        VN2CN5_sign => VN_sign_out(7163),
        codeword => codeword(1193),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1194 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7169 downto 7164),
        Din0 => VN1194_in0,
        Din1 => VN1194_in1,
        Din2 => VN1194_in2,
        Din3 => VN1194_in3,
        Din4 => VN1194_in4,
        Din5 => VN1194_in5,
        VN2CN0_bit => VN_data_out(7164),
        VN2CN1_bit => VN_data_out(7165),
        VN2CN2_bit => VN_data_out(7166),
        VN2CN3_bit => VN_data_out(7167),
        VN2CN4_bit => VN_data_out(7168),
        VN2CN5_bit => VN_data_out(7169),
        VN2CN0_sign => VN_sign_out(7164),
        VN2CN1_sign => VN_sign_out(7165),
        VN2CN2_sign => VN_sign_out(7166),
        VN2CN3_sign => VN_sign_out(7167),
        VN2CN4_sign => VN_sign_out(7168),
        VN2CN5_sign => VN_sign_out(7169),
        codeword => codeword(1194),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1195 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7175 downto 7170),
        Din0 => VN1195_in0,
        Din1 => VN1195_in1,
        Din2 => VN1195_in2,
        Din3 => VN1195_in3,
        Din4 => VN1195_in4,
        Din5 => VN1195_in5,
        VN2CN0_bit => VN_data_out(7170),
        VN2CN1_bit => VN_data_out(7171),
        VN2CN2_bit => VN_data_out(7172),
        VN2CN3_bit => VN_data_out(7173),
        VN2CN4_bit => VN_data_out(7174),
        VN2CN5_bit => VN_data_out(7175),
        VN2CN0_sign => VN_sign_out(7170),
        VN2CN1_sign => VN_sign_out(7171),
        VN2CN2_sign => VN_sign_out(7172),
        VN2CN3_sign => VN_sign_out(7173),
        VN2CN4_sign => VN_sign_out(7174),
        VN2CN5_sign => VN_sign_out(7175),
        codeword => codeword(1195),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1196 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7181 downto 7176),
        Din0 => VN1196_in0,
        Din1 => VN1196_in1,
        Din2 => VN1196_in2,
        Din3 => VN1196_in3,
        Din4 => VN1196_in4,
        Din5 => VN1196_in5,
        VN2CN0_bit => VN_data_out(7176),
        VN2CN1_bit => VN_data_out(7177),
        VN2CN2_bit => VN_data_out(7178),
        VN2CN3_bit => VN_data_out(7179),
        VN2CN4_bit => VN_data_out(7180),
        VN2CN5_bit => VN_data_out(7181),
        VN2CN0_sign => VN_sign_out(7176),
        VN2CN1_sign => VN_sign_out(7177),
        VN2CN2_sign => VN_sign_out(7178),
        VN2CN3_sign => VN_sign_out(7179),
        VN2CN4_sign => VN_sign_out(7180),
        VN2CN5_sign => VN_sign_out(7181),
        codeword => codeword(1196),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1197 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7187 downto 7182),
        Din0 => VN1197_in0,
        Din1 => VN1197_in1,
        Din2 => VN1197_in2,
        Din3 => VN1197_in3,
        Din4 => VN1197_in4,
        Din5 => VN1197_in5,
        VN2CN0_bit => VN_data_out(7182),
        VN2CN1_bit => VN_data_out(7183),
        VN2CN2_bit => VN_data_out(7184),
        VN2CN3_bit => VN_data_out(7185),
        VN2CN4_bit => VN_data_out(7186),
        VN2CN5_bit => VN_data_out(7187),
        VN2CN0_sign => VN_sign_out(7182),
        VN2CN1_sign => VN_sign_out(7183),
        VN2CN2_sign => VN_sign_out(7184),
        VN2CN3_sign => VN_sign_out(7185),
        VN2CN4_sign => VN_sign_out(7186),
        VN2CN5_sign => VN_sign_out(7187),
        codeword => codeword(1197),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1198 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7193 downto 7188),
        Din0 => VN1198_in0,
        Din1 => VN1198_in1,
        Din2 => VN1198_in2,
        Din3 => VN1198_in3,
        Din4 => VN1198_in4,
        Din5 => VN1198_in5,
        VN2CN0_bit => VN_data_out(7188),
        VN2CN1_bit => VN_data_out(7189),
        VN2CN2_bit => VN_data_out(7190),
        VN2CN3_bit => VN_data_out(7191),
        VN2CN4_bit => VN_data_out(7192),
        VN2CN5_bit => VN_data_out(7193),
        VN2CN0_sign => VN_sign_out(7188),
        VN2CN1_sign => VN_sign_out(7189),
        VN2CN2_sign => VN_sign_out(7190),
        VN2CN3_sign => VN_sign_out(7191),
        VN2CN4_sign => VN_sign_out(7192),
        VN2CN5_sign => VN_sign_out(7193),
        codeword => codeword(1198),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1199 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7199 downto 7194),
        Din0 => VN1199_in0,
        Din1 => VN1199_in1,
        Din2 => VN1199_in2,
        Din3 => VN1199_in3,
        Din4 => VN1199_in4,
        Din5 => VN1199_in5,
        VN2CN0_bit => VN_data_out(7194),
        VN2CN1_bit => VN_data_out(7195),
        VN2CN2_bit => VN_data_out(7196),
        VN2CN3_bit => VN_data_out(7197),
        VN2CN4_bit => VN_data_out(7198),
        VN2CN5_bit => VN_data_out(7199),
        VN2CN0_sign => VN_sign_out(7194),
        VN2CN1_sign => VN_sign_out(7195),
        VN2CN2_sign => VN_sign_out(7196),
        VN2CN3_sign => VN_sign_out(7197),
        VN2CN4_sign => VN_sign_out(7198),
        VN2CN5_sign => VN_sign_out(7199),
        codeword => codeword(1199),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1200 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7205 downto 7200),
        Din0 => VN1200_in0,
        Din1 => VN1200_in1,
        Din2 => VN1200_in2,
        Din3 => VN1200_in3,
        Din4 => VN1200_in4,
        Din5 => VN1200_in5,
        VN2CN0_bit => VN_data_out(7200),
        VN2CN1_bit => VN_data_out(7201),
        VN2CN2_bit => VN_data_out(7202),
        VN2CN3_bit => VN_data_out(7203),
        VN2CN4_bit => VN_data_out(7204),
        VN2CN5_bit => VN_data_out(7205),
        VN2CN0_sign => VN_sign_out(7200),
        VN2CN1_sign => VN_sign_out(7201),
        VN2CN2_sign => VN_sign_out(7202),
        VN2CN3_sign => VN_sign_out(7203),
        VN2CN4_sign => VN_sign_out(7204),
        VN2CN5_sign => VN_sign_out(7205),
        codeword => codeword(1200),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1201 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7211 downto 7206),
        Din0 => VN1201_in0,
        Din1 => VN1201_in1,
        Din2 => VN1201_in2,
        Din3 => VN1201_in3,
        Din4 => VN1201_in4,
        Din5 => VN1201_in5,
        VN2CN0_bit => VN_data_out(7206),
        VN2CN1_bit => VN_data_out(7207),
        VN2CN2_bit => VN_data_out(7208),
        VN2CN3_bit => VN_data_out(7209),
        VN2CN4_bit => VN_data_out(7210),
        VN2CN5_bit => VN_data_out(7211),
        VN2CN0_sign => VN_sign_out(7206),
        VN2CN1_sign => VN_sign_out(7207),
        VN2CN2_sign => VN_sign_out(7208),
        VN2CN3_sign => VN_sign_out(7209),
        VN2CN4_sign => VN_sign_out(7210),
        VN2CN5_sign => VN_sign_out(7211),
        codeword => codeword(1201),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1202 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7217 downto 7212),
        Din0 => VN1202_in0,
        Din1 => VN1202_in1,
        Din2 => VN1202_in2,
        Din3 => VN1202_in3,
        Din4 => VN1202_in4,
        Din5 => VN1202_in5,
        VN2CN0_bit => VN_data_out(7212),
        VN2CN1_bit => VN_data_out(7213),
        VN2CN2_bit => VN_data_out(7214),
        VN2CN3_bit => VN_data_out(7215),
        VN2CN4_bit => VN_data_out(7216),
        VN2CN5_bit => VN_data_out(7217),
        VN2CN0_sign => VN_sign_out(7212),
        VN2CN1_sign => VN_sign_out(7213),
        VN2CN2_sign => VN_sign_out(7214),
        VN2CN3_sign => VN_sign_out(7215),
        VN2CN4_sign => VN_sign_out(7216),
        VN2CN5_sign => VN_sign_out(7217),
        codeword => codeword(1202),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1203 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7223 downto 7218),
        Din0 => VN1203_in0,
        Din1 => VN1203_in1,
        Din2 => VN1203_in2,
        Din3 => VN1203_in3,
        Din4 => VN1203_in4,
        Din5 => VN1203_in5,
        VN2CN0_bit => VN_data_out(7218),
        VN2CN1_bit => VN_data_out(7219),
        VN2CN2_bit => VN_data_out(7220),
        VN2CN3_bit => VN_data_out(7221),
        VN2CN4_bit => VN_data_out(7222),
        VN2CN5_bit => VN_data_out(7223),
        VN2CN0_sign => VN_sign_out(7218),
        VN2CN1_sign => VN_sign_out(7219),
        VN2CN2_sign => VN_sign_out(7220),
        VN2CN3_sign => VN_sign_out(7221),
        VN2CN4_sign => VN_sign_out(7222),
        VN2CN5_sign => VN_sign_out(7223),
        codeword => codeword(1203),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1204 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7229 downto 7224),
        Din0 => VN1204_in0,
        Din1 => VN1204_in1,
        Din2 => VN1204_in2,
        Din3 => VN1204_in3,
        Din4 => VN1204_in4,
        Din5 => VN1204_in5,
        VN2CN0_bit => VN_data_out(7224),
        VN2CN1_bit => VN_data_out(7225),
        VN2CN2_bit => VN_data_out(7226),
        VN2CN3_bit => VN_data_out(7227),
        VN2CN4_bit => VN_data_out(7228),
        VN2CN5_bit => VN_data_out(7229),
        VN2CN0_sign => VN_sign_out(7224),
        VN2CN1_sign => VN_sign_out(7225),
        VN2CN2_sign => VN_sign_out(7226),
        VN2CN3_sign => VN_sign_out(7227),
        VN2CN4_sign => VN_sign_out(7228),
        VN2CN5_sign => VN_sign_out(7229),
        codeword => codeword(1204),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1205 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7235 downto 7230),
        Din0 => VN1205_in0,
        Din1 => VN1205_in1,
        Din2 => VN1205_in2,
        Din3 => VN1205_in3,
        Din4 => VN1205_in4,
        Din5 => VN1205_in5,
        VN2CN0_bit => VN_data_out(7230),
        VN2CN1_bit => VN_data_out(7231),
        VN2CN2_bit => VN_data_out(7232),
        VN2CN3_bit => VN_data_out(7233),
        VN2CN4_bit => VN_data_out(7234),
        VN2CN5_bit => VN_data_out(7235),
        VN2CN0_sign => VN_sign_out(7230),
        VN2CN1_sign => VN_sign_out(7231),
        VN2CN2_sign => VN_sign_out(7232),
        VN2CN3_sign => VN_sign_out(7233),
        VN2CN4_sign => VN_sign_out(7234),
        VN2CN5_sign => VN_sign_out(7235),
        codeword => codeword(1205),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1206 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7241 downto 7236),
        Din0 => VN1206_in0,
        Din1 => VN1206_in1,
        Din2 => VN1206_in2,
        Din3 => VN1206_in3,
        Din4 => VN1206_in4,
        Din5 => VN1206_in5,
        VN2CN0_bit => VN_data_out(7236),
        VN2CN1_bit => VN_data_out(7237),
        VN2CN2_bit => VN_data_out(7238),
        VN2CN3_bit => VN_data_out(7239),
        VN2CN4_bit => VN_data_out(7240),
        VN2CN5_bit => VN_data_out(7241),
        VN2CN0_sign => VN_sign_out(7236),
        VN2CN1_sign => VN_sign_out(7237),
        VN2CN2_sign => VN_sign_out(7238),
        VN2CN3_sign => VN_sign_out(7239),
        VN2CN4_sign => VN_sign_out(7240),
        VN2CN5_sign => VN_sign_out(7241),
        codeword => codeword(1206),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1207 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7247 downto 7242),
        Din0 => VN1207_in0,
        Din1 => VN1207_in1,
        Din2 => VN1207_in2,
        Din3 => VN1207_in3,
        Din4 => VN1207_in4,
        Din5 => VN1207_in5,
        VN2CN0_bit => VN_data_out(7242),
        VN2CN1_bit => VN_data_out(7243),
        VN2CN2_bit => VN_data_out(7244),
        VN2CN3_bit => VN_data_out(7245),
        VN2CN4_bit => VN_data_out(7246),
        VN2CN5_bit => VN_data_out(7247),
        VN2CN0_sign => VN_sign_out(7242),
        VN2CN1_sign => VN_sign_out(7243),
        VN2CN2_sign => VN_sign_out(7244),
        VN2CN3_sign => VN_sign_out(7245),
        VN2CN4_sign => VN_sign_out(7246),
        VN2CN5_sign => VN_sign_out(7247),
        codeword => codeword(1207),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1208 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7253 downto 7248),
        Din0 => VN1208_in0,
        Din1 => VN1208_in1,
        Din2 => VN1208_in2,
        Din3 => VN1208_in3,
        Din4 => VN1208_in4,
        Din5 => VN1208_in5,
        VN2CN0_bit => VN_data_out(7248),
        VN2CN1_bit => VN_data_out(7249),
        VN2CN2_bit => VN_data_out(7250),
        VN2CN3_bit => VN_data_out(7251),
        VN2CN4_bit => VN_data_out(7252),
        VN2CN5_bit => VN_data_out(7253),
        VN2CN0_sign => VN_sign_out(7248),
        VN2CN1_sign => VN_sign_out(7249),
        VN2CN2_sign => VN_sign_out(7250),
        VN2CN3_sign => VN_sign_out(7251),
        VN2CN4_sign => VN_sign_out(7252),
        VN2CN5_sign => VN_sign_out(7253),
        codeword => codeword(1208),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1209 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7259 downto 7254),
        Din0 => VN1209_in0,
        Din1 => VN1209_in1,
        Din2 => VN1209_in2,
        Din3 => VN1209_in3,
        Din4 => VN1209_in4,
        Din5 => VN1209_in5,
        VN2CN0_bit => VN_data_out(7254),
        VN2CN1_bit => VN_data_out(7255),
        VN2CN2_bit => VN_data_out(7256),
        VN2CN3_bit => VN_data_out(7257),
        VN2CN4_bit => VN_data_out(7258),
        VN2CN5_bit => VN_data_out(7259),
        VN2CN0_sign => VN_sign_out(7254),
        VN2CN1_sign => VN_sign_out(7255),
        VN2CN2_sign => VN_sign_out(7256),
        VN2CN3_sign => VN_sign_out(7257),
        VN2CN4_sign => VN_sign_out(7258),
        VN2CN5_sign => VN_sign_out(7259),
        codeword => codeword(1209),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1210 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7265 downto 7260),
        Din0 => VN1210_in0,
        Din1 => VN1210_in1,
        Din2 => VN1210_in2,
        Din3 => VN1210_in3,
        Din4 => VN1210_in4,
        Din5 => VN1210_in5,
        VN2CN0_bit => VN_data_out(7260),
        VN2CN1_bit => VN_data_out(7261),
        VN2CN2_bit => VN_data_out(7262),
        VN2CN3_bit => VN_data_out(7263),
        VN2CN4_bit => VN_data_out(7264),
        VN2CN5_bit => VN_data_out(7265),
        VN2CN0_sign => VN_sign_out(7260),
        VN2CN1_sign => VN_sign_out(7261),
        VN2CN2_sign => VN_sign_out(7262),
        VN2CN3_sign => VN_sign_out(7263),
        VN2CN4_sign => VN_sign_out(7264),
        VN2CN5_sign => VN_sign_out(7265),
        codeword => codeword(1210),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1211 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7271 downto 7266),
        Din0 => VN1211_in0,
        Din1 => VN1211_in1,
        Din2 => VN1211_in2,
        Din3 => VN1211_in3,
        Din4 => VN1211_in4,
        Din5 => VN1211_in5,
        VN2CN0_bit => VN_data_out(7266),
        VN2CN1_bit => VN_data_out(7267),
        VN2CN2_bit => VN_data_out(7268),
        VN2CN3_bit => VN_data_out(7269),
        VN2CN4_bit => VN_data_out(7270),
        VN2CN5_bit => VN_data_out(7271),
        VN2CN0_sign => VN_sign_out(7266),
        VN2CN1_sign => VN_sign_out(7267),
        VN2CN2_sign => VN_sign_out(7268),
        VN2CN3_sign => VN_sign_out(7269),
        VN2CN4_sign => VN_sign_out(7270),
        VN2CN5_sign => VN_sign_out(7271),
        codeword => codeword(1211),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1212 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7277 downto 7272),
        Din0 => VN1212_in0,
        Din1 => VN1212_in1,
        Din2 => VN1212_in2,
        Din3 => VN1212_in3,
        Din4 => VN1212_in4,
        Din5 => VN1212_in5,
        VN2CN0_bit => VN_data_out(7272),
        VN2CN1_bit => VN_data_out(7273),
        VN2CN2_bit => VN_data_out(7274),
        VN2CN3_bit => VN_data_out(7275),
        VN2CN4_bit => VN_data_out(7276),
        VN2CN5_bit => VN_data_out(7277),
        VN2CN0_sign => VN_sign_out(7272),
        VN2CN1_sign => VN_sign_out(7273),
        VN2CN2_sign => VN_sign_out(7274),
        VN2CN3_sign => VN_sign_out(7275),
        VN2CN4_sign => VN_sign_out(7276),
        VN2CN5_sign => VN_sign_out(7277),
        codeword => codeword(1212),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1213 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7283 downto 7278),
        Din0 => VN1213_in0,
        Din1 => VN1213_in1,
        Din2 => VN1213_in2,
        Din3 => VN1213_in3,
        Din4 => VN1213_in4,
        Din5 => VN1213_in5,
        VN2CN0_bit => VN_data_out(7278),
        VN2CN1_bit => VN_data_out(7279),
        VN2CN2_bit => VN_data_out(7280),
        VN2CN3_bit => VN_data_out(7281),
        VN2CN4_bit => VN_data_out(7282),
        VN2CN5_bit => VN_data_out(7283),
        VN2CN0_sign => VN_sign_out(7278),
        VN2CN1_sign => VN_sign_out(7279),
        VN2CN2_sign => VN_sign_out(7280),
        VN2CN3_sign => VN_sign_out(7281),
        VN2CN4_sign => VN_sign_out(7282),
        VN2CN5_sign => VN_sign_out(7283),
        codeword => codeword(1213),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1214 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7289 downto 7284),
        Din0 => VN1214_in0,
        Din1 => VN1214_in1,
        Din2 => VN1214_in2,
        Din3 => VN1214_in3,
        Din4 => VN1214_in4,
        Din5 => VN1214_in5,
        VN2CN0_bit => VN_data_out(7284),
        VN2CN1_bit => VN_data_out(7285),
        VN2CN2_bit => VN_data_out(7286),
        VN2CN3_bit => VN_data_out(7287),
        VN2CN4_bit => VN_data_out(7288),
        VN2CN5_bit => VN_data_out(7289),
        VN2CN0_sign => VN_sign_out(7284),
        VN2CN1_sign => VN_sign_out(7285),
        VN2CN2_sign => VN_sign_out(7286),
        VN2CN3_sign => VN_sign_out(7287),
        VN2CN4_sign => VN_sign_out(7288),
        VN2CN5_sign => VN_sign_out(7289),
        codeword => codeword(1214),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1215 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7295 downto 7290),
        Din0 => VN1215_in0,
        Din1 => VN1215_in1,
        Din2 => VN1215_in2,
        Din3 => VN1215_in3,
        Din4 => VN1215_in4,
        Din5 => VN1215_in5,
        VN2CN0_bit => VN_data_out(7290),
        VN2CN1_bit => VN_data_out(7291),
        VN2CN2_bit => VN_data_out(7292),
        VN2CN3_bit => VN_data_out(7293),
        VN2CN4_bit => VN_data_out(7294),
        VN2CN5_bit => VN_data_out(7295),
        VN2CN0_sign => VN_sign_out(7290),
        VN2CN1_sign => VN_sign_out(7291),
        VN2CN2_sign => VN_sign_out(7292),
        VN2CN3_sign => VN_sign_out(7293),
        VN2CN4_sign => VN_sign_out(7294),
        VN2CN5_sign => VN_sign_out(7295),
        codeword => codeword(1215),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1216 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7301 downto 7296),
        Din0 => VN1216_in0,
        Din1 => VN1216_in1,
        Din2 => VN1216_in2,
        Din3 => VN1216_in3,
        Din4 => VN1216_in4,
        Din5 => VN1216_in5,
        VN2CN0_bit => VN_data_out(7296),
        VN2CN1_bit => VN_data_out(7297),
        VN2CN2_bit => VN_data_out(7298),
        VN2CN3_bit => VN_data_out(7299),
        VN2CN4_bit => VN_data_out(7300),
        VN2CN5_bit => VN_data_out(7301),
        VN2CN0_sign => VN_sign_out(7296),
        VN2CN1_sign => VN_sign_out(7297),
        VN2CN2_sign => VN_sign_out(7298),
        VN2CN3_sign => VN_sign_out(7299),
        VN2CN4_sign => VN_sign_out(7300),
        VN2CN5_sign => VN_sign_out(7301),
        codeword => codeword(1216),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1217 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7307 downto 7302),
        Din0 => VN1217_in0,
        Din1 => VN1217_in1,
        Din2 => VN1217_in2,
        Din3 => VN1217_in3,
        Din4 => VN1217_in4,
        Din5 => VN1217_in5,
        VN2CN0_bit => VN_data_out(7302),
        VN2CN1_bit => VN_data_out(7303),
        VN2CN2_bit => VN_data_out(7304),
        VN2CN3_bit => VN_data_out(7305),
        VN2CN4_bit => VN_data_out(7306),
        VN2CN5_bit => VN_data_out(7307),
        VN2CN0_sign => VN_sign_out(7302),
        VN2CN1_sign => VN_sign_out(7303),
        VN2CN2_sign => VN_sign_out(7304),
        VN2CN3_sign => VN_sign_out(7305),
        VN2CN4_sign => VN_sign_out(7306),
        VN2CN5_sign => VN_sign_out(7307),
        codeword => codeword(1217),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1218 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7313 downto 7308),
        Din0 => VN1218_in0,
        Din1 => VN1218_in1,
        Din2 => VN1218_in2,
        Din3 => VN1218_in3,
        Din4 => VN1218_in4,
        Din5 => VN1218_in5,
        VN2CN0_bit => VN_data_out(7308),
        VN2CN1_bit => VN_data_out(7309),
        VN2CN2_bit => VN_data_out(7310),
        VN2CN3_bit => VN_data_out(7311),
        VN2CN4_bit => VN_data_out(7312),
        VN2CN5_bit => VN_data_out(7313),
        VN2CN0_sign => VN_sign_out(7308),
        VN2CN1_sign => VN_sign_out(7309),
        VN2CN2_sign => VN_sign_out(7310),
        VN2CN3_sign => VN_sign_out(7311),
        VN2CN4_sign => VN_sign_out(7312),
        VN2CN5_sign => VN_sign_out(7313),
        codeword => codeword(1218),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1219 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7319 downto 7314),
        Din0 => VN1219_in0,
        Din1 => VN1219_in1,
        Din2 => VN1219_in2,
        Din3 => VN1219_in3,
        Din4 => VN1219_in4,
        Din5 => VN1219_in5,
        VN2CN0_bit => VN_data_out(7314),
        VN2CN1_bit => VN_data_out(7315),
        VN2CN2_bit => VN_data_out(7316),
        VN2CN3_bit => VN_data_out(7317),
        VN2CN4_bit => VN_data_out(7318),
        VN2CN5_bit => VN_data_out(7319),
        VN2CN0_sign => VN_sign_out(7314),
        VN2CN1_sign => VN_sign_out(7315),
        VN2CN2_sign => VN_sign_out(7316),
        VN2CN3_sign => VN_sign_out(7317),
        VN2CN4_sign => VN_sign_out(7318),
        VN2CN5_sign => VN_sign_out(7319),
        codeword => codeword(1219),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1220 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7325 downto 7320),
        Din0 => VN1220_in0,
        Din1 => VN1220_in1,
        Din2 => VN1220_in2,
        Din3 => VN1220_in3,
        Din4 => VN1220_in4,
        Din5 => VN1220_in5,
        VN2CN0_bit => VN_data_out(7320),
        VN2CN1_bit => VN_data_out(7321),
        VN2CN2_bit => VN_data_out(7322),
        VN2CN3_bit => VN_data_out(7323),
        VN2CN4_bit => VN_data_out(7324),
        VN2CN5_bit => VN_data_out(7325),
        VN2CN0_sign => VN_sign_out(7320),
        VN2CN1_sign => VN_sign_out(7321),
        VN2CN2_sign => VN_sign_out(7322),
        VN2CN3_sign => VN_sign_out(7323),
        VN2CN4_sign => VN_sign_out(7324),
        VN2CN5_sign => VN_sign_out(7325),
        codeword => codeword(1220),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1221 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7331 downto 7326),
        Din0 => VN1221_in0,
        Din1 => VN1221_in1,
        Din2 => VN1221_in2,
        Din3 => VN1221_in3,
        Din4 => VN1221_in4,
        Din5 => VN1221_in5,
        VN2CN0_bit => VN_data_out(7326),
        VN2CN1_bit => VN_data_out(7327),
        VN2CN2_bit => VN_data_out(7328),
        VN2CN3_bit => VN_data_out(7329),
        VN2CN4_bit => VN_data_out(7330),
        VN2CN5_bit => VN_data_out(7331),
        VN2CN0_sign => VN_sign_out(7326),
        VN2CN1_sign => VN_sign_out(7327),
        VN2CN2_sign => VN_sign_out(7328),
        VN2CN3_sign => VN_sign_out(7329),
        VN2CN4_sign => VN_sign_out(7330),
        VN2CN5_sign => VN_sign_out(7331),
        codeword => codeword(1221),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1222 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7337 downto 7332),
        Din0 => VN1222_in0,
        Din1 => VN1222_in1,
        Din2 => VN1222_in2,
        Din3 => VN1222_in3,
        Din4 => VN1222_in4,
        Din5 => VN1222_in5,
        VN2CN0_bit => VN_data_out(7332),
        VN2CN1_bit => VN_data_out(7333),
        VN2CN2_bit => VN_data_out(7334),
        VN2CN3_bit => VN_data_out(7335),
        VN2CN4_bit => VN_data_out(7336),
        VN2CN5_bit => VN_data_out(7337),
        VN2CN0_sign => VN_sign_out(7332),
        VN2CN1_sign => VN_sign_out(7333),
        VN2CN2_sign => VN_sign_out(7334),
        VN2CN3_sign => VN_sign_out(7335),
        VN2CN4_sign => VN_sign_out(7336),
        VN2CN5_sign => VN_sign_out(7337),
        codeword => codeword(1222),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1223 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7343 downto 7338),
        Din0 => VN1223_in0,
        Din1 => VN1223_in1,
        Din2 => VN1223_in2,
        Din3 => VN1223_in3,
        Din4 => VN1223_in4,
        Din5 => VN1223_in5,
        VN2CN0_bit => VN_data_out(7338),
        VN2CN1_bit => VN_data_out(7339),
        VN2CN2_bit => VN_data_out(7340),
        VN2CN3_bit => VN_data_out(7341),
        VN2CN4_bit => VN_data_out(7342),
        VN2CN5_bit => VN_data_out(7343),
        VN2CN0_sign => VN_sign_out(7338),
        VN2CN1_sign => VN_sign_out(7339),
        VN2CN2_sign => VN_sign_out(7340),
        VN2CN3_sign => VN_sign_out(7341),
        VN2CN4_sign => VN_sign_out(7342),
        VN2CN5_sign => VN_sign_out(7343),
        codeword => codeword(1223),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1224 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7349 downto 7344),
        Din0 => VN1224_in0,
        Din1 => VN1224_in1,
        Din2 => VN1224_in2,
        Din3 => VN1224_in3,
        Din4 => VN1224_in4,
        Din5 => VN1224_in5,
        VN2CN0_bit => VN_data_out(7344),
        VN2CN1_bit => VN_data_out(7345),
        VN2CN2_bit => VN_data_out(7346),
        VN2CN3_bit => VN_data_out(7347),
        VN2CN4_bit => VN_data_out(7348),
        VN2CN5_bit => VN_data_out(7349),
        VN2CN0_sign => VN_sign_out(7344),
        VN2CN1_sign => VN_sign_out(7345),
        VN2CN2_sign => VN_sign_out(7346),
        VN2CN3_sign => VN_sign_out(7347),
        VN2CN4_sign => VN_sign_out(7348),
        VN2CN5_sign => VN_sign_out(7349),
        codeword => codeword(1224),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1225 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7355 downto 7350),
        Din0 => VN1225_in0,
        Din1 => VN1225_in1,
        Din2 => VN1225_in2,
        Din3 => VN1225_in3,
        Din4 => VN1225_in4,
        Din5 => VN1225_in5,
        VN2CN0_bit => VN_data_out(7350),
        VN2CN1_bit => VN_data_out(7351),
        VN2CN2_bit => VN_data_out(7352),
        VN2CN3_bit => VN_data_out(7353),
        VN2CN4_bit => VN_data_out(7354),
        VN2CN5_bit => VN_data_out(7355),
        VN2CN0_sign => VN_sign_out(7350),
        VN2CN1_sign => VN_sign_out(7351),
        VN2CN2_sign => VN_sign_out(7352),
        VN2CN3_sign => VN_sign_out(7353),
        VN2CN4_sign => VN_sign_out(7354),
        VN2CN5_sign => VN_sign_out(7355),
        codeword => codeword(1225),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1226 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7361 downto 7356),
        Din0 => VN1226_in0,
        Din1 => VN1226_in1,
        Din2 => VN1226_in2,
        Din3 => VN1226_in3,
        Din4 => VN1226_in4,
        Din5 => VN1226_in5,
        VN2CN0_bit => VN_data_out(7356),
        VN2CN1_bit => VN_data_out(7357),
        VN2CN2_bit => VN_data_out(7358),
        VN2CN3_bit => VN_data_out(7359),
        VN2CN4_bit => VN_data_out(7360),
        VN2CN5_bit => VN_data_out(7361),
        VN2CN0_sign => VN_sign_out(7356),
        VN2CN1_sign => VN_sign_out(7357),
        VN2CN2_sign => VN_sign_out(7358),
        VN2CN3_sign => VN_sign_out(7359),
        VN2CN4_sign => VN_sign_out(7360),
        VN2CN5_sign => VN_sign_out(7361),
        codeword => codeword(1226),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1227 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7367 downto 7362),
        Din0 => VN1227_in0,
        Din1 => VN1227_in1,
        Din2 => VN1227_in2,
        Din3 => VN1227_in3,
        Din4 => VN1227_in4,
        Din5 => VN1227_in5,
        VN2CN0_bit => VN_data_out(7362),
        VN2CN1_bit => VN_data_out(7363),
        VN2CN2_bit => VN_data_out(7364),
        VN2CN3_bit => VN_data_out(7365),
        VN2CN4_bit => VN_data_out(7366),
        VN2CN5_bit => VN_data_out(7367),
        VN2CN0_sign => VN_sign_out(7362),
        VN2CN1_sign => VN_sign_out(7363),
        VN2CN2_sign => VN_sign_out(7364),
        VN2CN3_sign => VN_sign_out(7365),
        VN2CN4_sign => VN_sign_out(7366),
        VN2CN5_sign => VN_sign_out(7367),
        codeword => codeword(1227),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1228 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7373 downto 7368),
        Din0 => VN1228_in0,
        Din1 => VN1228_in1,
        Din2 => VN1228_in2,
        Din3 => VN1228_in3,
        Din4 => VN1228_in4,
        Din5 => VN1228_in5,
        VN2CN0_bit => VN_data_out(7368),
        VN2CN1_bit => VN_data_out(7369),
        VN2CN2_bit => VN_data_out(7370),
        VN2CN3_bit => VN_data_out(7371),
        VN2CN4_bit => VN_data_out(7372),
        VN2CN5_bit => VN_data_out(7373),
        VN2CN0_sign => VN_sign_out(7368),
        VN2CN1_sign => VN_sign_out(7369),
        VN2CN2_sign => VN_sign_out(7370),
        VN2CN3_sign => VN_sign_out(7371),
        VN2CN4_sign => VN_sign_out(7372),
        VN2CN5_sign => VN_sign_out(7373),
        codeword => codeword(1228),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1229 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7379 downto 7374),
        Din0 => VN1229_in0,
        Din1 => VN1229_in1,
        Din2 => VN1229_in2,
        Din3 => VN1229_in3,
        Din4 => VN1229_in4,
        Din5 => VN1229_in5,
        VN2CN0_bit => VN_data_out(7374),
        VN2CN1_bit => VN_data_out(7375),
        VN2CN2_bit => VN_data_out(7376),
        VN2CN3_bit => VN_data_out(7377),
        VN2CN4_bit => VN_data_out(7378),
        VN2CN5_bit => VN_data_out(7379),
        VN2CN0_sign => VN_sign_out(7374),
        VN2CN1_sign => VN_sign_out(7375),
        VN2CN2_sign => VN_sign_out(7376),
        VN2CN3_sign => VN_sign_out(7377),
        VN2CN4_sign => VN_sign_out(7378),
        VN2CN5_sign => VN_sign_out(7379),
        codeword => codeword(1229),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1230 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7385 downto 7380),
        Din0 => VN1230_in0,
        Din1 => VN1230_in1,
        Din2 => VN1230_in2,
        Din3 => VN1230_in3,
        Din4 => VN1230_in4,
        Din5 => VN1230_in5,
        VN2CN0_bit => VN_data_out(7380),
        VN2CN1_bit => VN_data_out(7381),
        VN2CN2_bit => VN_data_out(7382),
        VN2CN3_bit => VN_data_out(7383),
        VN2CN4_bit => VN_data_out(7384),
        VN2CN5_bit => VN_data_out(7385),
        VN2CN0_sign => VN_sign_out(7380),
        VN2CN1_sign => VN_sign_out(7381),
        VN2CN2_sign => VN_sign_out(7382),
        VN2CN3_sign => VN_sign_out(7383),
        VN2CN4_sign => VN_sign_out(7384),
        VN2CN5_sign => VN_sign_out(7385),
        codeword => codeword(1230),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1231 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7391 downto 7386),
        Din0 => VN1231_in0,
        Din1 => VN1231_in1,
        Din2 => VN1231_in2,
        Din3 => VN1231_in3,
        Din4 => VN1231_in4,
        Din5 => VN1231_in5,
        VN2CN0_bit => VN_data_out(7386),
        VN2CN1_bit => VN_data_out(7387),
        VN2CN2_bit => VN_data_out(7388),
        VN2CN3_bit => VN_data_out(7389),
        VN2CN4_bit => VN_data_out(7390),
        VN2CN5_bit => VN_data_out(7391),
        VN2CN0_sign => VN_sign_out(7386),
        VN2CN1_sign => VN_sign_out(7387),
        VN2CN2_sign => VN_sign_out(7388),
        VN2CN3_sign => VN_sign_out(7389),
        VN2CN4_sign => VN_sign_out(7390),
        VN2CN5_sign => VN_sign_out(7391),
        codeword => codeword(1231),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1232 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7397 downto 7392),
        Din0 => VN1232_in0,
        Din1 => VN1232_in1,
        Din2 => VN1232_in2,
        Din3 => VN1232_in3,
        Din4 => VN1232_in4,
        Din5 => VN1232_in5,
        VN2CN0_bit => VN_data_out(7392),
        VN2CN1_bit => VN_data_out(7393),
        VN2CN2_bit => VN_data_out(7394),
        VN2CN3_bit => VN_data_out(7395),
        VN2CN4_bit => VN_data_out(7396),
        VN2CN5_bit => VN_data_out(7397),
        VN2CN0_sign => VN_sign_out(7392),
        VN2CN1_sign => VN_sign_out(7393),
        VN2CN2_sign => VN_sign_out(7394),
        VN2CN3_sign => VN_sign_out(7395),
        VN2CN4_sign => VN_sign_out(7396),
        VN2CN5_sign => VN_sign_out(7397),
        codeword => codeword(1232),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1233 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7403 downto 7398),
        Din0 => VN1233_in0,
        Din1 => VN1233_in1,
        Din2 => VN1233_in2,
        Din3 => VN1233_in3,
        Din4 => VN1233_in4,
        Din5 => VN1233_in5,
        VN2CN0_bit => VN_data_out(7398),
        VN2CN1_bit => VN_data_out(7399),
        VN2CN2_bit => VN_data_out(7400),
        VN2CN3_bit => VN_data_out(7401),
        VN2CN4_bit => VN_data_out(7402),
        VN2CN5_bit => VN_data_out(7403),
        VN2CN0_sign => VN_sign_out(7398),
        VN2CN1_sign => VN_sign_out(7399),
        VN2CN2_sign => VN_sign_out(7400),
        VN2CN3_sign => VN_sign_out(7401),
        VN2CN4_sign => VN_sign_out(7402),
        VN2CN5_sign => VN_sign_out(7403),
        codeword => codeword(1233),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1234 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7409 downto 7404),
        Din0 => VN1234_in0,
        Din1 => VN1234_in1,
        Din2 => VN1234_in2,
        Din3 => VN1234_in3,
        Din4 => VN1234_in4,
        Din5 => VN1234_in5,
        VN2CN0_bit => VN_data_out(7404),
        VN2CN1_bit => VN_data_out(7405),
        VN2CN2_bit => VN_data_out(7406),
        VN2CN3_bit => VN_data_out(7407),
        VN2CN4_bit => VN_data_out(7408),
        VN2CN5_bit => VN_data_out(7409),
        VN2CN0_sign => VN_sign_out(7404),
        VN2CN1_sign => VN_sign_out(7405),
        VN2CN2_sign => VN_sign_out(7406),
        VN2CN3_sign => VN_sign_out(7407),
        VN2CN4_sign => VN_sign_out(7408),
        VN2CN5_sign => VN_sign_out(7409),
        codeword => codeword(1234),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1235 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7415 downto 7410),
        Din0 => VN1235_in0,
        Din1 => VN1235_in1,
        Din2 => VN1235_in2,
        Din3 => VN1235_in3,
        Din4 => VN1235_in4,
        Din5 => VN1235_in5,
        VN2CN0_bit => VN_data_out(7410),
        VN2CN1_bit => VN_data_out(7411),
        VN2CN2_bit => VN_data_out(7412),
        VN2CN3_bit => VN_data_out(7413),
        VN2CN4_bit => VN_data_out(7414),
        VN2CN5_bit => VN_data_out(7415),
        VN2CN0_sign => VN_sign_out(7410),
        VN2CN1_sign => VN_sign_out(7411),
        VN2CN2_sign => VN_sign_out(7412),
        VN2CN3_sign => VN_sign_out(7413),
        VN2CN4_sign => VN_sign_out(7414),
        VN2CN5_sign => VN_sign_out(7415),
        codeword => codeword(1235),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1236 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7421 downto 7416),
        Din0 => VN1236_in0,
        Din1 => VN1236_in1,
        Din2 => VN1236_in2,
        Din3 => VN1236_in3,
        Din4 => VN1236_in4,
        Din5 => VN1236_in5,
        VN2CN0_bit => VN_data_out(7416),
        VN2CN1_bit => VN_data_out(7417),
        VN2CN2_bit => VN_data_out(7418),
        VN2CN3_bit => VN_data_out(7419),
        VN2CN4_bit => VN_data_out(7420),
        VN2CN5_bit => VN_data_out(7421),
        VN2CN0_sign => VN_sign_out(7416),
        VN2CN1_sign => VN_sign_out(7417),
        VN2CN2_sign => VN_sign_out(7418),
        VN2CN3_sign => VN_sign_out(7419),
        VN2CN4_sign => VN_sign_out(7420),
        VN2CN5_sign => VN_sign_out(7421),
        codeword => codeword(1236),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1237 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7427 downto 7422),
        Din0 => VN1237_in0,
        Din1 => VN1237_in1,
        Din2 => VN1237_in2,
        Din3 => VN1237_in3,
        Din4 => VN1237_in4,
        Din5 => VN1237_in5,
        VN2CN0_bit => VN_data_out(7422),
        VN2CN1_bit => VN_data_out(7423),
        VN2CN2_bit => VN_data_out(7424),
        VN2CN3_bit => VN_data_out(7425),
        VN2CN4_bit => VN_data_out(7426),
        VN2CN5_bit => VN_data_out(7427),
        VN2CN0_sign => VN_sign_out(7422),
        VN2CN1_sign => VN_sign_out(7423),
        VN2CN2_sign => VN_sign_out(7424),
        VN2CN3_sign => VN_sign_out(7425),
        VN2CN4_sign => VN_sign_out(7426),
        VN2CN5_sign => VN_sign_out(7427),
        codeword => codeword(1237),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1238 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7433 downto 7428),
        Din0 => VN1238_in0,
        Din1 => VN1238_in1,
        Din2 => VN1238_in2,
        Din3 => VN1238_in3,
        Din4 => VN1238_in4,
        Din5 => VN1238_in5,
        VN2CN0_bit => VN_data_out(7428),
        VN2CN1_bit => VN_data_out(7429),
        VN2CN2_bit => VN_data_out(7430),
        VN2CN3_bit => VN_data_out(7431),
        VN2CN4_bit => VN_data_out(7432),
        VN2CN5_bit => VN_data_out(7433),
        VN2CN0_sign => VN_sign_out(7428),
        VN2CN1_sign => VN_sign_out(7429),
        VN2CN2_sign => VN_sign_out(7430),
        VN2CN3_sign => VN_sign_out(7431),
        VN2CN4_sign => VN_sign_out(7432),
        VN2CN5_sign => VN_sign_out(7433),
        codeword => codeword(1238),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1239 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7439 downto 7434),
        Din0 => VN1239_in0,
        Din1 => VN1239_in1,
        Din2 => VN1239_in2,
        Din3 => VN1239_in3,
        Din4 => VN1239_in4,
        Din5 => VN1239_in5,
        VN2CN0_bit => VN_data_out(7434),
        VN2CN1_bit => VN_data_out(7435),
        VN2CN2_bit => VN_data_out(7436),
        VN2CN3_bit => VN_data_out(7437),
        VN2CN4_bit => VN_data_out(7438),
        VN2CN5_bit => VN_data_out(7439),
        VN2CN0_sign => VN_sign_out(7434),
        VN2CN1_sign => VN_sign_out(7435),
        VN2CN2_sign => VN_sign_out(7436),
        VN2CN3_sign => VN_sign_out(7437),
        VN2CN4_sign => VN_sign_out(7438),
        VN2CN5_sign => VN_sign_out(7439),
        codeword => codeword(1239),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1240 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7445 downto 7440),
        Din0 => VN1240_in0,
        Din1 => VN1240_in1,
        Din2 => VN1240_in2,
        Din3 => VN1240_in3,
        Din4 => VN1240_in4,
        Din5 => VN1240_in5,
        VN2CN0_bit => VN_data_out(7440),
        VN2CN1_bit => VN_data_out(7441),
        VN2CN2_bit => VN_data_out(7442),
        VN2CN3_bit => VN_data_out(7443),
        VN2CN4_bit => VN_data_out(7444),
        VN2CN5_bit => VN_data_out(7445),
        VN2CN0_sign => VN_sign_out(7440),
        VN2CN1_sign => VN_sign_out(7441),
        VN2CN2_sign => VN_sign_out(7442),
        VN2CN3_sign => VN_sign_out(7443),
        VN2CN4_sign => VN_sign_out(7444),
        VN2CN5_sign => VN_sign_out(7445),
        codeword => codeword(1240),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1241 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7451 downto 7446),
        Din0 => VN1241_in0,
        Din1 => VN1241_in1,
        Din2 => VN1241_in2,
        Din3 => VN1241_in3,
        Din4 => VN1241_in4,
        Din5 => VN1241_in5,
        VN2CN0_bit => VN_data_out(7446),
        VN2CN1_bit => VN_data_out(7447),
        VN2CN2_bit => VN_data_out(7448),
        VN2CN3_bit => VN_data_out(7449),
        VN2CN4_bit => VN_data_out(7450),
        VN2CN5_bit => VN_data_out(7451),
        VN2CN0_sign => VN_sign_out(7446),
        VN2CN1_sign => VN_sign_out(7447),
        VN2CN2_sign => VN_sign_out(7448),
        VN2CN3_sign => VN_sign_out(7449),
        VN2CN4_sign => VN_sign_out(7450),
        VN2CN5_sign => VN_sign_out(7451),
        codeword => codeword(1241),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1242 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7457 downto 7452),
        Din0 => VN1242_in0,
        Din1 => VN1242_in1,
        Din2 => VN1242_in2,
        Din3 => VN1242_in3,
        Din4 => VN1242_in4,
        Din5 => VN1242_in5,
        VN2CN0_bit => VN_data_out(7452),
        VN2CN1_bit => VN_data_out(7453),
        VN2CN2_bit => VN_data_out(7454),
        VN2CN3_bit => VN_data_out(7455),
        VN2CN4_bit => VN_data_out(7456),
        VN2CN5_bit => VN_data_out(7457),
        VN2CN0_sign => VN_sign_out(7452),
        VN2CN1_sign => VN_sign_out(7453),
        VN2CN2_sign => VN_sign_out(7454),
        VN2CN3_sign => VN_sign_out(7455),
        VN2CN4_sign => VN_sign_out(7456),
        VN2CN5_sign => VN_sign_out(7457),
        codeword => codeword(1242),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1243 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7463 downto 7458),
        Din0 => VN1243_in0,
        Din1 => VN1243_in1,
        Din2 => VN1243_in2,
        Din3 => VN1243_in3,
        Din4 => VN1243_in4,
        Din5 => VN1243_in5,
        VN2CN0_bit => VN_data_out(7458),
        VN2CN1_bit => VN_data_out(7459),
        VN2CN2_bit => VN_data_out(7460),
        VN2CN3_bit => VN_data_out(7461),
        VN2CN4_bit => VN_data_out(7462),
        VN2CN5_bit => VN_data_out(7463),
        VN2CN0_sign => VN_sign_out(7458),
        VN2CN1_sign => VN_sign_out(7459),
        VN2CN2_sign => VN_sign_out(7460),
        VN2CN3_sign => VN_sign_out(7461),
        VN2CN4_sign => VN_sign_out(7462),
        VN2CN5_sign => VN_sign_out(7463),
        codeword => codeword(1243),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1244 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7469 downto 7464),
        Din0 => VN1244_in0,
        Din1 => VN1244_in1,
        Din2 => VN1244_in2,
        Din3 => VN1244_in3,
        Din4 => VN1244_in4,
        Din5 => VN1244_in5,
        VN2CN0_bit => VN_data_out(7464),
        VN2CN1_bit => VN_data_out(7465),
        VN2CN2_bit => VN_data_out(7466),
        VN2CN3_bit => VN_data_out(7467),
        VN2CN4_bit => VN_data_out(7468),
        VN2CN5_bit => VN_data_out(7469),
        VN2CN0_sign => VN_sign_out(7464),
        VN2CN1_sign => VN_sign_out(7465),
        VN2CN2_sign => VN_sign_out(7466),
        VN2CN3_sign => VN_sign_out(7467),
        VN2CN4_sign => VN_sign_out(7468),
        VN2CN5_sign => VN_sign_out(7469),
        codeword => codeword(1244),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1245 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7475 downto 7470),
        Din0 => VN1245_in0,
        Din1 => VN1245_in1,
        Din2 => VN1245_in2,
        Din3 => VN1245_in3,
        Din4 => VN1245_in4,
        Din5 => VN1245_in5,
        VN2CN0_bit => VN_data_out(7470),
        VN2CN1_bit => VN_data_out(7471),
        VN2CN2_bit => VN_data_out(7472),
        VN2CN3_bit => VN_data_out(7473),
        VN2CN4_bit => VN_data_out(7474),
        VN2CN5_bit => VN_data_out(7475),
        VN2CN0_sign => VN_sign_out(7470),
        VN2CN1_sign => VN_sign_out(7471),
        VN2CN2_sign => VN_sign_out(7472),
        VN2CN3_sign => VN_sign_out(7473),
        VN2CN4_sign => VN_sign_out(7474),
        VN2CN5_sign => VN_sign_out(7475),
        codeword => codeword(1245),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1246 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7481 downto 7476),
        Din0 => VN1246_in0,
        Din1 => VN1246_in1,
        Din2 => VN1246_in2,
        Din3 => VN1246_in3,
        Din4 => VN1246_in4,
        Din5 => VN1246_in5,
        VN2CN0_bit => VN_data_out(7476),
        VN2CN1_bit => VN_data_out(7477),
        VN2CN2_bit => VN_data_out(7478),
        VN2CN3_bit => VN_data_out(7479),
        VN2CN4_bit => VN_data_out(7480),
        VN2CN5_bit => VN_data_out(7481),
        VN2CN0_sign => VN_sign_out(7476),
        VN2CN1_sign => VN_sign_out(7477),
        VN2CN2_sign => VN_sign_out(7478),
        VN2CN3_sign => VN_sign_out(7479),
        VN2CN4_sign => VN_sign_out(7480),
        VN2CN5_sign => VN_sign_out(7481),
        codeword => codeword(1246),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1247 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7487 downto 7482),
        Din0 => VN1247_in0,
        Din1 => VN1247_in1,
        Din2 => VN1247_in2,
        Din3 => VN1247_in3,
        Din4 => VN1247_in4,
        Din5 => VN1247_in5,
        VN2CN0_bit => VN_data_out(7482),
        VN2CN1_bit => VN_data_out(7483),
        VN2CN2_bit => VN_data_out(7484),
        VN2CN3_bit => VN_data_out(7485),
        VN2CN4_bit => VN_data_out(7486),
        VN2CN5_bit => VN_data_out(7487),
        VN2CN0_sign => VN_sign_out(7482),
        VN2CN1_sign => VN_sign_out(7483),
        VN2CN2_sign => VN_sign_out(7484),
        VN2CN3_sign => VN_sign_out(7485),
        VN2CN4_sign => VN_sign_out(7486),
        VN2CN5_sign => VN_sign_out(7487),
        codeword => codeword(1247),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1248 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7493 downto 7488),
        Din0 => VN1248_in0,
        Din1 => VN1248_in1,
        Din2 => VN1248_in2,
        Din3 => VN1248_in3,
        Din4 => VN1248_in4,
        Din5 => VN1248_in5,
        VN2CN0_bit => VN_data_out(7488),
        VN2CN1_bit => VN_data_out(7489),
        VN2CN2_bit => VN_data_out(7490),
        VN2CN3_bit => VN_data_out(7491),
        VN2CN4_bit => VN_data_out(7492),
        VN2CN5_bit => VN_data_out(7493),
        VN2CN0_sign => VN_sign_out(7488),
        VN2CN1_sign => VN_sign_out(7489),
        VN2CN2_sign => VN_sign_out(7490),
        VN2CN3_sign => VN_sign_out(7491),
        VN2CN4_sign => VN_sign_out(7492),
        VN2CN5_sign => VN_sign_out(7493),
        codeword => codeword(1248),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1249 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7499 downto 7494),
        Din0 => VN1249_in0,
        Din1 => VN1249_in1,
        Din2 => VN1249_in2,
        Din3 => VN1249_in3,
        Din4 => VN1249_in4,
        Din5 => VN1249_in5,
        VN2CN0_bit => VN_data_out(7494),
        VN2CN1_bit => VN_data_out(7495),
        VN2CN2_bit => VN_data_out(7496),
        VN2CN3_bit => VN_data_out(7497),
        VN2CN4_bit => VN_data_out(7498),
        VN2CN5_bit => VN_data_out(7499),
        VN2CN0_sign => VN_sign_out(7494),
        VN2CN1_sign => VN_sign_out(7495),
        VN2CN2_sign => VN_sign_out(7496),
        VN2CN3_sign => VN_sign_out(7497),
        VN2CN4_sign => VN_sign_out(7498),
        VN2CN5_sign => VN_sign_out(7499),
        codeword => codeword(1249),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1250 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7505 downto 7500),
        Din0 => VN1250_in0,
        Din1 => VN1250_in1,
        Din2 => VN1250_in2,
        Din3 => VN1250_in3,
        Din4 => VN1250_in4,
        Din5 => VN1250_in5,
        VN2CN0_bit => VN_data_out(7500),
        VN2CN1_bit => VN_data_out(7501),
        VN2CN2_bit => VN_data_out(7502),
        VN2CN3_bit => VN_data_out(7503),
        VN2CN4_bit => VN_data_out(7504),
        VN2CN5_bit => VN_data_out(7505),
        VN2CN0_sign => VN_sign_out(7500),
        VN2CN1_sign => VN_sign_out(7501),
        VN2CN2_sign => VN_sign_out(7502),
        VN2CN3_sign => VN_sign_out(7503),
        VN2CN4_sign => VN_sign_out(7504),
        VN2CN5_sign => VN_sign_out(7505),
        codeword => codeword(1250),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1251 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7511 downto 7506),
        Din0 => VN1251_in0,
        Din1 => VN1251_in1,
        Din2 => VN1251_in2,
        Din3 => VN1251_in3,
        Din4 => VN1251_in4,
        Din5 => VN1251_in5,
        VN2CN0_bit => VN_data_out(7506),
        VN2CN1_bit => VN_data_out(7507),
        VN2CN2_bit => VN_data_out(7508),
        VN2CN3_bit => VN_data_out(7509),
        VN2CN4_bit => VN_data_out(7510),
        VN2CN5_bit => VN_data_out(7511),
        VN2CN0_sign => VN_sign_out(7506),
        VN2CN1_sign => VN_sign_out(7507),
        VN2CN2_sign => VN_sign_out(7508),
        VN2CN3_sign => VN_sign_out(7509),
        VN2CN4_sign => VN_sign_out(7510),
        VN2CN5_sign => VN_sign_out(7511),
        codeword => codeword(1251),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1252 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7517 downto 7512),
        Din0 => VN1252_in0,
        Din1 => VN1252_in1,
        Din2 => VN1252_in2,
        Din3 => VN1252_in3,
        Din4 => VN1252_in4,
        Din5 => VN1252_in5,
        VN2CN0_bit => VN_data_out(7512),
        VN2CN1_bit => VN_data_out(7513),
        VN2CN2_bit => VN_data_out(7514),
        VN2CN3_bit => VN_data_out(7515),
        VN2CN4_bit => VN_data_out(7516),
        VN2CN5_bit => VN_data_out(7517),
        VN2CN0_sign => VN_sign_out(7512),
        VN2CN1_sign => VN_sign_out(7513),
        VN2CN2_sign => VN_sign_out(7514),
        VN2CN3_sign => VN_sign_out(7515),
        VN2CN4_sign => VN_sign_out(7516),
        VN2CN5_sign => VN_sign_out(7517),
        codeword => codeword(1252),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1253 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7523 downto 7518),
        Din0 => VN1253_in0,
        Din1 => VN1253_in1,
        Din2 => VN1253_in2,
        Din3 => VN1253_in3,
        Din4 => VN1253_in4,
        Din5 => VN1253_in5,
        VN2CN0_bit => VN_data_out(7518),
        VN2CN1_bit => VN_data_out(7519),
        VN2CN2_bit => VN_data_out(7520),
        VN2CN3_bit => VN_data_out(7521),
        VN2CN4_bit => VN_data_out(7522),
        VN2CN5_bit => VN_data_out(7523),
        VN2CN0_sign => VN_sign_out(7518),
        VN2CN1_sign => VN_sign_out(7519),
        VN2CN2_sign => VN_sign_out(7520),
        VN2CN3_sign => VN_sign_out(7521),
        VN2CN4_sign => VN_sign_out(7522),
        VN2CN5_sign => VN_sign_out(7523),
        codeword => codeword(1253),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1254 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7529 downto 7524),
        Din0 => VN1254_in0,
        Din1 => VN1254_in1,
        Din2 => VN1254_in2,
        Din3 => VN1254_in3,
        Din4 => VN1254_in4,
        Din5 => VN1254_in5,
        VN2CN0_bit => VN_data_out(7524),
        VN2CN1_bit => VN_data_out(7525),
        VN2CN2_bit => VN_data_out(7526),
        VN2CN3_bit => VN_data_out(7527),
        VN2CN4_bit => VN_data_out(7528),
        VN2CN5_bit => VN_data_out(7529),
        VN2CN0_sign => VN_sign_out(7524),
        VN2CN1_sign => VN_sign_out(7525),
        VN2CN2_sign => VN_sign_out(7526),
        VN2CN3_sign => VN_sign_out(7527),
        VN2CN4_sign => VN_sign_out(7528),
        VN2CN5_sign => VN_sign_out(7529),
        codeword => codeword(1254),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1255 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7535 downto 7530),
        Din0 => VN1255_in0,
        Din1 => VN1255_in1,
        Din2 => VN1255_in2,
        Din3 => VN1255_in3,
        Din4 => VN1255_in4,
        Din5 => VN1255_in5,
        VN2CN0_bit => VN_data_out(7530),
        VN2CN1_bit => VN_data_out(7531),
        VN2CN2_bit => VN_data_out(7532),
        VN2CN3_bit => VN_data_out(7533),
        VN2CN4_bit => VN_data_out(7534),
        VN2CN5_bit => VN_data_out(7535),
        VN2CN0_sign => VN_sign_out(7530),
        VN2CN1_sign => VN_sign_out(7531),
        VN2CN2_sign => VN_sign_out(7532),
        VN2CN3_sign => VN_sign_out(7533),
        VN2CN4_sign => VN_sign_out(7534),
        VN2CN5_sign => VN_sign_out(7535),
        codeword => codeword(1255),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1256 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7541 downto 7536),
        Din0 => VN1256_in0,
        Din1 => VN1256_in1,
        Din2 => VN1256_in2,
        Din3 => VN1256_in3,
        Din4 => VN1256_in4,
        Din5 => VN1256_in5,
        VN2CN0_bit => VN_data_out(7536),
        VN2CN1_bit => VN_data_out(7537),
        VN2CN2_bit => VN_data_out(7538),
        VN2CN3_bit => VN_data_out(7539),
        VN2CN4_bit => VN_data_out(7540),
        VN2CN5_bit => VN_data_out(7541),
        VN2CN0_sign => VN_sign_out(7536),
        VN2CN1_sign => VN_sign_out(7537),
        VN2CN2_sign => VN_sign_out(7538),
        VN2CN3_sign => VN_sign_out(7539),
        VN2CN4_sign => VN_sign_out(7540),
        VN2CN5_sign => VN_sign_out(7541),
        codeword => codeword(1256),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1257 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7547 downto 7542),
        Din0 => VN1257_in0,
        Din1 => VN1257_in1,
        Din2 => VN1257_in2,
        Din3 => VN1257_in3,
        Din4 => VN1257_in4,
        Din5 => VN1257_in5,
        VN2CN0_bit => VN_data_out(7542),
        VN2CN1_bit => VN_data_out(7543),
        VN2CN2_bit => VN_data_out(7544),
        VN2CN3_bit => VN_data_out(7545),
        VN2CN4_bit => VN_data_out(7546),
        VN2CN5_bit => VN_data_out(7547),
        VN2CN0_sign => VN_sign_out(7542),
        VN2CN1_sign => VN_sign_out(7543),
        VN2CN2_sign => VN_sign_out(7544),
        VN2CN3_sign => VN_sign_out(7545),
        VN2CN4_sign => VN_sign_out(7546),
        VN2CN5_sign => VN_sign_out(7547),
        codeword => codeword(1257),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1258 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7553 downto 7548),
        Din0 => VN1258_in0,
        Din1 => VN1258_in1,
        Din2 => VN1258_in2,
        Din3 => VN1258_in3,
        Din4 => VN1258_in4,
        Din5 => VN1258_in5,
        VN2CN0_bit => VN_data_out(7548),
        VN2CN1_bit => VN_data_out(7549),
        VN2CN2_bit => VN_data_out(7550),
        VN2CN3_bit => VN_data_out(7551),
        VN2CN4_bit => VN_data_out(7552),
        VN2CN5_bit => VN_data_out(7553),
        VN2CN0_sign => VN_sign_out(7548),
        VN2CN1_sign => VN_sign_out(7549),
        VN2CN2_sign => VN_sign_out(7550),
        VN2CN3_sign => VN_sign_out(7551),
        VN2CN4_sign => VN_sign_out(7552),
        VN2CN5_sign => VN_sign_out(7553),
        codeword => codeword(1258),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1259 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7559 downto 7554),
        Din0 => VN1259_in0,
        Din1 => VN1259_in1,
        Din2 => VN1259_in2,
        Din3 => VN1259_in3,
        Din4 => VN1259_in4,
        Din5 => VN1259_in5,
        VN2CN0_bit => VN_data_out(7554),
        VN2CN1_bit => VN_data_out(7555),
        VN2CN2_bit => VN_data_out(7556),
        VN2CN3_bit => VN_data_out(7557),
        VN2CN4_bit => VN_data_out(7558),
        VN2CN5_bit => VN_data_out(7559),
        VN2CN0_sign => VN_sign_out(7554),
        VN2CN1_sign => VN_sign_out(7555),
        VN2CN2_sign => VN_sign_out(7556),
        VN2CN3_sign => VN_sign_out(7557),
        VN2CN4_sign => VN_sign_out(7558),
        VN2CN5_sign => VN_sign_out(7559),
        codeword => codeword(1259),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1260 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7565 downto 7560),
        Din0 => VN1260_in0,
        Din1 => VN1260_in1,
        Din2 => VN1260_in2,
        Din3 => VN1260_in3,
        Din4 => VN1260_in4,
        Din5 => VN1260_in5,
        VN2CN0_bit => VN_data_out(7560),
        VN2CN1_bit => VN_data_out(7561),
        VN2CN2_bit => VN_data_out(7562),
        VN2CN3_bit => VN_data_out(7563),
        VN2CN4_bit => VN_data_out(7564),
        VN2CN5_bit => VN_data_out(7565),
        VN2CN0_sign => VN_sign_out(7560),
        VN2CN1_sign => VN_sign_out(7561),
        VN2CN2_sign => VN_sign_out(7562),
        VN2CN3_sign => VN_sign_out(7563),
        VN2CN4_sign => VN_sign_out(7564),
        VN2CN5_sign => VN_sign_out(7565),
        codeword => codeword(1260),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1261 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7571 downto 7566),
        Din0 => VN1261_in0,
        Din1 => VN1261_in1,
        Din2 => VN1261_in2,
        Din3 => VN1261_in3,
        Din4 => VN1261_in4,
        Din5 => VN1261_in5,
        VN2CN0_bit => VN_data_out(7566),
        VN2CN1_bit => VN_data_out(7567),
        VN2CN2_bit => VN_data_out(7568),
        VN2CN3_bit => VN_data_out(7569),
        VN2CN4_bit => VN_data_out(7570),
        VN2CN5_bit => VN_data_out(7571),
        VN2CN0_sign => VN_sign_out(7566),
        VN2CN1_sign => VN_sign_out(7567),
        VN2CN2_sign => VN_sign_out(7568),
        VN2CN3_sign => VN_sign_out(7569),
        VN2CN4_sign => VN_sign_out(7570),
        VN2CN5_sign => VN_sign_out(7571),
        codeword => codeword(1261),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1262 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7577 downto 7572),
        Din0 => VN1262_in0,
        Din1 => VN1262_in1,
        Din2 => VN1262_in2,
        Din3 => VN1262_in3,
        Din4 => VN1262_in4,
        Din5 => VN1262_in5,
        VN2CN0_bit => VN_data_out(7572),
        VN2CN1_bit => VN_data_out(7573),
        VN2CN2_bit => VN_data_out(7574),
        VN2CN3_bit => VN_data_out(7575),
        VN2CN4_bit => VN_data_out(7576),
        VN2CN5_bit => VN_data_out(7577),
        VN2CN0_sign => VN_sign_out(7572),
        VN2CN1_sign => VN_sign_out(7573),
        VN2CN2_sign => VN_sign_out(7574),
        VN2CN3_sign => VN_sign_out(7575),
        VN2CN4_sign => VN_sign_out(7576),
        VN2CN5_sign => VN_sign_out(7577),
        codeword => codeword(1262),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1263 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7583 downto 7578),
        Din0 => VN1263_in0,
        Din1 => VN1263_in1,
        Din2 => VN1263_in2,
        Din3 => VN1263_in3,
        Din4 => VN1263_in4,
        Din5 => VN1263_in5,
        VN2CN0_bit => VN_data_out(7578),
        VN2CN1_bit => VN_data_out(7579),
        VN2CN2_bit => VN_data_out(7580),
        VN2CN3_bit => VN_data_out(7581),
        VN2CN4_bit => VN_data_out(7582),
        VN2CN5_bit => VN_data_out(7583),
        VN2CN0_sign => VN_sign_out(7578),
        VN2CN1_sign => VN_sign_out(7579),
        VN2CN2_sign => VN_sign_out(7580),
        VN2CN3_sign => VN_sign_out(7581),
        VN2CN4_sign => VN_sign_out(7582),
        VN2CN5_sign => VN_sign_out(7583),
        codeword => codeword(1263),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1264 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7589 downto 7584),
        Din0 => VN1264_in0,
        Din1 => VN1264_in1,
        Din2 => VN1264_in2,
        Din3 => VN1264_in3,
        Din4 => VN1264_in4,
        Din5 => VN1264_in5,
        VN2CN0_bit => VN_data_out(7584),
        VN2CN1_bit => VN_data_out(7585),
        VN2CN2_bit => VN_data_out(7586),
        VN2CN3_bit => VN_data_out(7587),
        VN2CN4_bit => VN_data_out(7588),
        VN2CN5_bit => VN_data_out(7589),
        VN2CN0_sign => VN_sign_out(7584),
        VN2CN1_sign => VN_sign_out(7585),
        VN2CN2_sign => VN_sign_out(7586),
        VN2CN3_sign => VN_sign_out(7587),
        VN2CN4_sign => VN_sign_out(7588),
        VN2CN5_sign => VN_sign_out(7589),
        codeword => codeword(1264),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1265 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7595 downto 7590),
        Din0 => VN1265_in0,
        Din1 => VN1265_in1,
        Din2 => VN1265_in2,
        Din3 => VN1265_in3,
        Din4 => VN1265_in4,
        Din5 => VN1265_in5,
        VN2CN0_bit => VN_data_out(7590),
        VN2CN1_bit => VN_data_out(7591),
        VN2CN2_bit => VN_data_out(7592),
        VN2CN3_bit => VN_data_out(7593),
        VN2CN4_bit => VN_data_out(7594),
        VN2CN5_bit => VN_data_out(7595),
        VN2CN0_sign => VN_sign_out(7590),
        VN2CN1_sign => VN_sign_out(7591),
        VN2CN2_sign => VN_sign_out(7592),
        VN2CN3_sign => VN_sign_out(7593),
        VN2CN4_sign => VN_sign_out(7594),
        VN2CN5_sign => VN_sign_out(7595),
        codeword => codeword(1265),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1266 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7601 downto 7596),
        Din0 => VN1266_in0,
        Din1 => VN1266_in1,
        Din2 => VN1266_in2,
        Din3 => VN1266_in3,
        Din4 => VN1266_in4,
        Din5 => VN1266_in5,
        VN2CN0_bit => VN_data_out(7596),
        VN2CN1_bit => VN_data_out(7597),
        VN2CN2_bit => VN_data_out(7598),
        VN2CN3_bit => VN_data_out(7599),
        VN2CN4_bit => VN_data_out(7600),
        VN2CN5_bit => VN_data_out(7601),
        VN2CN0_sign => VN_sign_out(7596),
        VN2CN1_sign => VN_sign_out(7597),
        VN2CN2_sign => VN_sign_out(7598),
        VN2CN3_sign => VN_sign_out(7599),
        VN2CN4_sign => VN_sign_out(7600),
        VN2CN5_sign => VN_sign_out(7601),
        codeword => codeword(1266),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1267 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7607 downto 7602),
        Din0 => VN1267_in0,
        Din1 => VN1267_in1,
        Din2 => VN1267_in2,
        Din3 => VN1267_in3,
        Din4 => VN1267_in4,
        Din5 => VN1267_in5,
        VN2CN0_bit => VN_data_out(7602),
        VN2CN1_bit => VN_data_out(7603),
        VN2CN2_bit => VN_data_out(7604),
        VN2CN3_bit => VN_data_out(7605),
        VN2CN4_bit => VN_data_out(7606),
        VN2CN5_bit => VN_data_out(7607),
        VN2CN0_sign => VN_sign_out(7602),
        VN2CN1_sign => VN_sign_out(7603),
        VN2CN2_sign => VN_sign_out(7604),
        VN2CN3_sign => VN_sign_out(7605),
        VN2CN4_sign => VN_sign_out(7606),
        VN2CN5_sign => VN_sign_out(7607),
        codeword => codeword(1267),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1268 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7613 downto 7608),
        Din0 => VN1268_in0,
        Din1 => VN1268_in1,
        Din2 => VN1268_in2,
        Din3 => VN1268_in3,
        Din4 => VN1268_in4,
        Din5 => VN1268_in5,
        VN2CN0_bit => VN_data_out(7608),
        VN2CN1_bit => VN_data_out(7609),
        VN2CN2_bit => VN_data_out(7610),
        VN2CN3_bit => VN_data_out(7611),
        VN2CN4_bit => VN_data_out(7612),
        VN2CN5_bit => VN_data_out(7613),
        VN2CN0_sign => VN_sign_out(7608),
        VN2CN1_sign => VN_sign_out(7609),
        VN2CN2_sign => VN_sign_out(7610),
        VN2CN3_sign => VN_sign_out(7611),
        VN2CN4_sign => VN_sign_out(7612),
        VN2CN5_sign => VN_sign_out(7613),
        codeword => codeword(1268),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1269 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7619 downto 7614),
        Din0 => VN1269_in0,
        Din1 => VN1269_in1,
        Din2 => VN1269_in2,
        Din3 => VN1269_in3,
        Din4 => VN1269_in4,
        Din5 => VN1269_in5,
        VN2CN0_bit => VN_data_out(7614),
        VN2CN1_bit => VN_data_out(7615),
        VN2CN2_bit => VN_data_out(7616),
        VN2CN3_bit => VN_data_out(7617),
        VN2CN4_bit => VN_data_out(7618),
        VN2CN5_bit => VN_data_out(7619),
        VN2CN0_sign => VN_sign_out(7614),
        VN2CN1_sign => VN_sign_out(7615),
        VN2CN2_sign => VN_sign_out(7616),
        VN2CN3_sign => VN_sign_out(7617),
        VN2CN4_sign => VN_sign_out(7618),
        VN2CN5_sign => VN_sign_out(7619),
        codeword => codeword(1269),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1270 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7625 downto 7620),
        Din0 => VN1270_in0,
        Din1 => VN1270_in1,
        Din2 => VN1270_in2,
        Din3 => VN1270_in3,
        Din4 => VN1270_in4,
        Din5 => VN1270_in5,
        VN2CN0_bit => VN_data_out(7620),
        VN2CN1_bit => VN_data_out(7621),
        VN2CN2_bit => VN_data_out(7622),
        VN2CN3_bit => VN_data_out(7623),
        VN2CN4_bit => VN_data_out(7624),
        VN2CN5_bit => VN_data_out(7625),
        VN2CN0_sign => VN_sign_out(7620),
        VN2CN1_sign => VN_sign_out(7621),
        VN2CN2_sign => VN_sign_out(7622),
        VN2CN3_sign => VN_sign_out(7623),
        VN2CN4_sign => VN_sign_out(7624),
        VN2CN5_sign => VN_sign_out(7625),
        codeword => codeword(1270),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1271 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7631 downto 7626),
        Din0 => VN1271_in0,
        Din1 => VN1271_in1,
        Din2 => VN1271_in2,
        Din3 => VN1271_in3,
        Din4 => VN1271_in4,
        Din5 => VN1271_in5,
        VN2CN0_bit => VN_data_out(7626),
        VN2CN1_bit => VN_data_out(7627),
        VN2CN2_bit => VN_data_out(7628),
        VN2CN3_bit => VN_data_out(7629),
        VN2CN4_bit => VN_data_out(7630),
        VN2CN5_bit => VN_data_out(7631),
        VN2CN0_sign => VN_sign_out(7626),
        VN2CN1_sign => VN_sign_out(7627),
        VN2CN2_sign => VN_sign_out(7628),
        VN2CN3_sign => VN_sign_out(7629),
        VN2CN4_sign => VN_sign_out(7630),
        VN2CN5_sign => VN_sign_out(7631),
        codeword => codeword(1271),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1272 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7637 downto 7632),
        Din0 => VN1272_in0,
        Din1 => VN1272_in1,
        Din2 => VN1272_in2,
        Din3 => VN1272_in3,
        Din4 => VN1272_in4,
        Din5 => VN1272_in5,
        VN2CN0_bit => VN_data_out(7632),
        VN2CN1_bit => VN_data_out(7633),
        VN2CN2_bit => VN_data_out(7634),
        VN2CN3_bit => VN_data_out(7635),
        VN2CN4_bit => VN_data_out(7636),
        VN2CN5_bit => VN_data_out(7637),
        VN2CN0_sign => VN_sign_out(7632),
        VN2CN1_sign => VN_sign_out(7633),
        VN2CN2_sign => VN_sign_out(7634),
        VN2CN3_sign => VN_sign_out(7635),
        VN2CN4_sign => VN_sign_out(7636),
        VN2CN5_sign => VN_sign_out(7637),
        codeword => codeword(1272),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1273 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7643 downto 7638),
        Din0 => VN1273_in0,
        Din1 => VN1273_in1,
        Din2 => VN1273_in2,
        Din3 => VN1273_in3,
        Din4 => VN1273_in4,
        Din5 => VN1273_in5,
        VN2CN0_bit => VN_data_out(7638),
        VN2CN1_bit => VN_data_out(7639),
        VN2CN2_bit => VN_data_out(7640),
        VN2CN3_bit => VN_data_out(7641),
        VN2CN4_bit => VN_data_out(7642),
        VN2CN5_bit => VN_data_out(7643),
        VN2CN0_sign => VN_sign_out(7638),
        VN2CN1_sign => VN_sign_out(7639),
        VN2CN2_sign => VN_sign_out(7640),
        VN2CN3_sign => VN_sign_out(7641),
        VN2CN4_sign => VN_sign_out(7642),
        VN2CN5_sign => VN_sign_out(7643),
        codeword => codeword(1273),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1274 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7649 downto 7644),
        Din0 => VN1274_in0,
        Din1 => VN1274_in1,
        Din2 => VN1274_in2,
        Din3 => VN1274_in3,
        Din4 => VN1274_in4,
        Din5 => VN1274_in5,
        VN2CN0_bit => VN_data_out(7644),
        VN2CN1_bit => VN_data_out(7645),
        VN2CN2_bit => VN_data_out(7646),
        VN2CN3_bit => VN_data_out(7647),
        VN2CN4_bit => VN_data_out(7648),
        VN2CN5_bit => VN_data_out(7649),
        VN2CN0_sign => VN_sign_out(7644),
        VN2CN1_sign => VN_sign_out(7645),
        VN2CN2_sign => VN_sign_out(7646),
        VN2CN3_sign => VN_sign_out(7647),
        VN2CN4_sign => VN_sign_out(7648),
        VN2CN5_sign => VN_sign_out(7649),
        codeword => codeword(1274),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1275 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7655 downto 7650),
        Din0 => VN1275_in0,
        Din1 => VN1275_in1,
        Din2 => VN1275_in2,
        Din3 => VN1275_in3,
        Din4 => VN1275_in4,
        Din5 => VN1275_in5,
        VN2CN0_bit => VN_data_out(7650),
        VN2CN1_bit => VN_data_out(7651),
        VN2CN2_bit => VN_data_out(7652),
        VN2CN3_bit => VN_data_out(7653),
        VN2CN4_bit => VN_data_out(7654),
        VN2CN5_bit => VN_data_out(7655),
        VN2CN0_sign => VN_sign_out(7650),
        VN2CN1_sign => VN_sign_out(7651),
        VN2CN2_sign => VN_sign_out(7652),
        VN2CN3_sign => VN_sign_out(7653),
        VN2CN4_sign => VN_sign_out(7654),
        VN2CN5_sign => VN_sign_out(7655),
        codeword => codeword(1275),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1276 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7661 downto 7656),
        Din0 => VN1276_in0,
        Din1 => VN1276_in1,
        Din2 => VN1276_in2,
        Din3 => VN1276_in3,
        Din4 => VN1276_in4,
        Din5 => VN1276_in5,
        VN2CN0_bit => VN_data_out(7656),
        VN2CN1_bit => VN_data_out(7657),
        VN2CN2_bit => VN_data_out(7658),
        VN2CN3_bit => VN_data_out(7659),
        VN2CN4_bit => VN_data_out(7660),
        VN2CN5_bit => VN_data_out(7661),
        VN2CN0_sign => VN_sign_out(7656),
        VN2CN1_sign => VN_sign_out(7657),
        VN2CN2_sign => VN_sign_out(7658),
        VN2CN3_sign => VN_sign_out(7659),
        VN2CN4_sign => VN_sign_out(7660),
        VN2CN5_sign => VN_sign_out(7661),
        codeword => codeword(1276),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1277 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7667 downto 7662),
        Din0 => VN1277_in0,
        Din1 => VN1277_in1,
        Din2 => VN1277_in2,
        Din3 => VN1277_in3,
        Din4 => VN1277_in4,
        Din5 => VN1277_in5,
        VN2CN0_bit => VN_data_out(7662),
        VN2CN1_bit => VN_data_out(7663),
        VN2CN2_bit => VN_data_out(7664),
        VN2CN3_bit => VN_data_out(7665),
        VN2CN4_bit => VN_data_out(7666),
        VN2CN5_bit => VN_data_out(7667),
        VN2CN0_sign => VN_sign_out(7662),
        VN2CN1_sign => VN_sign_out(7663),
        VN2CN2_sign => VN_sign_out(7664),
        VN2CN3_sign => VN_sign_out(7665),
        VN2CN4_sign => VN_sign_out(7666),
        VN2CN5_sign => VN_sign_out(7667),
        codeword => codeword(1277),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1278 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7673 downto 7668),
        Din0 => VN1278_in0,
        Din1 => VN1278_in1,
        Din2 => VN1278_in2,
        Din3 => VN1278_in3,
        Din4 => VN1278_in4,
        Din5 => VN1278_in5,
        VN2CN0_bit => VN_data_out(7668),
        VN2CN1_bit => VN_data_out(7669),
        VN2CN2_bit => VN_data_out(7670),
        VN2CN3_bit => VN_data_out(7671),
        VN2CN4_bit => VN_data_out(7672),
        VN2CN5_bit => VN_data_out(7673),
        VN2CN0_sign => VN_sign_out(7668),
        VN2CN1_sign => VN_sign_out(7669),
        VN2CN2_sign => VN_sign_out(7670),
        VN2CN3_sign => VN_sign_out(7671),
        VN2CN4_sign => VN_sign_out(7672),
        VN2CN5_sign => VN_sign_out(7673),
        codeword => codeword(1278),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1279 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7679 downto 7674),
        Din0 => VN1279_in0,
        Din1 => VN1279_in1,
        Din2 => VN1279_in2,
        Din3 => VN1279_in3,
        Din4 => VN1279_in4,
        Din5 => VN1279_in5,
        VN2CN0_bit => VN_data_out(7674),
        VN2CN1_bit => VN_data_out(7675),
        VN2CN2_bit => VN_data_out(7676),
        VN2CN3_bit => VN_data_out(7677),
        VN2CN4_bit => VN_data_out(7678),
        VN2CN5_bit => VN_data_out(7679),
        VN2CN0_sign => VN_sign_out(7674),
        VN2CN1_sign => VN_sign_out(7675),
        VN2CN2_sign => VN_sign_out(7676),
        VN2CN3_sign => VN_sign_out(7677),
        VN2CN4_sign => VN_sign_out(7678),
        VN2CN5_sign => VN_sign_out(7679),
        codeword => codeword(1279),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1280 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7685 downto 7680),
        Din0 => VN1280_in0,
        Din1 => VN1280_in1,
        Din2 => VN1280_in2,
        Din3 => VN1280_in3,
        Din4 => VN1280_in4,
        Din5 => VN1280_in5,
        VN2CN0_bit => VN_data_out(7680),
        VN2CN1_bit => VN_data_out(7681),
        VN2CN2_bit => VN_data_out(7682),
        VN2CN3_bit => VN_data_out(7683),
        VN2CN4_bit => VN_data_out(7684),
        VN2CN5_bit => VN_data_out(7685),
        VN2CN0_sign => VN_sign_out(7680),
        VN2CN1_sign => VN_sign_out(7681),
        VN2CN2_sign => VN_sign_out(7682),
        VN2CN3_sign => VN_sign_out(7683),
        VN2CN4_sign => VN_sign_out(7684),
        VN2CN5_sign => VN_sign_out(7685),
        codeword => codeword(1280),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1281 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7691 downto 7686),
        Din0 => VN1281_in0,
        Din1 => VN1281_in1,
        Din2 => VN1281_in2,
        Din3 => VN1281_in3,
        Din4 => VN1281_in4,
        Din5 => VN1281_in5,
        VN2CN0_bit => VN_data_out(7686),
        VN2CN1_bit => VN_data_out(7687),
        VN2CN2_bit => VN_data_out(7688),
        VN2CN3_bit => VN_data_out(7689),
        VN2CN4_bit => VN_data_out(7690),
        VN2CN5_bit => VN_data_out(7691),
        VN2CN0_sign => VN_sign_out(7686),
        VN2CN1_sign => VN_sign_out(7687),
        VN2CN2_sign => VN_sign_out(7688),
        VN2CN3_sign => VN_sign_out(7689),
        VN2CN4_sign => VN_sign_out(7690),
        VN2CN5_sign => VN_sign_out(7691),
        codeword => codeword(1281),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1282 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7697 downto 7692),
        Din0 => VN1282_in0,
        Din1 => VN1282_in1,
        Din2 => VN1282_in2,
        Din3 => VN1282_in3,
        Din4 => VN1282_in4,
        Din5 => VN1282_in5,
        VN2CN0_bit => VN_data_out(7692),
        VN2CN1_bit => VN_data_out(7693),
        VN2CN2_bit => VN_data_out(7694),
        VN2CN3_bit => VN_data_out(7695),
        VN2CN4_bit => VN_data_out(7696),
        VN2CN5_bit => VN_data_out(7697),
        VN2CN0_sign => VN_sign_out(7692),
        VN2CN1_sign => VN_sign_out(7693),
        VN2CN2_sign => VN_sign_out(7694),
        VN2CN3_sign => VN_sign_out(7695),
        VN2CN4_sign => VN_sign_out(7696),
        VN2CN5_sign => VN_sign_out(7697),
        codeword => codeword(1282),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1283 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7703 downto 7698),
        Din0 => VN1283_in0,
        Din1 => VN1283_in1,
        Din2 => VN1283_in2,
        Din3 => VN1283_in3,
        Din4 => VN1283_in4,
        Din5 => VN1283_in5,
        VN2CN0_bit => VN_data_out(7698),
        VN2CN1_bit => VN_data_out(7699),
        VN2CN2_bit => VN_data_out(7700),
        VN2CN3_bit => VN_data_out(7701),
        VN2CN4_bit => VN_data_out(7702),
        VN2CN5_bit => VN_data_out(7703),
        VN2CN0_sign => VN_sign_out(7698),
        VN2CN1_sign => VN_sign_out(7699),
        VN2CN2_sign => VN_sign_out(7700),
        VN2CN3_sign => VN_sign_out(7701),
        VN2CN4_sign => VN_sign_out(7702),
        VN2CN5_sign => VN_sign_out(7703),
        codeword => codeword(1283),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1284 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7709 downto 7704),
        Din0 => VN1284_in0,
        Din1 => VN1284_in1,
        Din2 => VN1284_in2,
        Din3 => VN1284_in3,
        Din4 => VN1284_in4,
        Din5 => VN1284_in5,
        VN2CN0_bit => VN_data_out(7704),
        VN2CN1_bit => VN_data_out(7705),
        VN2CN2_bit => VN_data_out(7706),
        VN2CN3_bit => VN_data_out(7707),
        VN2CN4_bit => VN_data_out(7708),
        VN2CN5_bit => VN_data_out(7709),
        VN2CN0_sign => VN_sign_out(7704),
        VN2CN1_sign => VN_sign_out(7705),
        VN2CN2_sign => VN_sign_out(7706),
        VN2CN3_sign => VN_sign_out(7707),
        VN2CN4_sign => VN_sign_out(7708),
        VN2CN5_sign => VN_sign_out(7709),
        codeword => codeword(1284),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1285 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7715 downto 7710),
        Din0 => VN1285_in0,
        Din1 => VN1285_in1,
        Din2 => VN1285_in2,
        Din3 => VN1285_in3,
        Din4 => VN1285_in4,
        Din5 => VN1285_in5,
        VN2CN0_bit => VN_data_out(7710),
        VN2CN1_bit => VN_data_out(7711),
        VN2CN2_bit => VN_data_out(7712),
        VN2CN3_bit => VN_data_out(7713),
        VN2CN4_bit => VN_data_out(7714),
        VN2CN5_bit => VN_data_out(7715),
        VN2CN0_sign => VN_sign_out(7710),
        VN2CN1_sign => VN_sign_out(7711),
        VN2CN2_sign => VN_sign_out(7712),
        VN2CN3_sign => VN_sign_out(7713),
        VN2CN4_sign => VN_sign_out(7714),
        VN2CN5_sign => VN_sign_out(7715),
        codeword => codeword(1285),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1286 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7721 downto 7716),
        Din0 => VN1286_in0,
        Din1 => VN1286_in1,
        Din2 => VN1286_in2,
        Din3 => VN1286_in3,
        Din4 => VN1286_in4,
        Din5 => VN1286_in5,
        VN2CN0_bit => VN_data_out(7716),
        VN2CN1_bit => VN_data_out(7717),
        VN2CN2_bit => VN_data_out(7718),
        VN2CN3_bit => VN_data_out(7719),
        VN2CN4_bit => VN_data_out(7720),
        VN2CN5_bit => VN_data_out(7721),
        VN2CN0_sign => VN_sign_out(7716),
        VN2CN1_sign => VN_sign_out(7717),
        VN2CN2_sign => VN_sign_out(7718),
        VN2CN3_sign => VN_sign_out(7719),
        VN2CN4_sign => VN_sign_out(7720),
        VN2CN5_sign => VN_sign_out(7721),
        codeword => codeword(1286),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1287 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7727 downto 7722),
        Din0 => VN1287_in0,
        Din1 => VN1287_in1,
        Din2 => VN1287_in2,
        Din3 => VN1287_in3,
        Din4 => VN1287_in4,
        Din5 => VN1287_in5,
        VN2CN0_bit => VN_data_out(7722),
        VN2CN1_bit => VN_data_out(7723),
        VN2CN2_bit => VN_data_out(7724),
        VN2CN3_bit => VN_data_out(7725),
        VN2CN4_bit => VN_data_out(7726),
        VN2CN5_bit => VN_data_out(7727),
        VN2CN0_sign => VN_sign_out(7722),
        VN2CN1_sign => VN_sign_out(7723),
        VN2CN2_sign => VN_sign_out(7724),
        VN2CN3_sign => VN_sign_out(7725),
        VN2CN4_sign => VN_sign_out(7726),
        VN2CN5_sign => VN_sign_out(7727),
        codeword => codeword(1287),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1288 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7733 downto 7728),
        Din0 => VN1288_in0,
        Din1 => VN1288_in1,
        Din2 => VN1288_in2,
        Din3 => VN1288_in3,
        Din4 => VN1288_in4,
        Din5 => VN1288_in5,
        VN2CN0_bit => VN_data_out(7728),
        VN2CN1_bit => VN_data_out(7729),
        VN2CN2_bit => VN_data_out(7730),
        VN2CN3_bit => VN_data_out(7731),
        VN2CN4_bit => VN_data_out(7732),
        VN2CN5_bit => VN_data_out(7733),
        VN2CN0_sign => VN_sign_out(7728),
        VN2CN1_sign => VN_sign_out(7729),
        VN2CN2_sign => VN_sign_out(7730),
        VN2CN3_sign => VN_sign_out(7731),
        VN2CN4_sign => VN_sign_out(7732),
        VN2CN5_sign => VN_sign_out(7733),
        codeword => codeword(1288),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1289 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7739 downto 7734),
        Din0 => VN1289_in0,
        Din1 => VN1289_in1,
        Din2 => VN1289_in2,
        Din3 => VN1289_in3,
        Din4 => VN1289_in4,
        Din5 => VN1289_in5,
        VN2CN0_bit => VN_data_out(7734),
        VN2CN1_bit => VN_data_out(7735),
        VN2CN2_bit => VN_data_out(7736),
        VN2CN3_bit => VN_data_out(7737),
        VN2CN4_bit => VN_data_out(7738),
        VN2CN5_bit => VN_data_out(7739),
        VN2CN0_sign => VN_sign_out(7734),
        VN2CN1_sign => VN_sign_out(7735),
        VN2CN2_sign => VN_sign_out(7736),
        VN2CN3_sign => VN_sign_out(7737),
        VN2CN4_sign => VN_sign_out(7738),
        VN2CN5_sign => VN_sign_out(7739),
        codeword => codeword(1289),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1290 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7745 downto 7740),
        Din0 => VN1290_in0,
        Din1 => VN1290_in1,
        Din2 => VN1290_in2,
        Din3 => VN1290_in3,
        Din4 => VN1290_in4,
        Din5 => VN1290_in5,
        VN2CN0_bit => VN_data_out(7740),
        VN2CN1_bit => VN_data_out(7741),
        VN2CN2_bit => VN_data_out(7742),
        VN2CN3_bit => VN_data_out(7743),
        VN2CN4_bit => VN_data_out(7744),
        VN2CN5_bit => VN_data_out(7745),
        VN2CN0_sign => VN_sign_out(7740),
        VN2CN1_sign => VN_sign_out(7741),
        VN2CN2_sign => VN_sign_out(7742),
        VN2CN3_sign => VN_sign_out(7743),
        VN2CN4_sign => VN_sign_out(7744),
        VN2CN5_sign => VN_sign_out(7745),
        codeword => codeword(1290),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1291 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7751 downto 7746),
        Din0 => VN1291_in0,
        Din1 => VN1291_in1,
        Din2 => VN1291_in2,
        Din3 => VN1291_in3,
        Din4 => VN1291_in4,
        Din5 => VN1291_in5,
        VN2CN0_bit => VN_data_out(7746),
        VN2CN1_bit => VN_data_out(7747),
        VN2CN2_bit => VN_data_out(7748),
        VN2CN3_bit => VN_data_out(7749),
        VN2CN4_bit => VN_data_out(7750),
        VN2CN5_bit => VN_data_out(7751),
        VN2CN0_sign => VN_sign_out(7746),
        VN2CN1_sign => VN_sign_out(7747),
        VN2CN2_sign => VN_sign_out(7748),
        VN2CN3_sign => VN_sign_out(7749),
        VN2CN4_sign => VN_sign_out(7750),
        VN2CN5_sign => VN_sign_out(7751),
        codeword => codeword(1291),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1292 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7757 downto 7752),
        Din0 => VN1292_in0,
        Din1 => VN1292_in1,
        Din2 => VN1292_in2,
        Din3 => VN1292_in3,
        Din4 => VN1292_in4,
        Din5 => VN1292_in5,
        VN2CN0_bit => VN_data_out(7752),
        VN2CN1_bit => VN_data_out(7753),
        VN2CN2_bit => VN_data_out(7754),
        VN2CN3_bit => VN_data_out(7755),
        VN2CN4_bit => VN_data_out(7756),
        VN2CN5_bit => VN_data_out(7757),
        VN2CN0_sign => VN_sign_out(7752),
        VN2CN1_sign => VN_sign_out(7753),
        VN2CN2_sign => VN_sign_out(7754),
        VN2CN3_sign => VN_sign_out(7755),
        VN2CN4_sign => VN_sign_out(7756),
        VN2CN5_sign => VN_sign_out(7757),
        codeword => codeword(1292),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1293 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7763 downto 7758),
        Din0 => VN1293_in0,
        Din1 => VN1293_in1,
        Din2 => VN1293_in2,
        Din3 => VN1293_in3,
        Din4 => VN1293_in4,
        Din5 => VN1293_in5,
        VN2CN0_bit => VN_data_out(7758),
        VN2CN1_bit => VN_data_out(7759),
        VN2CN2_bit => VN_data_out(7760),
        VN2CN3_bit => VN_data_out(7761),
        VN2CN4_bit => VN_data_out(7762),
        VN2CN5_bit => VN_data_out(7763),
        VN2CN0_sign => VN_sign_out(7758),
        VN2CN1_sign => VN_sign_out(7759),
        VN2CN2_sign => VN_sign_out(7760),
        VN2CN3_sign => VN_sign_out(7761),
        VN2CN4_sign => VN_sign_out(7762),
        VN2CN5_sign => VN_sign_out(7763),
        codeword => codeword(1293),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1294 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7769 downto 7764),
        Din0 => VN1294_in0,
        Din1 => VN1294_in1,
        Din2 => VN1294_in2,
        Din3 => VN1294_in3,
        Din4 => VN1294_in4,
        Din5 => VN1294_in5,
        VN2CN0_bit => VN_data_out(7764),
        VN2CN1_bit => VN_data_out(7765),
        VN2CN2_bit => VN_data_out(7766),
        VN2CN3_bit => VN_data_out(7767),
        VN2CN4_bit => VN_data_out(7768),
        VN2CN5_bit => VN_data_out(7769),
        VN2CN0_sign => VN_sign_out(7764),
        VN2CN1_sign => VN_sign_out(7765),
        VN2CN2_sign => VN_sign_out(7766),
        VN2CN3_sign => VN_sign_out(7767),
        VN2CN4_sign => VN_sign_out(7768),
        VN2CN5_sign => VN_sign_out(7769),
        codeword => codeword(1294),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1295 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7775 downto 7770),
        Din0 => VN1295_in0,
        Din1 => VN1295_in1,
        Din2 => VN1295_in2,
        Din3 => VN1295_in3,
        Din4 => VN1295_in4,
        Din5 => VN1295_in5,
        VN2CN0_bit => VN_data_out(7770),
        VN2CN1_bit => VN_data_out(7771),
        VN2CN2_bit => VN_data_out(7772),
        VN2CN3_bit => VN_data_out(7773),
        VN2CN4_bit => VN_data_out(7774),
        VN2CN5_bit => VN_data_out(7775),
        VN2CN0_sign => VN_sign_out(7770),
        VN2CN1_sign => VN_sign_out(7771),
        VN2CN2_sign => VN_sign_out(7772),
        VN2CN3_sign => VN_sign_out(7773),
        VN2CN4_sign => VN_sign_out(7774),
        VN2CN5_sign => VN_sign_out(7775),
        codeword => codeword(1295),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1296 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7781 downto 7776),
        Din0 => VN1296_in0,
        Din1 => VN1296_in1,
        Din2 => VN1296_in2,
        Din3 => VN1296_in3,
        Din4 => VN1296_in4,
        Din5 => VN1296_in5,
        VN2CN0_bit => VN_data_out(7776),
        VN2CN1_bit => VN_data_out(7777),
        VN2CN2_bit => VN_data_out(7778),
        VN2CN3_bit => VN_data_out(7779),
        VN2CN4_bit => VN_data_out(7780),
        VN2CN5_bit => VN_data_out(7781),
        VN2CN0_sign => VN_sign_out(7776),
        VN2CN1_sign => VN_sign_out(7777),
        VN2CN2_sign => VN_sign_out(7778),
        VN2CN3_sign => VN_sign_out(7779),
        VN2CN4_sign => VN_sign_out(7780),
        VN2CN5_sign => VN_sign_out(7781),
        codeword => codeword(1296),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1297 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7787 downto 7782),
        Din0 => VN1297_in0,
        Din1 => VN1297_in1,
        Din2 => VN1297_in2,
        Din3 => VN1297_in3,
        Din4 => VN1297_in4,
        Din5 => VN1297_in5,
        VN2CN0_bit => VN_data_out(7782),
        VN2CN1_bit => VN_data_out(7783),
        VN2CN2_bit => VN_data_out(7784),
        VN2CN3_bit => VN_data_out(7785),
        VN2CN4_bit => VN_data_out(7786),
        VN2CN5_bit => VN_data_out(7787),
        VN2CN0_sign => VN_sign_out(7782),
        VN2CN1_sign => VN_sign_out(7783),
        VN2CN2_sign => VN_sign_out(7784),
        VN2CN3_sign => VN_sign_out(7785),
        VN2CN4_sign => VN_sign_out(7786),
        VN2CN5_sign => VN_sign_out(7787),
        codeword => codeword(1297),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1298 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7793 downto 7788),
        Din0 => VN1298_in0,
        Din1 => VN1298_in1,
        Din2 => VN1298_in2,
        Din3 => VN1298_in3,
        Din4 => VN1298_in4,
        Din5 => VN1298_in5,
        VN2CN0_bit => VN_data_out(7788),
        VN2CN1_bit => VN_data_out(7789),
        VN2CN2_bit => VN_data_out(7790),
        VN2CN3_bit => VN_data_out(7791),
        VN2CN4_bit => VN_data_out(7792),
        VN2CN5_bit => VN_data_out(7793),
        VN2CN0_sign => VN_sign_out(7788),
        VN2CN1_sign => VN_sign_out(7789),
        VN2CN2_sign => VN_sign_out(7790),
        VN2CN3_sign => VN_sign_out(7791),
        VN2CN4_sign => VN_sign_out(7792),
        VN2CN5_sign => VN_sign_out(7793),
        codeword => codeword(1298),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1299 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7799 downto 7794),
        Din0 => VN1299_in0,
        Din1 => VN1299_in1,
        Din2 => VN1299_in2,
        Din3 => VN1299_in3,
        Din4 => VN1299_in4,
        Din5 => VN1299_in5,
        VN2CN0_bit => VN_data_out(7794),
        VN2CN1_bit => VN_data_out(7795),
        VN2CN2_bit => VN_data_out(7796),
        VN2CN3_bit => VN_data_out(7797),
        VN2CN4_bit => VN_data_out(7798),
        VN2CN5_bit => VN_data_out(7799),
        VN2CN0_sign => VN_sign_out(7794),
        VN2CN1_sign => VN_sign_out(7795),
        VN2CN2_sign => VN_sign_out(7796),
        VN2CN3_sign => VN_sign_out(7797),
        VN2CN4_sign => VN_sign_out(7798),
        VN2CN5_sign => VN_sign_out(7799),
        codeword => codeword(1299),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1300 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7805 downto 7800),
        Din0 => VN1300_in0,
        Din1 => VN1300_in1,
        Din2 => VN1300_in2,
        Din3 => VN1300_in3,
        Din4 => VN1300_in4,
        Din5 => VN1300_in5,
        VN2CN0_bit => VN_data_out(7800),
        VN2CN1_bit => VN_data_out(7801),
        VN2CN2_bit => VN_data_out(7802),
        VN2CN3_bit => VN_data_out(7803),
        VN2CN4_bit => VN_data_out(7804),
        VN2CN5_bit => VN_data_out(7805),
        VN2CN0_sign => VN_sign_out(7800),
        VN2CN1_sign => VN_sign_out(7801),
        VN2CN2_sign => VN_sign_out(7802),
        VN2CN3_sign => VN_sign_out(7803),
        VN2CN4_sign => VN_sign_out(7804),
        VN2CN5_sign => VN_sign_out(7805),
        codeword => codeword(1300),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1301 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7811 downto 7806),
        Din0 => VN1301_in0,
        Din1 => VN1301_in1,
        Din2 => VN1301_in2,
        Din3 => VN1301_in3,
        Din4 => VN1301_in4,
        Din5 => VN1301_in5,
        VN2CN0_bit => VN_data_out(7806),
        VN2CN1_bit => VN_data_out(7807),
        VN2CN2_bit => VN_data_out(7808),
        VN2CN3_bit => VN_data_out(7809),
        VN2CN4_bit => VN_data_out(7810),
        VN2CN5_bit => VN_data_out(7811),
        VN2CN0_sign => VN_sign_out(7806),
        VN2CN1_sign => VN_sign_out(7807),
        VN2CN2_sign => VN_sign_out(7808),
        VN2CN3_sign => VN_sign_out(7809),
        VN2CN4_sign => VN_sign_out(7810),
        VN2CN5_sign => VN_sign_out(7811),
        codeword => codeword(1301),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1302 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7817 downto 7812),
        Din0 => VN1302_in0,
        Din1 => VN1302_in1,
        Din2 => VN1302_in2,
        Din3 => VN1302_in3,
        Din4 => VN1302_in4,
        Din5 => VN1302_in5,
        VN2CN0_bit => VN_data_out(7812),
        VN2CN1_bit => VN_data_out(7813),
        VN2CN2_bit => VN_data_out(7814),
        VN2CN3_bit => VN_data_out(7815),
        VN2CN4_bit => VN_data_out(7816),
        VN2CN5_bit => VN_data_out(7817),
        VN2CN0_sign => VN_sign_out(7812),
        VN2CN1_sign => VN_sign_out(7813),
        VN2CN2_sign => VN_sign_out(7814),
        VN2CN3_sign => VN_sign_out(7815),
        VN2CN4_sign => VN_sign_out(7816),
        VN2CN5_sign => VN_sign_out(7817),
        codeword => codeword(1302),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1303 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7823 downto 7818),
        Din0 => VN1303_in0,
        Din1 => VN1303_in1,
        Din2 => VN1303_in2,
        Din3 => VN1303_in3,
        Din4 => VN1303_in4,
        Din5 => VN1303_in5,
        VN2CN0_bit => VN_data_out(7818),
        VN2CN1_bit => VN_data_out(7819),
        VN2CN2_bit => VN_data_out(7820),
        VN2CN3_bit => VN_data_out(7821),
        VN2CN4_bit => VN_data_out(7822),
        VN2CN5_bit => VN_data_out(7823),
        VN2CN0_sign => VN_sign_out(7818),
        VN2CN1_sign => VN_sign_out(7819),
        VN2CN2_sign => VN_sign_out(7820),
        VN2CN3_sign => VN_sign_out(7821),
        VN2CN4_sign => VN_sign_out(7822),
        VN2CN5_sign => VN_sign_out(7823),
        codeword => codeword(1303),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1304 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7829 downto 7824),
        Din0 => VN1304_in0,
        Din1 => VN1304_in1,
        Din2 => VN1304_in2,
        Din3 => VN1304_in3,
        Din4 => VN1304_in4,
        Din5 => VN1304_in5,
        VN2CN0_bit => VN_data_out(7824),
        VN2CN1_bit => VN_data_out(7825),
        VN2CN2_bit => VN_data_out(7826),
        VN2CN3_bit => VN_data_out(7827),
        VN2CN4_bit => VN_data_out(7828),
        VN2CN5_bit => VN_data_out(7829),
        VN2CN0_sign => VN_sign_out(7824),
        VN2CN1_sign => VN_sign_out(7825),
        VN2CN2_sign => VN_sign_out(7826),
        VN2CN3_sign => VN_sign_out(7827),
        VN2CN4_sign => VN_sign_out(7828),
        VN2CN5_sign => VN_sign_out(7829),
        codeword => codeword(1304),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1305 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7835 downto 7830),
        Din0 => VN1305_in0,
        Din1 => VN1305_in1,
        Din2 => VN1305_in2,
        Din3 => VN1305_in3,
        Din4 => VN1305_in4,
        Din5 => VN1305_in5,
        VN2CN0_bit => VN_data_out(7830),
        VN2CN1_bit => VN_data_out(7831),
        VN2CN2_bit => VN_data_out(7832),
        VN2CN3_bit => VN_data_out(7833),
        VN2CN4_bit => VN_data_out(7834),
        VN2CN5_bit => VN_data_out(7835),
        VN2CN0_sign => VN_sign_out(7830),
        VN2CN1_sign => VN_sign_out(7831),
        VN2CN2_sign => VN_sign_out(7832),
        VN2CN3_sign => VN_sign_out(7833),
        VN2CN4_sign => VN_sign_out(7834),
        VN2CN5_sign => VN_sign_out(7835),
        codeword => codeword(1305),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1306 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7841 downto 7836),
        Din0 => VN1306_in0,
        Din1 => VN1306_in1,
        Din2 => VN1306_in2,
        Din3 => VN1306_in3,
        Din4 => VN1306_in4,
        Din5 => VN1306_in5,
        VN2CN0_bit => VN_data_out(7836),
        VN2CN1_bit => VN_data_out(7837),
        VN2CN2_bit => VN_data_out(7838),
        VN2CN3_bit => VN_data_out(7839),
        VN2CN4_bit => VN_data_out(7840),
        VN2CN5_bit => VN_data_out(7841),
        VN2CN0_sign => VN_sign_out(7836),
        VN2CN1_sign => VN_sign_out(7837),
        VN2CN2_sign => VN_sign_out(7838),
        VN2CN3_sign => VN_sign_out(7839),
        VN2CN4_sign => VN_sign_out(7840),
        VN2CN5_sign => VN_sign_out(7841),
        codeword => codeword(1306),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1307 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7847 downto 7842),
        Din0 => VN1307_in0,
        Din1 => VN1307_in1,
        Din2 => VN1307_in2,
        Din3 => VN1307_in3,
        Din4 => VN1307_in4,
        Din5 => VN1307_in5,
        VN2CN0_bit => VN_data_out(7842),
        VN2CN1_bit => VN_data_out(7843),
        VN2CN2_bit => VN_data_out(7844),
        VN2CN3_bit => VN_data_out(7845),
        VN2CN4_bit => VN_data_out(7846),
        VN2CN5_bit => VN_data_out(7847),
        VN2CN0_sign => VN_sign_out(7842),
        VN2CN1_sign => VN_sign_out(7843),
        VN2CN2_sign => VN_sign_out(7844),
        VN2CN3_sign => VN_sign_out(7845),
        VN2CN4_sign => VN_sign_out(7846),
        VN2CN5_sign => VN_sign_out(7847),
        codeword => codeword(1307),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1308 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7853 downto 7848),
        Din0 => VN1308_in0,
        Din1 => VN1308_in1,
        Din2 => VN1308_in2,
        Din3 => VN1308_in3,
        Din4 => VN1308_in4,
        Din5 => VN1308_in5,
        VN2CN0_bit => VN_data_out(7848),
        VN2CN1_bit => VN_data_out(7849),
        VN2CN2_bit => VN_data_out(7850),
        VN2CN3_bit => VN_data_out(7851),
        VN2CN4_bit => VN_data_out(7852),
        VN2CN5_bit => VN_data_out(7853),
        VN2CN0_sign => VN_sign_out(7848),
        VN2CN1_sign => VN_sign_out(7849),
        VN2CN2_sign => VN_sign_out(7850),
        VN2CN3_sign => VN_sign_out(7851),
        VN2CN4_sign => VN_sign_out(7852),
        VN2CN5_sign => VN_sign_out(7853),
        codeword => codeword(1308),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1309 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7859 downto 7854),
        Din0 => VN1309_in0,
        Din1 => VN1309_in1,
        Din2 => VN1309_in2,
        Din3 => VN1309_in3,
        Din4 => VN1309_in4,
        Din5 => VN1309_in5,
        VN2CN0_bit => VN_data_out(7854),
        VN2CN1_bit => VN_data_out(7855),
        VN2CN2_bit => VN_data_out(7856),
        VN2CN3_bit => VN_data_out(7857),
        VN2CN4_bit => VN_data_out(7858),
        VN2CN5_bit => VN_data_out(7859),
        VN2CN0_sign => VN_sign_out(7854),
        VN2CN1_sign => VN_sign_out(7855),
        VN2CN2_sign => VN_sign_out(7856),
        VN2CN3_sign => VN_sign_out(7857),
        VN2CN4_sign => VN_sign_out(7858),
        VN2CN5_sign => VN_sign_out(7859),
        codeword => codeword(1309),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1310 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7865 downto 7860),
        Din0 => VN1310_in0,
        Din1 => VN1310_in1,
        Din2 => VN1310_in2,
        Din3 => VN1310_in3,
        Din4 => VN1310_in4,
        Din5 => VN1310_in5,
        VN2CN0_bit => VN_data_out(7860),
        VN2CN1_bit => VN_data_out(7861),
        VN2CN2_bit => VN_data_out(7862),
        VN2CN3_bit => VN_data_out(7863),
        VN2CN4_bit => VN_data_out(7864),
        VN2CN5_bit => VN_data_out(7865),
        VN2CN0_sign => VN_sign_out(7860),
        VN2CN1_sign => VN_sign_out(7861),
        VN2CN2_sign => VN_sign_out(7862),
        VN2CN3_sign => VN_sign_out(7863),
        VN2CN4_sign => VN_sign_out(7864),
        VN2CN5_sign => VN_sign_out(7865),
        codeword => codeword(1310),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1311 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7871 downto 7866),
        Din0 => VN1311_in0,
        Din1 => VN1311_in1,
        Din2 => VN1311_in2,
        Din3 => VN1311_in3,
        Din4 => VN1311_in4,
        Din5 => VN1311_in5,
        VN2CN0_bit => VN_data_out(7866),
        VN2CN1_bit => VN_data_out(7867),
        VN2CN2_bit => VN_data_out(7868),
        VN2CN3_bit => VN_data_out(7869),
        VN2CN4_bit => VN_data_out(7870),
        VN2CN5_bit => VN_data_out(7871),
        VN2CN0_sign => VN_sign_out(7866),
        VN2CN1_sign => VN_sign_out(7867),
        VN2CN2_sign => VN_sign_out(7868),
        VN2CN3_sign => VN_sign_out(7869),
        VN2CN4_sign => VN_sign_out(7870),
        VN2CN5_sign => VN_sign_out(7871),
        codeword => codeword(1311),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1312 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7877 downto 7872),
        Din0 => VN1312_in0,
        Din1 => VN1312_in1,
        Din2 => VN1312_in2,
        Din3 => VN1312_in3,
        Din4 => VN1312_in4,
        Din5 => VN1312_in5,
        VN2CN0_bit => VN_data_out(7872),
        VN2CN1_bit => VN_data_out(7873),
        VN2CN2_bit => VN_data_out(7874),
        VN2CN3_bit => VN_data_out(7875),
        VN2CN4_bit => VN_data_out(7876),
        VN2CN5_bit => VN_data_out(7877),
        VN2CN0_sign => VN_sign_out(7872),
        VN2CN1_sign => VN_sign_out(7873),
        VN2CN2_sign => VN_sign_out(7874),
        VN2CN3_sign => VN_sign_out(7875),
        VN2CN4_sign => VN_sign_out(7876),
        VN2CN5_sign => VN_sign_out(7877),
        codeword => codeword(1312),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1313 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7883 downto 7878),
        Din0 => VN1313_in0,
        Din1 => VN1313_in1,
        Din2 => VN1313_in2,
        Din3 => VN1313_in3,
        Din4 => VN1313_in4,
        Din5 => VN1313_in5,
        VN2CN0_bit => VN_data_out(7878),
        VN2CN1_bit => VN_data_out(7879),
        VN2CN2_bit => VN_data_out(7880),
        VN2CN3_bit => VN_data_out(7881),
        VN2CN4_bit => VN_data_out(7882),
        VN2CN5_bit => VN_data_out(7883),
        VN2CN0_sign => VN_sign_out(7878),
        VN2CN1_sign => VN_sign_out(7879),
        VN2CN2_sign => VN_sign_out(7880),
        VN2CN3_sign => VN_sign_out(7881),
        VN2CN4_sign => VN_sign_out(7882),
        VN2CN5_sign => VN_sign_out(7883),
        codeword => codeword(1313),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1314 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7889 downto 7884),
        Din0 => VN1314_in0,
        Din1 => VN1314_in1,
        Din2 => VN1314_in2,
        Din3 => VN1314_in3,
        Din4 => VN1314_in4,
        Din5 => VN1314_in5,
        VN2CN0_bit => VN_data_out(7884),
        VN2CN1_bit => VN_data_out(7885),
        VN2CN2_bit => VN_data_out(7886),
        VN2CN3_bit => VN_data_out(7887),
        VN2CN4_bit => VN_data_out(7888),
        VN2CN5_bit => VN_data_out(7889),
        VN2CN0_sign => VN_sign_out(7884),
        VN2CN1_sign => VN_sign_out(7885),
        VN2CN2_sign => VN_sign_out(7886),
        VN2CN3_sign => VN_sign_out(7887),
        VN2CN4_sign => VN_sign_out(7888),
        VN2CN5_sign => VN_sign_out(7889),
        codeword => codeword(1314),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1315 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7895 downto 7890),
        Din0 => VN1315_in0,
        Din1 => VN1315_in1,
        Din2 => VN1315_in2,
        Din3 => VN1315_in3,
        Din4 => VN1315_in4,
        Din5 => VN1315_in5,
        VN2CN0_bit => VN_data_out(7890),
        VN2CN1_bit => VN_data_out(7891),
        VN2CN2_bit => VN_data_out(7892),
        VN2CN3_bit => VN_data_out(7893),
        VN2CN4_bit => VN_data_out(7894),
        VN2CN5_bit => VN_data_out(7895),
        VN2CN0_sign => VN_sign_out(7890),
        VN2CN1_sign => VN_sign_out(7891),
        VN2CN2_sign => VN_sign_out(7892),
        VN2CN3_sign => VN_sign_out(7893),
        VN2CN4_sign => VN_sign_out(7894),
        VN2CN5_sign => VN_sign_out(7895),
        codeword => codeword(1315),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1316 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7901 downto 7896),
        Din0 => VN1316_in0,
        Din1 => VN1316_in1,
        Din2 => VN1316_in2,
        Din3 => VN1316_in3,
        Din4 => VN1316_in4,
        Din5 => VN1316_in5,
        VN2CN0_bit => VN_data_out(7896),
        VN2CN1_bit => VN_data_out(7897),
        VN2CN2_bit => VN_data_out(7898),
        VN2CN3_bit => VN_data_out(7899),
        VN2CN4_bit => VN_data_out(7900),
        VN2CN5_bit => VN_data_out(7901),
        VN2CN0_sign => VN_sign_out(7896),
        VN2CN1_sign => VN_sign_out(7897),
        VN2CN2_sign => VN_sign_out(7898),
        VN2CN3_sign => VN_sign_out(7899),
        VN2CN4_sign => VN_sign_out(7900),
        VN2CN5_sign => VN_sign_out(7901),
        codeword => codeword(1316),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1317 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7907 downto 7902),
        Din0 => VN1317_in0,
        Din1 => VN1317_in1,
        Din2 => VN1317_in2,
        Din3 => VN1317_in3,
        Din4 => VN1317_in4,
        Din5 => VN1317_in5,
        VN2CN0_bit => VN_data_out(7902),
        VN2CN1_bit => VN_data_out(7903),
        VN2CN2_bit => VN_data_out(7904),
        VN2CN3_bit => VN_data_out(7905),
        VN2CN4_bit => VN_data_out(7906),
        VN2CN5_bit => VN_data_out(7907),
        VN2CN0_sign => VN_sign_out(7902),
        VN2CN1_sign => VN_sign_out(7903),
        VN2CN2_sign => VN_sign_out(7904),
        VN2CN3_sign => VN_sign_out(7905),
        VN2CN4_sign => VN_sign_out(7906),
        VN2CN5_sign => VN_sign_out(7907),
        codeword => codeword(1317),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1318 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7913 downto 7908),
        Din0 => VN1318_in0,
        Din1 => VN1318_in1,
        Din2 => VN1318_in2,
        Din3 => VN1318_in3,
        Din4 => VN1318_in4,
        Din5 => VN1318_in5,
        VN2CN0_bit => VN_data_out(7908),
        VN2CN1_bit => VN_data_out(7909),
        VN2CN2_bit => VN_data_out(7910),
        VN2CN3_bit => VN_data_out(7911),
        VN2CN4_bit => VN_data_out(7912),
        VN2CN5_bit => VN_data_out(7913),
        VN2CN0_sign => VN_sign_out(7908),
        VN2CN1_sign => VN_sign_out(7909),
        VN2CN2_sign => VN_sign_out(7910),
        VN2CN3_sign => VN_sign_out(7911),
        VN2CN4_sign => VN_sign_out(7912),
        VN2CN5_sign => VN_sign_out(7913),
        codeword => codeword(1318),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1319 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7919 downto 7914),
        Din0 => VN1319_in0,
        Din1 => VN1319_in1,
        Din2 => VN1319_in2,
        Din3 => VN1319_in3,
        Din4 => VN1319_in4,
        Din5 => VN1319_in5,
        VN2CN0_bit => VN_data_out(7914),
        VN2CN1_bit => VN_data_out(7915),
        VN2CN2_bit => VN_data_out(7916),
        VN2CN3_bit => VN_data_out(7917),
        VN2CN4_bit => VN_data_out(7918),
        VN2CN5_bit => VN_data_out(7919),
        VN2CN0_sign => VN_sign_out(7914),
        VN2CN1_sign => VN_sign_out(7915),
        VN2CN2_sign => VN_sign_out(7916),
        VN2CN3_sign => VN_sign_out(7917),
        VN2CN4_sign => VN_sign_out(7918),
        VN2CN5_sign => VN_sign_out(7919),
        codeword => codeword(1319),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1320 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7925 downto 7920),
        Din0 => VN1320_in0,
        Din1 => VN1320_in1,
        Din2 => VN1320_in2,
        Din3 => VN1320_in3,
        Din4 => VN1320_in4,
        Din5 => VN1320_in5,
        VN2CN0_bit => VN_data_out(7920),
        VN2CN1_bit => VN_data_out(7921),
        VN2CN2_bit => VN_data_out(7922),
        VN2CN3_bit => VN_data_out(7923),
        VN2CN4_bit => VN_data_out(7924),
        VN2CN5_bit => VN_data_out(7925),
        VN2CN0_sign => VN_sign_out(7920),
        VN2CN1_sign => VN_sign_out(7921),
        VN2CN2_sign => VN_sign_out(7922),
        VN2CN3_sign => VN_sign_out(7923),
        VN2CN4_sign => VN_sign_out(7924),
        VN2CN5_sign => VN_sign_out(7925),
        codeword => codeword(1320),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1321 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7931 downto 7926),
        Din0 => VN1321_in0,
        Din1 => VN1321_in1,
        Din2 => VN1321_in2,
        Din3 => VN1321_in3,
        Din4 => VN1321_in4,
        Din5 => VN1321_in5,
        VN2CN0_bit => VN_data_out(7926),
        VN2CN1_bit => VN_data_out(7927),
        VN2CN2_bit => VN_data_out(7928),
        VN2CN3_bit => VN_data_out(7929),
        VN2CN4_bit => VN_data_out(7930),
        VN2CN5_bit => VN_data_out(7931),
        VN2CN0_sign => VN_sign_out(7926),
        VN2CN1_sign => VN_sign_out(7927),
        VN2CN2_sign => VN_sign_out(7928),
        VN2CN3_sign => VN_sign_out(7929),
        VN2CN4_sign => VN_sign_out(7930),
        VN2CN5_sign => VN_sign_out(7931),
        codeword => codeword(1321),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1322 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7937 downto 7932),
        Din0 => VN1322_in0,
        Din1 => VN1322_in1,
        Din2 => VN1322_in2,
        Din3 => VN1322_in3,
        Din4 => VN1322_in4,
        Din5 => VN1322_in5,
        VN2CN0_bit => VN_data_out(7932),
        VN2CN1_bit => VN_data_out(7933),
        VN2CN2_bit => VN_data_out(7934),
        VN2CN3_bit => VN_data_out(7935),
        VN2CN4_bit => VN_data_out(7936),
        VN2CN5_bit => VN_data_out(7937),
        VN2CN0_sign => VN_sign_out(7932),
        VN2CN1_sign => VN_sign_out(7933),
        VN2CN2_sign => VN_sign_out(7934),
        VN2CN3_sign => VN_sign_out(7935),
        VN2CN4_sign => VN_sign_out(7936),
        VN2CN5_sign => VN_sign_out(7937),
        codeword => codeword(1322),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1323 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7943 downto 7938),
        Din0 => VN1323_in0,
        Din1 => VN1323_in1,
        Din2 => VN1323_in2,
        Din3 => VN1323_in3,
        Din4 => VN1323_in4,
        Din5 => VN1323_in5,
        VN2CN0_bit => VN_data_out(7938),
        VN2CN1_bit => VN_data_out(7939),
        VN2CN2_bit => VN_data_out(7940),
        VN2CN3_bit => VN_data_out(7941),
        VN2CN4_bit => VN_data_out(7942),
        VN2CN5_bit => VN_data_out(7943),
        VN2CN0_sign => VN_sign_out(7938),
        VN2CN1_sign => VN_sign_out(7939),
        VN2CN2_sign => VN_sign_out(7940),
        VN2CN3_sign => VN_sign_out(7941),
        VN2CN4_sign => VN_sign_out(7942),
        VN2CN5_sign => VN_sign_out(7943),
        codeword => codeword(1323),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1324 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7949 downto 7944),
        Din0 => VN1324_in0,
        Din1 => VN1324_in1,
        Din2 => VN1324_in2,
        Din3 => VN1324_in3,
        Din4 => VN1324_in4,
        Din5 => VN1324_in5,
        VN2CN0_bit => VN_data_out(7944),
        VN2CN1_bit => VN_data_out(7945),
        VN2CN2_bit => VN_data_out(7946),
        VN2CN3_bit => VN_data_out(7947),
        VN2CN4_bit => VN_data_out(7948),
        VN2CN5_bit => VN_data_out(7949),
        VN2CN0_sign => VN_sign_out(7944),
        VN2CN1_sign => VN_sign_out(7945),
        VN2CN2_sign => VN_sign_out(7946),
        VN2CN3_sign => VN_sign_out(7947),
        VN2CN4_sign => VN_sign_out(7948),
        VN2CN5_sign => VN_sign_out(7949),
        codeword => codeword(1324),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1325 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7955 downto 7950),
        Din0 => VN1325_in0,
        Din1 => VN1325_in1,
        Din2 => VN1325_in2,
        Din3 => VN1325_in3,
        Din4 => VN1325_in4,
        Din5 => VN1325_in5,
        VN2CN0_bit => VN_data_out(7950),
        VN2CN1_bit => VN_data_out(7951),
        VN2CN2_bit => VN_data_out(7952),
        VN2CN3_bit => VN_data_out(7953),
        VN2CN4_bit => VN_data_out(7954),
        VN2CN5_bit => VN_data_out(7955),
        VN2CN0_sign => VN_sign_out(7950),
        VN2CN1_sign => VN_sign_out(7951),
        VN2CN2_sign => VN_sign_out(7952),
        VN2CN3_sign => VN_sign_out(7953),
        VN2CN4_sign => VN_sign_out(7954),
        VN2CN5_sign => VN_sign_out(7955),
        codeword => codeword(1325),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1326 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7961 downto 7956),
        Din0 => VN1326_in0,
        Din1 => VN1326_in1,
        Din2 => VN1326_in2,
        Din3 => VN1326_in3,
        Din4 => VN1326_in4,
        Din5 => VN1326_in5,
        VN2CN0_bit => VN_data_out(7956),
        VN2CN1_bit => VN_data_out(7957),
        VN2CN2_bit => VN_data_out(7958),
        VN2CN3_bit => VN_data_out(7959),
        VN2CN4_bit => VN_data_out(7960),
        VN2CN5_bit => VN_data_out(7961),
        VN2CN0_sign => VN_sign_out(7956),
        VN2CN1_sign => VN_sign_out(7957),
        VN2CN2_sign => VN_sign_out(7958),
        VN2CN3_sign => VN_sign_out(7959),
        VN2CN4_sign => VN_sign_out(7960),
        VN2CN5_sign => VN_sign_out(7961),
        codeword => codeword(1326),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1327 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7967 downto 7962),
        Din0 => VN1327_in0,
        Din1 => VN1327_in1,
        Din2 => VN1327_in2,
        Din3 => VN1327_in3,
        Din4 => VN1327_in4,
        Din5 => VN1327_in5,
        VN2CN0_bit => VN_data_out(7962),
        VN2CN1_bit => VN_data_out(7963),
        VN2CN2_bit => VN_data_out(7964),
        VN2CN3_bit => VN_data_out(7965),
        VN2CN4_bit => VN_data_out(7966),
        VN2CN5_bit => VN_data_out(7967),
        VN2CN0_sign => VN_sign_out(7962),
        VN2CN1_sign => VN_sign_out(7963),
        VN2CN2_sign => VN_sign_out(7964),
        VN2CN3_sign => VN_sign_out(7965),
        VN2CN4_sign => VN_sign_out(7966),
        VN2CN5_sign => VN_sign_out(7967),
        codeword => codeword(1327),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1328 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7973 downto 7968),
        Din0 => VN1328_in0,
        Din1 => VN1328_in1,
        Din2 => VN1328_in2,
        Din3 => VN1328_in3,
        Din4 => VN1328_in4,
        Din5 => VN1328_in5,
        VN2CN0_bit => VN_data_out(7968),
        VN2CN1_bit => VN_data_out(7969),
        VN2CN2_bit => VN_data_out(7970),
        VN2CN3_bit => VN_data_out(7971),
        VN2CN4_bit => VN_data_out(7972),
        VN2CN5_bit => VN_data_out(7973),
        VN2CN0_sign => VN_sign_out(7968),
        VN2CN1_sign => VN_sign_out(7969),
        VN2CN2_sign => VN_sign_out(7970),
        VN2CN3_sign => VN_sign_out(7971),
        VN2CN4_sign => VN_sign_out(7972),
        VN2CN5_sign => VN_sign_out(7973),
        codeword => codeword(1328),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1329 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7979 downto 7974),
        Din0 => VN1329_in0,
        Din1 => VN1329_in1,
        Din2 => VN1329_in2,
        Din3 => VN1329_in3,
        Din4 => VN1329_in4,
        Din5 => VN1329_in5,
        VN2CN0_bit => VN_data_out(7974),
        VN2CN1_bit => VN_data_out(7975),
        VN2CN2_bit => VN_data_out(7976),
        VN2CN3_bit => VN_data_out(7977),
        VN2CN4_bit => VN_data_out(7978),
        VN2CN5_bit => VN_data_out(7979),
        VN2CN0_sign => VN_sign_out(7974),
        VN2CN1_sign => VN_sign_out(7975),
        VN2CN2_sign => VN_sign_out(7976),
        VN2CN3_sign => VN_sign_out(7977),
        VN2CN4_sign => VN_sign_out(7978),
        VN2CN5_sign => VN_sign_out(7979),
        codeword => codeword(1329),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1330 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7985 downto 7980),
        Din0 => VN1330_in0,
        Din1 => VN1330_in1,
        Din2 => VN1330_in2,
        Din3 => VN1330_in3,
        Din4 => VN1330_in4,
        Din5 => VN1330_in5,
        VN2CN0_bit => VN_data_out(7980),
        VN2CN1_bit => VN_data_out(7981),
        VN2CN2_bit => VN_data_out(7982),
        VN2CN3_bit => VN_data_out(7983),
        VN2CN4_bit => VN_data_out(7984),
        VN2CN5_bit => VN_data_out(7985),
        VN2CN0_sign => VN_sign_out(7980),
        VN2CN1_sign => VN_sign_out(7981),
        VN2CN2_sign => VN_sign_out(7982),
        VN2CN3_sign => VN_sign_out(7983),
        VN2CN4_sign => VN_sign_out(7984),
        VN2CN5_sign => VN_sign_out(7985),
        codeword => codeword(1330),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1331 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7991 downto 7986),
        Din0 => VN1331_in0,
        Din1 => VN1331_in1,
        Din2 => VN1331_in2,
        Din3 => VN1331_in3,
        Din4 => VN1331_in4,
        Din5 => VN1331_in5,
        VN2CN0_bit => VN_data_out(7986),
        VN2CN1_bit => VN_data_out(7987),
        VN2CN2_bit => VN_data_out(7988),
        VN2CN3_bit => VN_data_out(7989),
        VN2CN4_bit => VN_data_out(7990),
        VN2CN5_bit => VN_data_out(7991),
        VN2CN0_sign => VN_sign_out(7986),
        VN2CN1_sign => VN_sign_out(7987),
        VN2CN2_sign => VN_sign_out(7988),
        VN2CN3_sign => VN_sign_out(7989),
        VN2CN4_sign => VN_sign_out(7990),
        VN2CN5_sign => VN_sign_out(7991),
        codeword => codeword(1331),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1332 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(7997 downto 7992),
        Din0 => VN1332_in0,
        Din1 => VN1332_in1,
        Din2 => VN1332_in2,
        Din3 => VN1332_in3,
        Din4 => VN1332_in4,
        Din5 => VN1332_in5,
        VN2CN0_bit => VN_data_out(7992),
        VN2CN1_bit => VN_data_out(7993),
        VN2CN2_bit => VN_data_out(7994),
        VN2CN3_bit => VN_data_out(7995),
        VN2CN4_bit => VN_data_out(7996),
        VN2CN5_bit => VN_data_out(7997),
        VN2CN0_sign => VN_sign_out(7992),
        VN2CN1_sign => VN_sign_out(7993),
        VN2CN2_sign => VN_sign_out(7994),
        VN2CN3_sign => VN_sign_out(7995),
        VN2CN4_sign => VN_sign_out(7996),
        VN2CN5_sign => VN_sign_out(7997),
        codeword => codeword(1332),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1333 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8003 downto 7998),
        Din0 => VN1333_in0,
        Din1 => VN1333_in1,
        Din2 => VN1333_in2,
        Din3 => VN1333_in3,
        Din4 => VN1333_in4,
        Din5 => VN1333_in5,
        VN2CN0_bit => VN_data_out(7998),
        VN2CN1_bit => VN_data_out(7999),
        VN2CN2_bit => VN_data_out(8000),
        VN2CN3_bit => VN_data_out(8001),
        VN2CN4_bit => VN_data_out(8002),
        VN2CN5_bit => VN_data_out(8003),
        VN2CN0_sign => VN_sign_out(7998),
        VN2CN1_sign => VN_sign_out(7999),
        VN2CN2_sign => VN_sign_out(8000),
        VN2CN3_sign => VN_sign_out(8001),
        VN2CN4_sign => VN_sign_out(8002),
        VN2CN5_sign => VN_sign_out(8003),
        codeword => codeword(1333),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1334 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8009 downto 8004),
        Din0 => VN1334_in0,
        Din1 => VN1334_in1,
        Din2 => VN1334_in2,
        Din3 => VN1334_in3,
        Din4 => VN1334_in4,
        Din5 => VN1334_in5,
        VN2CN0_bit => VN_data_out(8004),
        VN2CN1_bit => VN_data_out(8005),
        VN2CN2_bit => VN_data_out(8006),
        VN2CN3_bit => VN_data_out(8007),
        VN2CN4_bit => VN_data_out(8008),
        VN2CN5_bit => VN_data_out(8009),
        VN2CN0_sign => VN_sign_out(8004),
        VN2CN1_sign => VN_sign_out(8005),
        VN2CN2_sign => VN_sign_out(8006),
        VN2CN3_sign => VN_sign_out(8007),
        VN2CN4_sign => VN_sign_out(8008),
        VN2CN5_sign => VN_sign_out(8009),
        codeword => codeword(1334),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1335 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8015 downto 8010),
        Din0 => VN1335_in0,
        Din1 => VN1335_in1,
        Din2 => VN1335_in2,
        Din3 => VN1335_in3,
        Din4 => VN1335_in4,
        Din5 => VN1335_in5,
        VN2CN0_bit => VN_data_out(8010),
        VN2CN1_bit => VN_data_out(8011),
        VN2CN2_bit => VN_data_out(8012),
        VN2CN3_bit => VN_data_out(8013),
        VN2CN4_bit => VN_data_out(8014),
        VN2CN5_bit => VN_data_out(8015),
        VN2CN0_sign => VN_sign_out(8010),
        VN2CN1_sign => VN_sign_out(8011),
        VN2CN2_sign => VN_sign_out(8012),
        VN2CN3_sign => VN_sign_out(8013),
        VN2CN4_sign => VN_sign_out(8014),
        VN2CN5_sign => VN_sign_out(8015),
        codeword => codeword(1335),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1336 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8021 downto 8016),
        Din0 => VN1336_in0,
        Din1 => VN1336_in1,
        Din2 => VN1336_in2,
        Din3 => VN1336_in3,
        Din4 => VN1336_in4,
        Din5 => VN1336_in5,
        VN2CN0_bit => VN_data_out(8016),
        VN2CN1_bit => VN_data_out(8017),
        VN2CN2_bit => VN_data_out(8018),
        VN2CN3_bit => VN_data_out(8019),
        VN2CN4_bit => VN_data_out(8020),
        VN2CN5_bit => VN_data_out(8021),
        VN2CN0_sign => VN_sign_out(8016),
        VN2CN1_sign => VN_sign_out(8017),
        VN2CN2_sign => VN_sign_out(8018),
        VN2CN3_sign => VN_sign_out(8019),
        VN2CN4_sign => VN_sign_out(8020),
        VN2CN5_sign => VN_sign_out(8021),
        codeword => codeword(1336),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1337 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8027 downto 8022),
        Din0 => VN1337_in0,
        Din1 => VN1337_in1,
        Din2 => VN1337_in2,
        Din3 => VN1337_in3,
        Din4 => VN1337_in4,
        Din5 => VN1337_in5,
        VN2CN0_bit => VN_data_out(8022),
        VN2CN1_bit => VN_data_out(8023),
        VN2CN2_bit => VN_data_out(8024),
        VN2CN3_bit => VN_data_out(8025),
        VN2CN4_bit => VN_data_out(8026),
        VN2CN5_bit => VN_data_out(8027),
        VN2CN0_sign => VN_sign_out(8022),
        VN2CN1_sign => VN_sign_out(8023),
        VN2CN2_sign => VN_sign_out(8024),
        VN2CN3_sign => VN_sign_out(8025),
        VN2CN4_sign => VN_sign_out(8026),
        VN2CN5_sign => VN_sign_out(8027),
        codeword => codeword(1337),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1338 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8033 downto 8028),
        Din0 => VN1338_in0,
        Din1 => VN1338_in1,
        Din2 => VN1338_in2,
        Din3 => VN1338_in3,
        Din4 => VN1338_in4,
        Din5 => VN1338_in5,
        VN2CN0_bit => VN_data_out(8028),
        VN2CN1_bit => VN_data_out(8029),
        VN2CN2_bit => VN_data_out(8030),
        VN2CN3_bit => VN_data_out(8031),
        VN2CN4_bit => VN_data_out(8032),
        VN2CN5_bit => VN_data_out(8033),
        VN2CN0_sign => VN_sign_out(8028),
        VN2CN1_sign => VN_sign_out(8029),
        VN2CN2_sign => VN_sign_out(8030),
        VN2CN3_sign => VN_sign_out(8031),
        VN2CN4_sign => VN_sign_out(8032),
        VN2CN5_sign => VN_sign_out(8033),
        codeword => codeword(1338),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1339 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8039 downto 8034),
        Din0 => VN1339_in0,
        Din1 => VN1339_in1,
        Din2 => VN1339_in2,
        Din3 => VN1339_in3,
        Din4 => VN1339_in4,
        Din5 => VN1339_in5,
        VN2CN0_bit => VN_data_out(8034),
        VN2CN1_bit => VN_data_out(8035),
        VN2CN2_bit => VN_data_out(8036),
        VN2CN3_bit => VN_data_out(8037),
        VN2CN4_bit => VN_data_out(8038),
        VN2CN5_bit => VN_data_out(8039),
        VN2CN0_sign => VN_sign_out(8034),
        VN2CN1_sign => VN_sign_out(8035),
        VN2CN2_sign => VN_sign_out(8036),
        VN2CN3_sign => VN_sign_out(8037),
        VN2CN4_sign => VN_sign_out(8038),
        VN2CN5_sign => VN_sign_out(8039),
        codeword => codeword(1339),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1340 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8045 downto 8040),
        Din0 => VN1340_in0,
        Din1 => VN1340_in1,
        Din2 => VN1340_in2,
        Din3 => VN1340_in3,
        Din4 => VN1340_in4,
        Din5 => VN1340_in5,
        VN2CN0_bit => VN_data_out(8040),
        VN2CN1_bit => VN_data_out(8041),
        VN2CN2_bit => VN_data_out(8042),
        VN2CN3_bit => VN_data_out(8043),
        VN2CN4_bit => VN_data_out(8044),
        VN2CN5_bit => VN_data_out(8045),
        VN2CN0_sign => VN_sign_out(8040),
        VN2CN1_sign => VN_sign_out(8041),
        VN2CN2_sign => VN_sign_out(8042),
        VN2CN3_sign => VN_sign_out(8043),
        VN2CN4_sign => VN_sign_out(8044),
        VN2CN5_sign => VN_sign_out(8045),
        codeword => codeword(1340),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1341 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8051 downto 8046),
        Din0 => VN1341_in0,
        Din1 => VN1341_in1,
        Din2 => VN1341_in2,
        Din3 => VN1341_in3,
        Din4 => VN1341_in4,
        Din5 => VN1341_in5,
        VN2CN0_bit => VN_data_out(8046),
        VN2CN1_bit => VN_data_out(8047),
        VN2CN2_bit => VN_data_out(8048),
        VN2CN3_bit => VN_data_out(8049),
        VN2CN4_bit => VN_data_out(8050),
        VN2CN5_bit => VN_data_out(8051),
        VN2CN0_sign => VN_sign_out(8046),
        VN2CN1_sign => VN_sign_out(8047),
        VN2CN2_sign => VN_sign_out(8048),
        VN2CN3_sign => VN_sign_out(8049),
        VN2CN4_sign => VN_sign_out(8050),
        VN2CN5_sign => VN_sign_out(8051),
        codeword => codeword(1341),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1342 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8057 downto 8052),
        Din0 => VN1342_in0,
        Din1 => VN1342_in1,
        Din2 => VN1342_in2,
        Din3 => VN1342_in3,
        Din4 => VN1342_in4,
        Din5 => VN1342_in5,
        VN2CN0_bit => VN_data_out(8052),
        VN2CN1_bit => VN_data_out(8053),
        VN2CN2_bit => VN_data_out(8054),
        VN2CN3_bit => VN_data_out(8055),
        VN2CN4_bit => VN_data_out(8056),
        VN2CN5_bit => VN_data_out(8057),
        VN2CN0_sign => VN_sign_out(8052),
        VN2CN1_sign => VN_sign_out(8053),
        VN2CN2_sign => VN_sign_out(8054),
        VN2CN3_sign => VN_sign_out(8055),
        VN2CN4_sign => VN_sign_out(8056),
        VN2CN5_sign => VN_sign_out(8057),
        codeword => codeword(1342),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1343 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8063 downto 8058),
        Din0 => VN1343_in0,
        Din1 => VN1343_in1,
        Din2 => VN1343_in2,
        Din3 => VN1343_in3,
        Din4 => VN1343_in4,
        Din5 => VN1343_in5,
        VN2CN0_bit => VN_data_out(8058),
        VN2CN1_bit => VN_data_out(8059),
        VN2CN2_bit => VN_data_out(8060),
        VN2CN3_bit => VN_data_out(8061),
        VN2CN4_bit => VN_data_out(8062),
        VN2CN5_bit => VN_data_out(8063),
        VN2CN0_sign => VN_sign_out(8058),
        VN2CN1_sign => VN_sign_out(8059),
        VN2CN2_sign => VN_sign_out(8060),
        VN2CN3_sign => VN_sign_out(8061),
        VN2CN4_sign => VN_sign_out(8062),
        VN2CN5_sign => VN_sign_out(8063),
        codeword => codeword(1343),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1344 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8069 downto 8064),
        Din0 => VN1344_in0,
        Din1 => VN1344_in1,
        Din2 => VN1344_in2,
        Din3 => VN1344_in3,
        Din4 => VN1344_in4,
        Din5 => VN1344_in5,
        VN2CN0_bit => VN_data_out(8064),
        VN2CN1_bit => VN_data_out(8065),
        VN2CN2_bit => VN_data_out(8066),
        VN2CN3_bit => VN_data_out(8067),
        VN2CN4_bit => VN_data_out(8068),
        VN2CN5_bit => VN_data_out(8069),
        VN2CN0_sign => VN_sign_out(8064),
        VN2CN1_sign => VN_sign_out(8065),
        VN2CN2_sign => VN_sign_out(8066),
        VN2CN3_sign => VN_sign_out(8067),
        VN2CN4_sign => VN_sign_out(8068),
        VN2CN5_sign => VN_sign_out(8069),
        codeword => codeword(1344),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1345 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8075 downto 8070),
        Din0 => VN1345_in0,
        Din1 => VN1345_in1,
        Din2 => VN1345_in2,
        Din3 => VN1345_in3,
        Din4 => VN1345_in4,
        Din5 => VN1345_in5,
        VN2CN0_bit => VN_data_out(8070),
        VN2CN1_bit => VN_data_out(8071),
        VN2CN2_bit => VN_data_out(8072),
        VN2CN3_bit => VN_data_out(8073),
        VN2CN4_bit => VN_data_out(8074),
        VN2CN5_bit => VN_data_out(8075),
        VN2CN0_sign => VN_sign_out(8070),
        VN2CN1_sign => VN_sign_out(8071),
        VN2CN2_sign => VN_sign_out(8072),
        VN2CN3_sign => VN_sign_out(8073),
        VN2CN4_sign => VN_sign_out(8074),
        VN2CN5_sign => VN_sign_out(8075),
        codeword => codeword(1345),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1346 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8081 downto 8076),
        Din0 => VN1346_in0,
        Din1 => VN1346_in1,
        Din2 => VN1346_in2,
        Din3 => VN1346_in3,
        Din4 => VN1346_in4,
        Din5 => VN1346_in5,
        VN2CN0_bit => VN_data_out(8076),
        VN2CN1_bit => VN_data_out(8077),
        VN2CN2_bit => VN_data_out(8078),
        VN2CN3_bit => VN_data_out(8079),
        VN2CN4_bit => VN_data_out(8080),
        VN2CN5_bit => VN_data_out(8081),
        VN2CN0_sign => VN_sign_out(8076),
        VN2CN1_sign => VN_sign_out(8077),
        VN2CN2_sign => VN_sign_out(8078),
        VN2CN3_sign => VN_sign_out(8079),
        VN2CN4_sign => VN_sign_out(8080),
        VN2CN5_sign => VN_sign_out(8081),
        codeword => codeword(1346),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1347 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8087 downto 8082),
        Din0 => VN1347_in0,
        Din1 => VN1347_in1,
        Din2 => VN1347_in2,
        Din3 => VN1347_in3,
        Din4 => VN1347_in4,
        Din5 => VN1347_in5,
        VN2CN0_bit => VN_data_out(8082),
        VN2CN1_bit => VN_data_out(8083),
        VN2CN2_bit => VN_data_out(8084),
        VN2CN3_bit => VN_data_out(8085),
        VN2CN4_bit => VN_data_out(8086),
        VN2CN5_bit => VN_data_out(8087),
        VN2CN0_sign => VN_sign_out(8082),
        VN2CN1_sign => VN_sign_out(8083),
        VN2CN2_sign => VN_sign_out(8084),
        VN2CN3_sign => VN_sign_out(8085),
        VN2CN4_sign => VN_sign_out(8086),
        VN2CN5_sign => VN_sign_out(8087),
        codeword => codeword(1347),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1348 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8093 downto 8088),
        Din0 => VN1348_in0,
        Din1 => VN1348_in1,
        Din2 => VN1348_in2,
        Din3 => VN1348_in3,
        Din4 => VN1348_in4,
        Din5 => VN1348_in5,
        VN2CN0_bit => VN_data_out(8088),
        VN2CN1_bit => VN_data_out(8089),
        VN2CN2_bit => VN_data_out(8090),
        VN2CN3_bit => VN_data_out(8091),
        VN2CN4_bit => VN_data_out(8092),
        VN2CN5_bit => VN_data_out(8093),
        VN2CN0_sign => VN_sign_out(8088),
        VN2CN1_sign => VN_sign_out(8089),
        VN2CN2_sign => VN_sign_out(8090),
        VN2CN3_sign => VN_sign_out(8091),
        VN2CN4_sign => VN_sign_out(8092),
        VN2CN5_sign => VN_sign_out(8093),
        codeword => codeword(1348),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1349 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8099 downto 8094),
        Din0 => VN1349_in0,
        Din1 => VN1349_in1,
        Din2 => VN1349_in2,
        Din3 => VN1349_in3,
        Din4 => VN1349_in4,
        Din5 => VN1349_in5,
        VN2CN0_bit => VN_data_out(8094),
        VN2CN1_bit => VN_data_out(8095),
        VN2CN2_bit => VN_data_out(8096),
        VN2CN3_bit => VN_data_out(8097),
        VN2CN4_bit => VN_data_out(8098),
        VN2CN5_bit => VN_data_out(8099),
        VN2CN0_sign => VN_sign_out(8094),
        VN2CN1_sign => VN_sign_out(8095),
        VN2CN2_sign => VN_sign_out(8096),
        VN2CN3_sign => VN_sign_out(8097),
        VN2CN4_sign => VN_sign_out(8098),
        VN2CN5_sign => VN_sign_out(8099),
        codeword => codeword(1349),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1350 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8105 downto 8100),
        Din0 => VN1350_in0,
        Din1 => VN1350_in1,
        Din2 => VN1350_in2,
        Din3 => VN1350_in3,
        Din4 => VN1350_in4,
        Din5 => VN1350_in5,
        VN2CN0_bit => VN_data_out(8100),
        VN2CN1_bit => VN_data_out(8101),
        VN2CN2_bit => VN_data_out(8102),
        VN2CN3_bit => VN_data_out(8103),
        VN2CN4_bit => VN_data_out(8104),
        VN2CN5_bit => VN_data_out(8105),
        VN2CN0_sign => VN_sign_out(8100),
        VN2CN1_sign => VN_sign_out(8101),
        VN2CN2_sign => VN_sign_out(8102),
        VN2CN3_sign => VN_sign_out(8103),
        VN2CN4_sign => VN_sign_out(8104),
        VN2CN5_sign => VN_sign_out(8105),
        codeword => codeword(1350),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1351 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8111 downto 8106),
        Din0 => VN1351_in0,
        Din1 => VN1351_in1,
        Din2 => VN1351_in2,
        Din3 => VN1351_in3,
        Din4 => VN1351_in4,
        Din5 => VN1351_in5,
        VN2CN0_bit => VN_data_out(8106),
        VN2CN1_bit => VN_data_out(8107),
        VN2CN2_bit => VN_data_out(8108),
        VN2CN3_bit => VN_data_out(8109),
        VN2CN4_bit => VN_data_out(8110),
        VN2CN5_bit => VN_data_out(8111),
        VN2CN0_sign => VN_sign_out(8106),
        VN2CN1_sign => VN_sign_out(8107),
        VN2CN2_sign => VN_sign_out(8108),
        VN2CN3_sign => VN_sign_out(8109),
        VN2CN4_sign => VN_sign_out(8110),
        VN2CN5_sign => VN_sign_out(8111),
        codeword => codeword(1351),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1352 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8117 downto 8112),
        Din0 => VN1352_in0,
        Din1 => VN1352_in1,
        Din2 => VN1352_in2,
        Din3 => VN1352_in3,
        Din4 => VN1352_in4,
        Din5 => VN1352_in5,
        VN2CN0_bit => VN_data_out(8112),
        VN2CN1_bit => VN_data_out(8113),
        VN2CN2_bit => VN_data_out(8114),
        VN2CN3_bit => VN_data_out(8115),
        VN2CN4_bit => VN_data_out(8116),
        VN2CN5_bit => VN_data_out(8117),
        VN2CN0_sign => VN_sign_out(8112),
        VN2CN1_sign => VN_sign_out(8113),
        VN2CN2_sign => VN_sign_out(8114),
        VN2CN3_sign => VN_sign_out(8115),
        VN2CN4_sign => VN_sign_out(8116),
        VN2CN5_sign => VN_sign_out(8117),
        codeword => codeword(1352),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1353 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8123 downto 8118),
        Din0 => VN1353_in0,
        Din1 => VN1353_in1,
        Din2 => VN1353_in2,
        Din3 => VN1353_in3,
        Din4 => VN1353_in4,
        Din5 => VN1353_in5,
        VN2CN0_bit => VN_data_out(8118),
        VN2CN1_bit => VN_data_out(8119),
        VN2CN2_bit => VN_data_out(8120),
        VN2CN3_bit => VN_data_out(8121),
        VN2CN4_bit => VN_data_out(8122),
        VN2CN5_bit => VN_data_out(8123),
        VN2CN0_sign => VN_sign_out(8118),
        VN2CN1_sign => VN_sign_out(8119),
        VN2CN2_sign => VN_sign_out(8120),
        VN2CN3_sign => VN_sign_out(8121),
        VN2CN4_sign => VN_sign_out(8122),
        VN2CN5_sign => VN_sign_out(8123),
        codeword => codeword(1353),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1354 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8129 downto 8124),
        Din0 => VN1354_in0,
        Din1 => VN1354_in1,
        Din2 => VN1354_in2,
        Din3 => VN1354_in3,
        Din4 => VN1354_in4,
        Din5 => VN1354_in5,
        VN2CN0_bit => VN_data_out(8124),
        VN2CN1_bit => VN_data_out(8125),
        VN2CN2_bit => VN_data_out(8126),
        VN2CN3_bit => VN_data_out(8127),
        VN2CN4_bit => VN_data_out(8128),
        VN2CN5_bit => VN_data_out(8129),
        VN2CN0_sign => VN_sign_out(8124),
        VN2CN1_sign => VN_sign_out(8125),
        VN2CN2_sign => VN_sign_out(8126),
        VN2CN3_sign => VN_sign_out(8127),
        VN2CN4_sign => VN_sign_out(8128),
        VN2CN5_sign => VN_sign_out(8129),
        codeword => codeword(1354),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1355 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8135 downto 8130),
        Din0 => VN1355_in0,
        Din1 => VN1355_in1,
        Din2 => VN1355_in2,
        Din3 => VN1355_in3,
        Din4 => VN1355_in4,
        Din5 => VN1355_in5,
        VN2CN0_bit => VN_data_out(8130),
        VN2CN1_bit => VN_data_out(8131),
        VN2CN2_bit => VN_data_out(8132),
        VN2CN3_bit => VN_data_out(8133),
        VN2CN4_bit => VN_data_out(8134),
        VN2CN5_bit => VN_data_out(8135),
        VN2CN0_sign => VN_sign_out(8130),
        VN2CN1_sign => VN_sign_out(8131),
        VN2CN2_sign => VN_sign_out(8132),
        VN2CN3_sign => VN_sign_out(8133),
        VN2CN4_sign => VN_sign_out(8134),
        VN2CN5_sign => VN_sign_out(8135),
        codeword => codeword(1355),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1356 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8141 downto 8136),
        Din0 => VN1356_in0,
        Din1 => VN1356_in1,
        Din2 => VN1356_in2,
        Din3 => VN1356_in3,
        Din4 => VN1356_in4,
        Din5 => VN1356_in5,
        VN2CN0_bit => VN_data_out(8136),
        VN2CN1_bit => VN_data_out(8137),
        VN2CN2_bit => VN_data_out(8138),
        VN2CN3_bit => VN_data_out(8139),
        VN2CN4_bit => VN_data_out(8140),
        VN2CN5_bit => VN_data_out(8141),
        VN2CN0_sign => VN_sign_out(8136),
        VN2CN1_sign => VN_sign_out(8137),
        VN2CN2_sign => VN_sign_out(8138),
        VN2CN3_sign => VN_sign_out(8139),
        VN2CN4_sign => VN_sign_out(8140),
        VN2CN5_sign => VN_sign_out(8141),
        codeword => codeword(1356),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1357 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8147 downto 8142),
        Din0 => VN1357_in0,
        Din1 => VN1357_in1,
        Din2 => VN1357_in2,
        Din3 => VN1357_in3,
        Din4 => VN1357_in4,
        Din5 => VN1357_in5,
        VN2CN0_bit => VN_data_out(8142),
        VN2CN1_bit => VN_data_out(8143),
        VN2CN2_bit => VN_data_out(8144),
        VN2CN3_bit => VN_data_out(8145),
        VN2CN4_bit => VN_data_out(8146),
        VN2CN5_bit => VN_data_out(8147),
        VN2CN0_sign => VN_sign_out(8142),
        VN2CN1_sign => VN_sign_out(8143),
        VN2CN2_sign => VN_sign_out(8144),
        VN2CN3_sign => VN_sign_out(8145),
        VN2CN4_sign => VN_sign_out(8146),
        VN2CN5_sign => VN_sign_out(8147),
        codeword => codeword(1357),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1358 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8153 downto 8148),
        Din0 => VN1358_in0,
        Din1 => VN1358_in1,
        Din2 => VN1358_in2,
        Din3 => VN1358_in3,
        Din4 => VN1358_in4,
        Din5 => VN1358_in5,
        VN2CN0_bit => VN_data_out(8148),
        VN2CN1_bit => VN_data_out(8149),
        VN2CN2_bit => VN_data_out(8150),
        VN2CN3_bit => VN_data_out(8151),
        VN2CN4_bit => VN_data_out(8152),
        VN2CN5_bit => VN_data_out(8153),
        VN2CN0_sign => VN_sign_out(8148),
        VN2CN1_sign => VN_sign_out(8149),
        VN2CN2_sign => VN_sign_out(8150),
        VN2CN3_sign => VN_sign_out(8151),
        VN2CN4_sign => VN_sign_out(8152),
        VN2CN5_sign => VN_sign_out(8153),
        codeword => codeword(1358),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1359 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8159 downto 8154),
        Din0 => VN1359_in0,
        Din1 => VN1359_in1,
        Din2 => VN1359_in2,
        Din3 => VN1359_in3,
        Din4 => VN1359_in4,
        Din5 => VN1359_in5,
        VN2CN0_bit => VN_data_out(8154),
        VN2CN1_bit => VN_data_out(8155),
        VN2CN2_bit => VN_data_out(8156),
        VN2CN3_bit => VN_data_out(8157),
        VN2CN4_bit => VN_data_out(8158),
        VN2CN5_bit => VN_data_out(8159),
        VN2CN0_sign => VN_sign_out(8154),
        VN2CN1_sign => VN_sign_out(8155),
        VN2CN2_sign => VN_sign_out(8156),
        VN2CN3_sign => VN_sign_out(8157),
        VN2CN4_sign => VN_sign_out(8158),
        VN2CN5_sign => VN_sign_out(8159),
        codeword => codeword(1359),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1360 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8165 downto 8160),
        Din0 => VN1360_in0,
        Din1 => VN1360_in1,
        Din2 => VN1360_in2,
        Din3 => VN1360_in3,
        Din4 => VN1360_in4,
        Din5 => VN1360_in5,
        VN2CN0_bit => VN_data_out(8160),
        VN2CN1_bit => VN_data_out(8161),
        VN2CN2_bit => VN_data_out(8162),
        VN2CN3_bit => VN_data_out(8163),
        VN2CN4_bit => VN_data_out(8164),
        VN2CN5_bit => VN_data_out(8165),
        VN2CN0_sign => VN_sign_out(8160),
        VN2CN1_sign => VN_sign_out(8161),
        VN2CN2_sign => VN_sign_out(8162),
        VN2CN3_sign => VN_sign_out(8163),
        VN2CN4_sign => VN_sign_out(8164),
        VN2CN5_sign => VN_sign_out(8165),
        codeword => codeword(1360),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1361 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8171 downto 8166),
        Din0 => VN1361_in0,
        Din1 => VN1361_in1,
        Din2 => VN1361_in2,
        Din3 => VN1361_in3,
        Din4 => VN1361_in4,
        Din5 => VN1361_in5,
        VN2CN0_bit => VN_data_out(8166),
        VN2CN1_bit => VN_data_out(8167),
        VN2CN2_bit => VN_data_out(8168),
        VN2CN3_bit => VN_data_out(8169),
        VN2CN4_bit => VN_data_out(8170),
        VN2CN5_bit => VN_data_out(8171),
        VN2CN0_sign => VN_sign_out(8166),
        VN2CN1_sign => VN_sign_out(8167),
        VN2CN2_sign => VN_sign_out(8168),
        VN2CN3_sign => VN_sign_out(8169),
        VN2CN4_sign => VN_sign_out(8170),
        VN2CN5_sign => VN_sign_out(8171),
        codeword => codeword(1361),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1362 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8177 downto 8172),
        Din0 => VN1362_in0,
        Din1 => VN1362_in1,
        Din2 => VN1362_in2,
        Din3 => VN1362_in3,
        Din4 => VN1362_in4,
        Din5 => VN1362_in5,
        VN2CN0_bit => VN_data_out(8172),
        VN2CN1_bit => VN_data_out(8173),
        VN2CN2_bit => VN_data_out(8174),
        VN2CN3_bit => VN_data_out(8175),
        VN2CN4_bit => VN_data_out(8176),
        VN2CN5_bit => VN_data_out(8177),
        VN2CN0_sign => VN_sign_out(8172),
        VN2CN1_sign => VN_sign_out(8173),
        VN2CN2_sign => VN_sign_out(8174),
        VN2CN3_sign => VN_sign_out(8175),
        VN2CN4_sign => VN_sign_out(8176),
        VN2CN5_sign => VN_sign_out(8177),
        codeword => codeword(1362),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1363 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8183 downto 8178),
        Din0 => VN1363_in0,
        Din1 => VN1363_in1,
        Din2 => VN1363_in2,
        Din3 => VN1363_in3,
        Din4 => VN1363_in4,
        Din5 => VN1363_in5,
        VN2CN0_bit => VN_data_out(8178),
        VN2CN1_bit => VN_data_out(8179),
        VN2CN2_bit => VN_data_out(8180),
        VN2CN3_bit => VN_data_out(8181),
        VN2CN4_bit => VN_data_out(8182),
        VN2CN5_bit => VN_data_out(8183),
        VN2CN0_sign => VN_sign_out(8178),
        VN2CN1_sign => VN_sign_out(8179),
        VN2CN2_sign => VN_sign_out(8180),
        VN2CN3_sign => VN_sign_out(8181),
        VN2CN4_sign => VN_sign_out(8182),
        VN2CN5_sign => VN_sign_out(8183),
        codeword => codeword(1363),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1364 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8189 downto 8184),
        Din0 => VN1364_in0,
        Din1 => VN1364_in1,
        Din2 => VN1364_in2,
        Din3 => VN1364_in3,
        Din4 => VN1364_in4,
        Din5 => VN1364_in5,
        VN2CN0_bit => VN_data_out(8184),
        VN2CN1_bit => VN_data_out(8185),
        VN2CN2_bit => VN_data_out(8186),
        VN2CN3_bit => VN_data_out(8187),
        VN2CN4_bit => VN_data_out(8188),
        VN2CN5_bit => VN_data_out(8189),
        VN2CN0_sign => VN_sign_out(8184),
        VN2CN1_sign => VN_sign_out(8185),
        VN2CN2_sign => VN_sign_out(8186),
        VN2CN3_sign => VN_sign_out(8187),
        VN2CN4_sign => VN_sign_out(8188),
        VN2CN5_sign => VN_sign_out(8189),
        codeword => codeword(1364),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1365 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8195 downto 8190),
        Din0 => VN1365_in0,
        Din1 => VN1365_in1,
        Din2 => VN1365_in2,
        Din3 => VN1365_in3,
        Din4 => VN1365_in4,
        Din5 => VN1365_in5,
        VN2CN0_bit => VN_data_out(8190),
        VN2CN1_bit => VN_data_out(8191),
        VN2CN2_bit => VN_data_out(8192),
        VN2CN3_bit => VN_data_out(8193),
        VN2CN4_bit => VN_data_out(8194),
        VN2CN5_bit => VN_data_out(8195),
        VN2CN0_sign => VN_sign_out(8190),
        VN2CN1_sign => VN_sign_out(8191),
        VN2CN2_sign => VN_sign_out(8192),
        VN2CN3_sign => VN_sign_out(8193),
        VN2CN4_sign => VN_sign_out(8194),
        VN2CN5_sign => VN_sign_out(8195),
        codeword => codeword(1365),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1366 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8201 downto 8196),
        Din0 => VN1366_in0,
        Din1 => VN1366_in1,
        Din2 => VN1366_in2,
        Din3 => VN1366_in3,
        Din4 => VN1366_in4,
        Din5 => VN1366_in5,
        VN2CN0_bit => VN_data_out(8196),
        VN2CN1_bit => VN_data_out(8197),
        VN2CN2_bit => VN_data_out(8198),
        VN2CN3_bit => VN_data_out(8199),
        VN2CN4_bit => VN_data_out(8200),
        VN2CN5_bit => VN_data_out(8201),
        VN2CN0_sign => VN_sign_out(8196),
        VN2CN1_sign => VN_sign_out(8197),
        VN2CN2_sign => VN_sign_out(8198),
        VN2CN3_sign => VN_sign_out(8199),
        VN2CN4_sign => VN_sign_out(8200),
        VN2CN5_sign => VN_sign_out(8201),
        codeword => codeword(1366),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1367 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8207 downto 8202),
        Din0 => VN1367_in0,
        Din1 => VN1367_in1,
        Din2 => VN1367_in2,
        Din3 => VN1367_in3,
        Din4 => VN1367_in4,
        Din5 => VN1367_in5,
        VN2CN0_bit => VN_data_out(8202),
        VN2CN1_bit => VN_data_out(8203),
        VN2CN2_bit => VN_data_out(8204),
        VN2CN3_bit => VN_data_out(8205),
        VN2CN4_bit => VN_data_out(8206),
        VN2CN5_bit => VN_data_out(8207),
        VN2CN0_sign => VN_sign_out(8202),
        VN2CN1_sign => VN_sign_out(8203),
        VN2CN2_sign => VN_sign_out(8204),
        VN2CN3_sign => VN_sign_out(8205),
        VN2CN4_sign => VN_sign_out(8206),
        VN2CN5_sign => VN_sign_out(8207),
        codeword => codeword(1367),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1368 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8213 downto 8208),
        Din0 => VN1368_in0,
        Din1 => VN1368_in1,
        Din2 => VN1368_in2,
        Din3 => VN1368_in3,
        Din4 => VN1368_in4,
        Din5 => VN1368_in5,
        VN2CN0_bit => VN_data_out(8208),
        VN2CN1_bit => VN_data_out(8209),
        VN2CN2_bit => VN_data_out(8210),
        VN2CN3_bit => VN_data_out(8211),
        VN2CN4_bit => VN_data_out(8212),
        VN2CN5_bit => VN_data_out(8213),
        VN2CN0_sign => VN_sign_out(8208),
        VN2CN1_sign => VN_sign_out(8209),
        VN2CN2_sign => VN_sign_out(8210),
        VN2CN3_sign => VN_sign_out(8211),
        VN2CN4_sign => VN_sign_out(8212),
        VN2CN5_sign => VN_sign_out(8213),
        codeword => codeword(1368),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1369 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8219 downto 8214),
        Din0 => VN1369_in0,
        Din1 => VN1369_in1,
        Din2 => VN1369_in2,
        Din3 => VN1369_in3,
        Din4 => VN1369_in4,
        Din5 => VN1369_in5,
        VN2CN0_bit => VN_data_out(8214),
        VN2CN1_bit => VN_data_out(8215),
        VN2CN2_bit => VN_data_out(8216),
        VN2CN3_bit => VN_data_out(8217),
        VN2CN4_bit => VN_data_out(8218),
        VN2CN5_bit => VN_data_out(8219),
        VN2CN0_sign => VN_sign_out(8214),
        VN2CN1_sign => VN_sign_out(8215),
        VN2CN2_sign => VN_sign_out(8216),
        VN2CN3_sign => VN_sign_out(8217),
        VN2CN4_sign => VN_sign_out(8218),
        VN2CN5_sign => VN_sign_out(8219),
        codeword => codeword(1369),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1370 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8225 downto 8220),
        Din0 => VN1370_in0,
        Din1 => VN1370_in1,
        Din2 => VN1370_in2,
        Din3 => VN1370_in3,
        Din4 => VN1370_in4,
        Din5 => VN1370_in5,
        VN2CN0_bit => VN_data_out(8220),
        VN2CN1_bit => VN_data_out(8221),
        VN2CN2_bit => VN_data_out(8222),
        VN2CN3_bit => VN_data_out(8223),
        VN2CN4_bit => VN_data_out(8224),
        VN2CN5_bit => VN_data_out(8225),
        VN2CN0_sign => VN_sign_out(8220),
        VN2CN1_sign => VN_sign_out(8221),
        VN2CN2_sign => VN_sign_out(8222),
        VN2CN3_sign => VN_sign_out(8223),
        VN2CN4_sign => VN_sign_out(8224),
        VN2CN5_sign => VN_sign_out(8225),
        codeword => codeword(1370),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1371 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8231 downto 8226),
        Din0 => VN1371_in0,
        Din1 => VN1371_in1,
        Din2 => VN1371_in2,
        Din3 => VN1371_in3,
        Din4 => VN1371_in4,
        Din5 => VN1371_in5,
        VN2CN0_bit => VN_data_out(8226),
        VN2CN1_bit => VN_data_out(8227),
        VN2CN2_bit => VN_data_out(8228),
        VN2CN3_bit => VN_data_out(8229),
        VN2CN4_bit => VN_data_out(8230),
        VN2CN5_bit => VN_data_out(8231),
        VN2CN0_sign => VN_sign_out(8226),
        VN2CN1_sign => VN_sign_out(8227),
        VN2CN2_sign => VN_sign_out(8228),
        VN2CN3_sign => VN_sign_out(8229),
        VN2CN4_sign => VN_sign_out(8230),
        VN2CN5_sign => VN_sign_out(8231),
        codeword => codeword(1371),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1372 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8237 downto 8232),
        Din0 => VN1372_in0,
        Din1 => VN1372_in1,
        Din2 => VN1372_in2,
        Din3 => VN1372_in3,
        Din4 => VN1372_in4,
        Din5 => VN1372_in5,
        VN2CN0_bit => VN_data_out(8232),
        VN2CN1_bit => VN_data_out(8233),
        VN2CN2_bit => VN_data_out(8234),
        VN2CN3_bit => VN_data_out(8235),
        VN2CN4_bit => VN_data_out(8236),
        VN2CN5_bit => VN_data_out(8237),
        VN2CN0_sign => VN_sign_out(8232),
        VN2CN1_sign => VN_sign_out(8233),
        VN2CN2_sign => VN_sign_out(8234),
        VN2CN3_sign => VN_sign_out(8235),
        VN2CN4_sign => VN_sign_out(8236),
        VN2CN5_sign => VN_sign_out(8237),
        codeword => codeword(1372),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1373 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8243 downto 8238),
        Din0 => VN1373_in0,
        Din1 => VN1373_in1,
        Din2 => VN1373_in2,
        Din3 => VN1373_in3,
        Din4 => VN1373_in4,
        Din5 => VN1373_in5,
        VN2CN0_bit => VN_data_out(8238),
        VN2CN1_bit => VN_data_out(8239),
        VN2CN2_bit => VN_data_out(8240),
        VN2CN3_bit => VN_data_out(8241),
        VN2CN4_bit => VN_data_out(8242),
        VN2CN5_bit => VN_data_out(8243),
        VN2CN0_sign => VN_sign_out(8238),
        VN2CN1_sign => VN_sign_out(8239),
        VN2CN2_sign => VN_sign_out(8240),
        VN2CN3_sign => VN_sign_out(8241),
        VN2CN4_sign => VN_sign_out(8242),
        VN2CN5_sign => VN_sign_out(8243),
        codeword => codeword(1373),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1374 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8249 downto 8244),
        Din0 => VN1374_in0,
        Din1 => VN1374_in1,
        Din2 => VN1374_in2,
        Din3 => VN1374_in3,
        Din4 => VN1374_in4,
        Din5 => VN1374_in5,
        VN2CN0_bit => VN_data_out(8244),
        VN2CN1_bit => VN_data_out(8245),
        VN2CN2_bit => VN_data_out(8246),
        VN2CN3_bit => VN_data_out(8247),
        VN2CN4_bit => VN_data_out(8248),
        VN2CN5_bit => VN_data_out(8249),
        VN2CN0_sign => VN_sign_out(8244),
        VN2CN1_sign => VN_sign_out(8245),
        VN2CN2_sign => VN_sign_out(8246),
        VN2CN3_sign => VN_sign_out(8247),
        VN2CN4_sign => VN_sign_out(8248),
        VN2CN5_sign => VN_sign_out(8249),
        codeword => codeword(1374),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1375 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8255 downto 8250),
        Din0 => VN1375_in0,
        Din1 => VN1375_in1,
        Din2 => VN1375_in2,
        Din3 => VN1375_in3,
        Din4 => VN1375_in4,
        Din5 => VN1375_in5,
        VN2CN0_bit => VN_data_out(8250),
        VN2CN1_bit => VN_data_out(8251),
        VN2CN2_bit => VN_data_out(8252),
        VN2CN3_bit => VN_data_out(8253),
        VN2CN4_bit => VN_data_out(8254),
        VN2CN5_bit => VN_data_out(8255),
        VN2CN0_sign => VN_sign_out(8250),
        VN2CN1_sign => VN_sign_out(8251),
        VN2CN2_sign => VN_sign_out(8252),
        VN2CN3_sign => VN_sign_out(8253),
        VN2CN4_sign => VN_sign_out(8254),
        VN2CN5_sign => VN_sign_out(8255),
        codeword => codeword(1375),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1376 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8261 downto 8256),
        Din0 => VN1376_in0,
        Din1 => VN1376_in1,
        Din2 => VN1376_in2,
        Din3 => VN1376_in3,
        Din4 => VN1376_in4,
        Din5 => VN1376_in5,
        VN2CN0_bit => VN_data_out(8256),
        VN2CN1_bit => VN_data_out(8257),
        VN2CN2_bit => VN_data_out(8258),
        VN2CN3_bit => VN_data_out(8259),
        VN2CN4_bit => VN_data_out(8260),
        VN2CN5_bit => VN_data_out(8261),
        VN2CN0_sign => VN_sign_out(8256),
        VN2CN1_sign => VN_sign_out(8257),
        VN2CN2_sign => VN_sign_out(8258),
        VN2CN3_sign => VN_sign_out(8259),
        VN2CN4_sign => VN_sign_out(8260),
        VN2CN5_sign => VN_sign_out(8261),
        codeword => codeword(1376),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1377 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8267 downto 8262),
        Din0 => VN1377_in0,
        Din1 => VN1377_in1,
        Din2 => VN1377_in2,
        Din3 => VN1377_in3,
        Din4 => VN1377_in4,
        Din5 => VN1377_in5,
        VN2CN0_bit => VN_data_out(8262),
        VN2CN1_bit => VN_data_out(8263),
        VN2CN2_bit => VN_data_out(8264),
        VN2CN3_bit => VN_data_out(8265),
        VN2CN4_bit => VN_data_out(8266),
        VN2CN5_bit => VN_data_out(8267),
        VN2CN0_sign => VN_sign_out(8262),
        VN2CN1_sign => VN_sign_out(8263),
        VN2CN2_sign => VN_sign_out(8264),
        VN2CN3_sign => VN_sign_out(8265),
        VN2CN4_sign => VN_sign_out(8266),
        VN2CN5_sign => VN_sign_out(8267),
        codeword => codeword(1377),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1378 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8273 downto 8268),
        Din0 => VN1378_in0,
        Din1 => VN1378_in1,
        Din2 => VN1378_in2,
        Din3 => VN1378_in3,
        Din4 => VN1378_in4,
        Din5 => VN1378_in5,
        VN2CN0_bit => VN_data_out(8268),
        VN2CN1_bit => VN_data_out(8269),
        VN2CN2_bit => VN_data_out(8270),
        VN2CN3_bit => VN_data_out(8271),
        VN2CN4_bit => VN_data_out(8272),
        VN2CN5_bit => VN_data_out(8273),
        VN2CN0_sign => VN_sign_out(8268),
        VN2CN1_sign => VN_sign_out(8269),
        VN2CN2_sign => VN_sign_out(8270),
        VN2CN3_sign => VN_sign_out(8271),
        VN2CN4_sign => VN_sign_out(8272),
        VN2CN5_sign => VN_sign_out(8273),
        codeword => codeword(1378),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1379 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8279 downto 8274),
        Din0 => VN1379_in0,
        Din1 => VN1379_in1,
        Din2 => VN1379_in2,
        Din3 => VN1379_in3,
        Din4 => VN1379_in4,
        Din5 => VN1379_in5,
        VN2CN0_bit => VN_data_out(8274),
        VN2CN1_bit => VN_data_out(8275),
        VN2CN2_bit => VN_data_out(8276),
        VN2CN3_bit => VN_data_out(8277),
        VN2CN4_bit => VN_data_out(8278),
        VN2CN5_bit => VN_data_out(8279),
        VN2CN0_sign => VN_sign_out(8274),
        VN2CN1_sign => VN_sign_out(8275),
        VN2CN2_sign => VN_sign_out(8276),
        VN2CN3_sign => VN_sign_out(8277),
        VN2CN4_sign => VN_sign_out(8278),
        VN2CN5_sign => VN_sign_out(8279),
        codeword => codeword(1379),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1380 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8285 downto 8280),
        Din0 => VN1380_in0,
        Din1 => VN1380_in1,
        Din2 => VN1380_in2,
        Din3 => VN1380_in3,
        Din4 => VN1380_in4,
        Din5 => VN1380_in5,
        VN2CN0_bit => VN_data_out(8280),
        VN2CN1_bit => VN_data_out(8281),
        VN2CN2_bit => VN_data_out(8282),
        VN2CN3_bit => VN_data_out(8283),
        VN2CN4_bit => VN_data_out(8284),
        VN2CN5_bit => VN_data_out(8285),
        VN2CN0_sign => VN_sign_out(8280),
        VN2CN1_sign => VN_sign_out(8281),
        VN2CN2_sign => VN_sign_out(8282),
        VN2CN3_sign => VN_sign_out(8283),
        VN2CN4_sign => VN_sign_out(8284),
        VN2CN5_sign => VN_sign_out(8285),
        codeword => codeword(1380),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1381 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8291 downto 8286),
        Din0 => VN1381_in0,
        Din1 => VN1381_in1,
        Din2 => VN1381_in2,
        Din3 => VN1381_in3,
        Din4 => VN1381_in4,
        Din5 => VN1381_in5,
        VN2CN0_bit => VN_data_out(8286),
        VN2CN1_bit => VN_data_out(8287),
        VN2CN2_bit => VN_data_out(8288),
        VN2CN3_bit => VN_data_out(8289),
        VN2CN4_bit => VN_data_out(8290),
        VN2CN5_bit => VN_data_out(8291),
        VN2CN0_sign => VN_sign_out(8286),
        VN2CN1_sign => VN_sign_out(8287),
        VN2CN2_sign => VN_sign_out(8288),
        VN2CN3_sign => VN_sign_out(8289),
        VN2CN4_sign => VN_sign_out(8290),
        VN2CN5_sign => VN_sign_out(8291),
        codeword => codeword(1381),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1382 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8297 downto 8292),
        Din0 => VN1382_in0,
        Din1 => VN1382_in1,
        Din2 => VN1382_in2,
        Din3 => VN1382_in3,
        Din4 => VN1382_in4,
        Din5 => VN1382_in5,
        VN2CN0_bit => VN_data_out(8292),
        VN2CN1_bit => VN_data_out(8293),
        VN2CN2_bit => VN_data_out(8294),
        VN2CN3_bit => VN_data_out(8295),
        VN2CN4_bit => VN_data_out(8296),
        VN2CN5_bit => VN_data_out(8297),
        VN2CN0_sign => VN_sign_out(8292),
        VN2CN1_sign => VN_sign_out(8293),
        VN2CN2_sign => VN_sign_out(8294),
        VN2CN3_sign => VN_sign_out(8295),
        VN2CN4_sign => VN_sign_out(8296),
        VN2CN5_sign => VN_sign_out(8297),
        codeword => codeword(1382),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1383 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8303 downto 8298),
        Din0 => VN1383_in0,
        Din1 => VN1383_in1,
        Din2 => VN1383_in2,
        Din3 => VN1383_in3,
        Din4 => VN1383_in4,
        Din5 => VN1383_in5,
        VN2CN0_bit => VN_data_out(8298),
        VN2CN1_bit => VN_data_out(8299),
        VN2CN2_bit => VN_data_out(8300),
        VN2CN3_bit => VN_data_out(8301),
        VN2CN4_bit => VN_data_out(8302),
        VN2CN5_bit => VN_data_out(8303),
        VN2CN0_sign => VN_sign_out(8298),
        VN2CN1_sign => VN_sign_out(8299),
        VN2CN2_sign => VN_sign_out(8300),
        VN2CN3_sign => VN_sign_out(8301),
        VN2CN4_sign => VN_sign_out(8302),
        VN2CN5_sign => VN_sign_out(8303),
        codeword => codeword(1383),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1384 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8309 downto 8304),
        Din0 => VN1384_in0,
        Din1 => VN1384_in1,
        Din2 => VN1384_in2,
        Din3 => VN1384_in3,
        Din4 => VN1384_in4,
        Din5 => VN1384_in5,
        VN2CN0_bit => VN_data_out(8304),
        VN2CN1_bit => VN_data_out(8305),
        VN2CN2_bit => VN_data_out(8306),
        VN2CN3_bit => VN_data_out(8307),
        VN2CN4_bit => VN_data_out(8308),
        VN2CN5_bit => VN_data_out(8309),
        VN2CN0_sign => VN_sign_out(8304),
        VN2CN1_sign => VN_sign_out(8305),
        VN2CN2_sign => VN_sign_out(8306),
        VN2CN3_sign => VN_sign_out(8307),
        VN2CN4_sign => VN_sign_out(8308),
        VN2CN5_sign => VN_sign_out(8309),
        codeword => codeword(1384),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1385 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8315 downto 8310),
        Din0 => VN1385_in0,
        Din1 => VN1385_in1,
        Din2 => VN1385_in2,
        Din3 => VN1385_in3,
        Din4 => VN1385_in4,
        Din5 => VN1385_in5,
        VN2CN0_bit => VN_data_out(8310),
        VN2CN1_bit => VN_data_out(8311),
        VN2CN2_bit => VN_data_out(8312),
        VN2CN3_bit => VN_data_out(8313),
        VN2CN4_bit => VN_data_out(8314),
        VN2CN5_bit => VN_data_out(8315),
        VN2CN0_sign => VN_sign_out(8310),
        VN2CN1_sign => VN_sign_out(8311),
        VN2CN2_sign => VN_sign_out(8312),
        VN2CN3_sign => VN_sign_out(8313),
        VN2CN4_sign => VN_sign_out(8314),
        VN2CN5_sign => VN_sign_out(8315),
        codeword => codeword(1385),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1386 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8321 downto 8316),
        Din0 => VN1386_in0,
        Din1 => VN1386_in1,
        Din2 => VN1386_in2,
        Din3 => VN1386_in3,
        Din4 => VN1386_in4,
        Din5 => VN1386_in5,
        VN2CN0_bit => VN_data_out(8316),
        VN2CN1_bit => VN_data_out(8317),
        VN2CN2_bit => VN_data_out(8318),
        VN2CN3_bit => VN_data_out(8319),
        VN2CN4_bit => VN_data_out(8320),
        VN2CN5_bit => VN_data_out(8321),
        VN2CN0_sign => VN_sign_out(8316),
        VN2CN1_sign => VN_sign_out(8317),
        VN2CN2_sign => VN_sign_out(8318),
        VN2CN3_sign => VN_sign_out(8319),
        VN2CN4_sign => VN_sign_out(8320),
        VN2CN5_sign => VN_sign_out(8321),
        codeword => codeword(1386),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1387 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8327 downto 8322),
        Din0 => VN1387_in0,
        Din1 => VN1387_in1,
        Din2 => VN1387_in2,
        Din3 => VN1387_in3,
        Din4 => VN1387_in4,
        Din5 => VN1387_in5,
        VN2CN0_bit => VN_data_out(8322),
        VN2CN1_bit => VN_data_out(8323),
        VN2CN2_bit => VN_data_out(8324),
        VN2CN3_bit => VN_data_out(8325),
        VN2CN4_bit => VN_data_out(8326),
        VN2CN5_bit => VN_data_out(8327),
        VN2CN0_sign => VN_sign_out(8322),
        VN2CN1_sign => VN_sign_out(8323),
        VN2CN2_sign => VN_sign_out(8324),
        VN2CN3_sign => VN_sign_out(8325),
        VN2CN4_sign => VN_sign_out(8326),
        VN2CN5_sign => VN_sign_out(8327),
        codeword => codeword(1387),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1388 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8333 downto 8328),
        Din0 => VN1388_in0,
        Din1 => VN1388_in1,
        Din2 => VN1388_in2,
        Din3 => VN1388_in3,
        Din4 => VN1388_in4,
        Din5 => VN1388_in5,
        VN2CN0_bit => VN_data_out(8328),
        VN2CN1_bit => VN_data_out(8329),
        VN2CN2_bit => VN_data_out(8330),
        VN2CN3_bit => VN_data_out(8331),
        VN2CN4_bit => VN_data_out(8332),
        VN2CN5_bit => VN_data_out(8333),
        VN2CN0_sign => VN_sign_out(8328),
        VN2CN1_sign => VN_sign_out(8329),
        VN2CN2_sign => VN_sign_out(8330),
        VN2CN3_sign => VN_sign_out(8331),
        VN2CN4_sign => VN_sign_out(8332),
        VN2CN5_sign => VN_sign_out(8333),
        codeword => codeword(1388),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1389 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8339 downto 8334),
        Din0 => VN1389_in0,
        Din1 => VN1389_in1,
        Din2 => VN1389_in2,
        Din3 => VN1389_in3,
        Din4 => VN1389_in4,
        Din5 => VN1389_in5,
        VN2CN0_bit => VN_data_out(8334),
        VN2CN1_bit => VN_data_out(8335),
        VN2CN2_bit => VN_data_out(8336),
        VN2CN3_bit => VN_data_out(8337),
        VN2CN4_bit => VN_data_out(8338),
        VN2CN5_bit => VN_data_out(8339),
        VN2CN0_sign => VN_sign_out(8334),
        VN2CN1_sign => VN_sign_out(8335),
        VN2CN2_sign => VN_sign_out(8336),
        VN2CN3_sign => VN_sign_out(8337),
        VN2CN4_sign => VN_sign_out(8338),
        VN2CN5_sign => VN_sign_out(8339),
        codeword => codeword(1389),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1390 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8345 downto 8340),
        Din0 => VN1390_in0,
        Din1 => VN1390_in1,
        Din2 => VN1390_in2,
        Din3 => VN1390_in3,
        Din4 => VN1390_in4,
        Din5 => VN1390_in5,
        VN2CN0_bit => VN_data_out(8340),
        VN2CN1_bit => VN_data_out(8341),
        VN2CN2_bit => VN_data_out(8342),
        VN2CN3_bit => VN_data_out(8343),
        VN2CN4_bit => VN_data_out(8344),
        VN2CN5_bit => VN_data_out(8345),
        VN2CN0_sign => VN_sign_out(8340),
        VN2CN1_sign => VN_sign_out(8341),
        VN2CN2_sign => VN_sign_out(8342),
        VN2CN3_sign => VN_sign_out(8343),
        VN2CN4_sign => VN_sign_out(8344),
        VN2CN5_sign => VN_sign_out(8345),
        codeword => codeword(1390),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1391 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8351 downto 8346),
        Din0 => VN1391_in0,
        Din1 => VN1391_in1,
        Din2 => VN1391_in2,
        Din3 => VN1391_in3,
        Din4 => VN1391_in4,
        Din5 => VN1391_in5,
        VN2CN0_bit => VN_data_out(8346),
        VN2CN1_bit => VN_data_out(8347),
        VN2CN2_bit => VN_data_out(8348),
        VN2CN3_bit => VN_data_out(8349),
        VN2CN4_bit => VN_data_out(8350),
        VN2CN5_bit => VN_data_out(8351),
        VN2CN0_sign => VN_sign_out(8346),
        VN2CN1_sign => VN_sign_out(8347),
        VN2CN2_sign => VN_sign_out(8348),
        VN2CN3_sign => VN_sign_out(8349),
        VN2CN4_sign => VN_sign_out(8350),
        VN2CN5_sign => VN_sign_out(8351),
        codeword => codeword(1391),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1392 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8357 downto 8352),
        Din0 => VN1392_in0,
        Din1 => VN1392_in1,
        Din2 => VN1392_in2,
        Din3 => VN1392_in3,
        Din4 => VN1392_in4,
        Din5 => VN1392_in5,
        VN2CN0_bit => VN_data_out(8352),
        VN2CN1_bit => VN_data_out(8353),
        VN2CN2_bit => VN_data_out(8354),
        VN2CN3_bit => VN_data_out(8355),
        VN2CN4_bit => VN_data_out(8356),
        VN2CN5_bit => VN_data_out(8357),
        VN2CN0_sign => VN_sign_out(8352),
        VN2CN1_sign => VN_sign_out(8353),
        VN2CN2_sign => VN_sign_out(8354),
        VN2CN3_sign => VN_sign_out(8355),
        VN2CN4_sign => VN_sign_out(8356),
        VN2CN5_sign => VN_sign_out(8357),
        codeword => codeword(1392),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1393 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8363 downto 8358),
        Din0 => VN1393_in0,
        Din1 => VN1393_in1,
        Din2 => VN1393_in2,
        Din3 => VN1393_in3,
        Din4 => VN1393_in4,
        Din5 => VN1393_in5,
        VN2CN0_bit => VN_data_out(8358),
        VN2CN1_bit => VN_data_out(8359),
        VN2CN2_bit => VN_data_out(8360),
        VN2CN3_bit => VN_data_out(8361),
        VN2CN4_bit => VN_data_out(8362),
        VN2CN5_bit => VN_data_out(8363),
        VN2CN0_sign => VN_sign_out(8358),
        VN2CN1_sign => VN_sign_out(8359),
        VN2CN2_sign => VN_sign_out(8360),
        VN2CN3_sign => VN_sign_out(8361),
        VN2CN4_sign => VN_sign_out(8362),
        VN2CN5_sign => VN_sign_out(8363),
        codeword => codeword(1393),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1394 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8369 downto 8364),
        Din0 => VN1394_in0,
        Din1 => VN1394_in1,
        Din2 => VN1394_in2,
        Din3 => VN1394_in3,
        Din4 => VN1394_in4,
        Din5 => VN1394_in5,
        VN2CN0_bit => VN_data_out(8364),
        VN2CN1_bit => VN_data_out(8365),
        VN2CN2_bit => VN_data_out(8366),
        VN2CN3_bit => VN_data_out(8367),
        VN2CN4_bit => VN_data_out(8368),
        VN2CN5_bit => VN_data_out(8369),
        VN2CN0_sign => VN_sign_out(8364),
        VN2CN1_sign => VN_sign_out(8365),
        VN2CN2_sign => VN_sign_out(8366),
        VN2CN3_sign => VN_sign_out(8367),
        VN2CN4_sign => VN_sign_out(8368),
        VN2CN5_sign => VN_sign_out(8369),
        codeword => codeword(1394),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1395 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8375 downto 8370),
        Din0 => VN1395_in0,
        Din1 => VN1395_in1,
        Din2 => VN1395_in2,
        Din3 => VN1395_in3,
        Din4 => VN1395_in4,
        Din5 => VN1395_in5,
        VN2CN0_bit => VN_data_out(8370),
        VN2CN1_bit => VN_data_out(8371),
        VN2CN2_bit => VN_data_out(8372),
        VN2CN3_bit => VN_data_out(8373),
        VN2CN4_bit => VN_data_out(8374),
        VN2CN5_bit => VN_data_out(8375),
        VN2CN0_sign => VN_sign_out(8370),
        VN2CN1_sign => VN_sign_out(8371),
        VN2CN2_sign => VN_sign_out(8372),
        VN2CN3_sign => VN_sign_out(8373),
        VN2CN4_sign => VN_sign_out(8374),
        VN2CN5_sign => VN_sign_out(8375),
        codeword => codeword(1395),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1396 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8381 downto 8376),
        Din0 => VN1396_in0,
        Din1 => VN1396_in1,
        Din2 => VN1396_in2,
        Din3 => VN1396_in3,
        Din4 => VN1396_in4,
        Din5 => VN1396_in5,
        VN2CN0_bit => VN_data_out(8376),
        VN2CN1_bit => VN_data_out(8377),
        VN2CN2_bit => VN_data_out(8378),
        VN2CN3_bit => VN_data_out(8379),
        VN2CN4_bit => VN_data_out(8380),
        VN2CN5_bit => VN_data_out(8381),
        VN2CN0_sign => VN_sign_out(8376),
        VN2CN1_sign => VN_sign_out(8377),
        VN2CN2_sign => VN_sign_out(8378),
        VN2CN3_sign => VN_sign_out(8379),
        VN2CN4_sign => VN_sign_out(8380),
        VN2CN5_sign => VN_sign_out(8381),
        codeword => codeword(1396),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1397 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8387 downto 8382),
        Din0 => VN1397_in0,
        Din1 => VN1397_in1,
        Din2 => VN1397_in2,
        Din3 => VN1397_in3,
        Din4 => VN1397_in4,
        Din5 => VN1397_in5,
        VN2CN0_bit => VN_data_out(8382),
        VN2CN1_bit => VN_data_out(8383),
        VN2CN2_bit => VN_data_out(8384),
        VN2CN3_bit => VN_data_out(8385),
        VN2CN4_bit => VN_data_out(8386),
        VN2CN5_bit => VN_data_out(8387),
        VN2CN0_sign => VN_sign_out(8382),
        VN2CN1_sign => VN_sign_out(8383),
        VN2CN2_sign => VN_sign_out(8384),
        VN2CN3_sign => VN_sign_out(8385),
        VN2CN4_sign => VN_sign_out(8386),
        VN2CN5_sign => VN_sign_out(8387),
        codeword => codeword(1397),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1398 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8393 downto 8388),
        Din0 => VN1398_in0,
        Din1 => VN1398_in1,
        Din2 => VN1398_in2,
        Din3 => VN1398_in3,
        Din4 => VN1398_in4,
        Din5 => VN1398_in5,
        VN2CN0_bit => VN_data_out(8388),
        VN2CN1_bit => VN_data_out(8389),
        VN2CN2_bit => VN_data_out(8390),
        VN2CN3_bit => VN_data_out(8391),
        VN2CN4_bit => VN_data_out(8392),
        VN2CN5_bit => VN_data_out(8393),
        VN2CN0_sign => VN_sign_out(8388),
        VN2CN1_sign => VN_sign_out(8389),
        VN2CN2_sign => VN_sign_out(8390),
        VN2CN3_sign => VN_sign_out(8391),
        VN2CN4_sign => VN_sign_out(8392),
        VN2CN5_sign => VN_sign_out(8393),
        codeword => codeword(1398),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1399 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8399 downto 8394),
        Din0 => VN1399_in0,
        Din1 => VN1399_in1,
        Din2 => VN1399_in2,
        Din3 => VN1399_in3,
        Din4 => VN1399_in4,
        Din5 => VN1399_in5,
        VN2CN0_bit => VN_data_out(8394),
        VN2CN1_bit => VN_data_out(8395),
        VN2CN2_bit => VN_data_out(8396),
        VN2CN3_bit => VN_data_out(8397),
        VN2CN4_bit => VN_data_out(8398),
        VN2CN5_bit => VN_data_out(8399),
        VN2CN0_sign => VN_sign_out(8394),
        VN2CN1_sign => VN_sign_out(8395),
        VN2CN2_sign => VN_sign_out(8396),
        VN2CN3_sign => VN_sign_out(8397),
        VN2CN4_sign => VN_sign_out(8398),
        VN2CN5_sign => VN_sign_out(8399),
        codeword => codeword(1399),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1400 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8405 downto 8400),
        Din0 => VN1400_in0,
        Din1 => VN1400_in1,
        Din2 => VN1400_in2,
        Din3 => VN1400_in3,
        Din4 => VN1400_in4,
        Din5 => VN1400_in5,
        VN2CN0_bit => VN_data_out(8400),
        VN2CN1_bit => VN_data_out(8401),
        VN2CN2_bit => VN_data_out(8402),
        VN2CN3_bit => VN_data_out(8403),
        VN2CN4_bit => VN_data_out(8404),
        VN2CN5_bit => VN_data_out(8405),
        VN2CN0_sign => VN_sign_out(8400),
        VN2CN1_sign => VN_sign_out(8401),
        VN2CN2_sign => VN_sign_out(8402),
        VN2CN3_sign => VN_sign_out(8403),
        VN2CN4_sign => VN_sign_out(8404),
        VN2CN5_sign => VN_sign_out(8405),
        codeword => codeword(1400),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1401 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8411 downto 8406),
        Din0 => VN1401_in0,
        Din1 => VN1401_in1,
        Din2 => VN1401_in2,
        Din3 => VN1401_in3,
        Din4 => VN1401_in4,
        Din5 => VN1401_in5,
        VN2CN0_bit => VN_data_out(8406),
        VN2CN1_bit => VN_data_out(8407),
        VN2CN2_bit => VN_data_out(8408),
        VN2CN3_bit => VN_data_out(8409),
        VN2CN4_bit => VN_data_out(8410),
        VN2CN5_bit => VN_data_out(8411),
        VN2CN0_sign => VN_sign_out(8406),
        VN2CN1_sign => VN_sign_out(8407),
        VN2CN2_sign => VN_sign_out(8408),
        VN2CN3_sign => VN_sign_out(8409),
        VN2CN4_sign => VN_sign_out(8410),
        VN2CN5_sign => VN_sign_out(8411),
        codeword => codeword(1401),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1402 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8417 downto 8412),
        Din0 => VN1402_in0,
        Din1 => VN1402_in1,
        Din2 => VN1402_in2,
        Din3 => VN1402_in3,
        Din4 => VN1402_in4,
        Din5 => VN1402_in5,
        VN2CN0_bit => VN_data_out(8412),
        VN2CN1_bit => VN_data_out(8413),
        VN2CN2_bit => VN_data_out(8414),
        VN2CN3_bit => VN_data_out(8415),
        VN2CN4_bit => VN_data_out(8416),
        VN2CN5_bit => VN_data_out(8417),
        VN2CN0_sign => VN_sign_out(8412),
        VN2CN1_sign => VN_sign_out(8413),
        VN2CN2_sign => VN_sign_out(8414),
        VN2CN3_sign => VN_sign_out(8415),
        VN2CN4_sign => VN_sign_out(8416),
        VN2CN5_sign => VN_sign_out(8417),
        codeword => codeword(1402),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1403 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8423 downto 8418),
        Din0 => VN1403_in0,
        Din1 => VN1403_in1,
        Din2 => VN1403_in2,
        Din3 => VN1403_in3,
        Din4 => VN1403_in4,
        Din5 => VN1403_in5,
        VN2CN0_bit => VN_data_out(8418),
        VN2CN1_bit => VN_data_out(8419),
        VN2CN2_bit => VN_data_out(8420),
        VN2CN3_bit => VN_data_out(8421),
        VN2CN4_bit => VN_data_out(8422),
        VN2CN5_bit => VN_data_out(8423),
        VN2CN0_sign => VN_sign_out(8418),
        VN2CN1_sign => VN_sign_out(8419),
        VN2CN2_sign => VN_sign_out(8420),
        VN2CN3_sign => VN_sign_out(8421),
        VN2CN4_sign => VN_sign_out(8422),
        VN2CN5_sign => VN_sign_out(8423),
        codeword => codeword(1403),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1404 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8429 downto 8424),
        Din0 => VN1404_in0,
        Din1 => VN1404_in1,
        Din2 => VN1404_in2,
        Din3 => VN1404_in3,
        Din4 => VN1404_in4,
        Din5 => VN1404_in5,
        VN2CN0_bit => VN_data_out(8424),
        VN2CN1_bit => VN_data_out(8425),
        VN2CN2_bit => VN_data_out(8426),
        VN2CN3_bit => VN_data_out(8427),
        VN2CN4_bit => VN_data_out(8428),
        VN2CN5_bit => VN_data_out(8429),
        VN2CN0_sign => VN_sign_out(8424),
        VN2CN1_sign => VN_sign_out(8425),
        VN2CN2_sign => VN_sign_out(8426),
        VN2CN3_sign => VN_sign_out(8427),
        VN2CN4_sign => VN_sign_out(8428),
        VN2CN5_sign => VN_sign_out(8429),
        codeword => codeword(1404),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1405 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8435 downto 8430),
        Din0 => VN1405_in0,
        Din1 => VN1405_in1,
        Din2 => VN1405_in2,
        Din3 => VN1405_in3,
        Din4 => VN1405_in4,
        Din5 => VN1405_in5,
        VN2CN0_bit => VN_data_out(8430),
        VN2CN1_bit => VN_data_out(8431),
        VN2CN2_bit => VN_data_out(8432),
        VN2CN3_bit => VN_data_out(8433),
        VN2CN4_bit => VN_data_out(8434),
        VN2CN5_bit => VN_data_out(8435),
        VN2CN0_sign => VN_sign_out(8430),
        VN2CN1_sign => VN_sign_out(8431),
        VN2CN2_sign => VN_sign_out(8432),
        VN2CN3_sign => VN_sign_out(8433),
        VN2CN4_sign => VN_sign_out(8434),
        VN2CN5_sign => VN_sign_out(8435),
        codeword => codeword(1405),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1406 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8441 downto 8436),
        Din0 => VN1406_in0,
        Din1 => VN1406_in1,
        Din2 => VN1406_in2,
        Din3 => VN1406_in3,
        Din4 => VN1406_in4,
        Din5 => VN1406_in5,
        VN2CN0_bit => VN_data_out(8436),
        VN2CN1_bit => VN_data_out(8437),
        VN2CN2_bit => VN_data_out(8438),
        VN2CN3_bit => VN_data_out(8439),
        VN2CN4_bit => VN_data_out(8440),
        VN2CN5_bit => VN_data_out(8441),
        VN2CN0_sign => VN_sign_out(8436),
        VN2CN1_sign => VN_sign_out(8437),
        VN2CN2_sign => VN_sign_out(8438),
        VN2CN3_sign => VN_sign_out(8439),
        VN2CN4_sign => VN_sign_out(8440),
        VN2CN5_sign => VN_sign_out(8441),
        codeword => codeword(1406),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1407 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8447 downto 8442),
        Din0 => VN1407_in0,
        Din1 => VN1407_in1,
        Din2 => VN1407_in2,
        Din3 => VN1407_in3,
        Din4 => VN1407_in4,
        Din5 => VN1407_in5,
        VN2CN0_bit => VN_data_out(8442),
        VN2CN1_bit => VN_data_out(8443),
        VN2CN2_bit => VN_data_out(8444),
        VN2CN3_bit => VN_data_out(8445),
        VN2CN4_bit => VN_data_out(8446),
        VN2CN5_bit => VN_data_out(8447),
        VN2CN0_sign => VN_sign_out(8442),
        VN2CN1_sign => VN_sign_out(8443),
        VN2CN2_sign => VN_sign_out(8444),
        VN2CN3_sign => VN_sign_out(8445),
        VN2CN4_sign => VN_sign_out(8446),
        VN2CN5_sign => VN_sign_out(8447),
        codeword => codeword(1407),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1408 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8453 downto 8448),
        Din0 => VN1408_in0,
        Din1 => VN1408_in1,
        Din2 => VN1408_in2,
        Din3 => VN1408_in3,
        Din4 => VN1408_in4,
        Din5 => VN1408_in5,
        VN2CN0_bit => VN_data_out(8448),
        VN2CN1_bit => VN_data_out(8449),
        VN2CN2_bit => VN_data_out(8450),
        VN2CN3_bit => VN_data_out(8451),
        VN2CN4_bit => VN_data_out(8452),
        VN2CN5_bit => VN_data_out(8453),
        VN2CN0_sign => VN_sign_out(8448),
        VN2CN1_sign => VN_sign_out(8449),
        VN2CN2_sign => VN_sign_out(8450),
        VN2CN3_sign => VN_sign_out(8451),
        VN2CN4_sign => VN_sign_out(8452),
        VN2CN5_sign => VN_sign_out(8453),
        codeword => codeword(1408),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1409 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8459 downto 8454),
        Din0 => VN1409_in0,
        Din1 => VN1409_in1,
        Din2 => VN1409_in2,
        Din3 => VN1409_in3,
        Din4 => VN1409_in4,
        Din5 => VN1409_in5,
        VN2CN0_bit => VN_data_out(8454),
        VN2CN1_bit => VN_data_out(8455),
        VN2CN2_bit => VN_data_out(8456),
        VN2CN3_bit => VN_data_out(8457),
        VN2CN4_bit => VN_data_out(8458),
        VN2CN5_bit => VN_data_out(8459),
        VN2CN0_sign => VN_sign_out(8454),
        VN2CN1_sign => VN_sign_out(8455),
        VN2CN2_sign => VN_sign_out(8456),
        VN2CN3_sign => VN_sign_out(8457),
        VN2CN4_sign => VN_sign_out(8458),
        VN2CN5_sign => VN_sign_out(8459),
        codeword => codeword(1409),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1410 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8465 downto 8460),
        Din0 => VN1410_in0,
        Din1 => VN1410_in1,
        Din2 => VN1410_in2,
        Din3 => VN1410_in3,
        Din4 => VN1410_in4,
        Din5 => VN1410_in5,
        VN2CN0_bit => VN_data_out(8460),
        VN2CN1_bit => VN_data_out(8461),
        VN2CN2_bit => VN_data_out(8462),
        VN2CN3_bit => VN_data_out(8463),
        VN2CN4_bit => VN_data_out(8464),
        VN2CN5_bit => VN_data_out(8465),
        VN2CN0_sign => VN_sign_out(8460),
        VN2CN1_sign => VN_sign_out(8461),
        VN2CN2_sign => VN_sign_out(8462),
        VN2CN3_sign => VN_sign_out(8463),
        VN2CN4_sign => VN_sign_out(8464),
        VN2CN5_sign => VN_sign_out(8465),
        codeword => codeword(1410),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1411 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8471 downto 8466),
        Din0 => VN1411_in0,
        Din1 => VN1411_in1,
        Din2 => VN1411_in2,
        Din3 => VN1411_in3,
        Din4 => VN1411_in4,
        Din5 => VN1411_in5,
        VN2CN0_bit => VN_data_out(8466),
        VN2CN1_bit => VN_data_out(8467),
        VN2CN2_bit => VN_data_out(8468),
        VN2CN3_bit => VN_data_out(8469),
        VN2CN4_bit => VN_data_out(8470),
        VN2CN5_bit => VN_data_out(8471),
        VN2CN0_sign => VN_sign_out(8466),
        VN2CN1_sign => VN_sign_out(8467),
        VN2CN2_sign => VN_sign_out(8468),
        VN2CN3_sign => VN_sign_out(8469),
        VN2CN4_sign => VN_sign_out(8470),
        VN2CN5_sign => VN_sign_out(8471),
        codeword => codeword(1411),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1412 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8477 downto 8472),
        Din0 => VN1412_in0,
        Din1 => VN1412_in1,
        Din2 => VN1412_in2,
        Din3 => VN1412_in3,
        Din4 => VN1412_in4,
        Din5 => VN1412_in5,
        VN2CN0_bit => VN_data_out(8472),
        VN2CN1_bit => VN_data_out(8473),
        VN2CN2_bit => VN_data_out(8474),
        VN2CN3_bit => VN_data_out(8475),
        VN2CN4_bit => VN_data_out(8476),
        VN2CN5_bit => VN_data_out(8477),
        VN2CN0_sign => VN_sign_out(8472),
        VN2CN1_sign => VN_sign_out(8473),
        VN2CN2_sign => VN_sign_out(8474),
        VN2CN3_sign => VN_sign_out(8475),
        VN2CN4_sign => VN_sign_out(8476),
        VN2CN5_sign => VN_sign_out(8477),
        codeword => codeword(1412),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1413 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8483 downto 8478),
        Din0 => VN1413_in0,
        Din1 => VN1413_in1,
        Din2 => VN1413_in2,
        Din3 => VN1413_in3,
        Din4 => VN1413_in4,
        Din5 => VN1413_in5,
        VN2CN0_bit => VN_data_out(8478),
        VN2CN1_bit => VN_data_out(8479),
        VN2CN2_bit => VN_data_out(8480),
        VN2CN3_bit => VN_data_out(8481),
        VN2CN4_bit => VN_data_out(8482),
        VN2CN5_bit => VN_data_out(8483),
        VN2CN0_sign => VN_sign_out(8478),
        VN2CN1_sign => VN_sign_out(8479),
        VN2CN2_sign => VN_sign_out(8480),
        VN2CN3_sign => VN_sign_out(8481),
        VN2CN4_sign => VN_sign_out(8482),
        VN2CN5_sign => VN_sign_out(8483),
        codeword => codeword(1413),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1414 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8489 downto 8484),
        Din0 => VN1414_in0,
        Din1 => VN1414_in1,
        Din2 => VN1414_in2,
        Din3 => VN1414_in3,
        Din4 => VN1414_in4,
        Din5 => VN1414_in5,
        VN2CN0_bit => VN_data_out(8484),
        VN2CN1_bit => VN_data_out(8485),
        VN2CN2_bit => VN_data_out(8486),
        VN2CN3_bit => VN_data_out(8487),
        VN2CN4_bit => VN_data_out(8488),
        VN2CN5_bit => VN_data_out(8489),
        VN2CN0_sign => VN_sign_out(8484),
        VN2CN1_sign => VN_sign_out(8485),
        VN2CN2_sign => VN_sign_out(8486),
        VN2CN3_sign => VN_sign_out(8487),
        VN2CN4_sign => VN_sign_out(8488),
        VN2CN5_sign => VN_sign_out(8489),
        codeword => codeword(1414),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1415 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8495 downto 8490),
        Din0 => VN1415_in0,
        Din1 => VN1415_in1,
        Din2 => VN1415_in2,
        Din3 => VN1415_in3,
        Din4 => VN1415_in4,
        Din5 => VN1415_in5,
        VN2CN0_bit => VN_data_out(8490),
        VN2CN1_bit => VN_data_out(8491),
        VN2CN2_bit => VN_data_out(8492),
        VN2CN3_bit => VN_data_out(8493),
        VN2CN4_bit => VN_data_out(8494),
        VN2CN5_bit => VN_data_out(8495),
        VN2CN0_sign => VN_sign_out(8490),
        VN2CN1_sign => VN_sign_out(8491),
        VN2CN2_sign => VN_sign_out(8492),
        VN2CN3_sign => VN_sign_out(8493),
        VN2CN4_sign => VN_sign_out(8494),
        VN2CN5_sign => VN_sign_out(8495),
        codeword => codeword(1415),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1416 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8501 downto 8496),
        Din0 => VN1416_in0,
        Din1 => VN1416_in1,
        Din2 => VN1416_in2,
        Din3 => VN1416_in3,
        Din4 => VN1416_in4,
        Din5 => VN1416_in5,
        VN2CN0_bit => VN_data_out(8496),
        VN2CN1_bit => VN_data_out(8497),
        VN2CN2_bit => VN_data_out(8498),
        VN2CN3_bit => VN_data_out(8499),
        VN2CN4_bit => VN_data_out(8500),
        VN2CN5_bit => VN_data_out(8501),
        VN2CN0_sign => VN_sign_out(8496),
        VN2CN1_sign => VN_sign_out(8497),
        VN2CN2_sign => VN_sign_out(8498),
        VN2CN3_sign => VN_sign_out(8499),
        VN2CN4_sign => VN_sign_out(8500),
        VN2CN5_sign => VN_sign_out(8501),
        codeword => codeword(1416),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1417 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8507 downto 8502),
        Din0 => VN1417_in0,
        Din1 => VN1417_in1,
        Din2 => VN1417_in2,
        Din3 => VN1417_in3,
        Din4 => VN1417_in4,
        Din5 => VN1417_in5,
        VN2CN0_bit => VN_data_out(8502),
        VN2CN1_bit => VN_data_out(8503),
        VN2CN2_bit => VN_data_out(8504),
        VN2CN3_bit => VN_data_out(8505),
        VN2CN4_bit => VN_data_out(8506),
        VN2CN5_bit => VN_data_out(8507),
        VN2CN0_sign => VN_sign_out(8502),
        VN2CN1_sign => VN_sign_out(8503),
        VN2CN2_sign => VN_sign_out(8504),
        VN2CN3_sign => VN_sign_out(8505),
        VN2CN4_sign => VN_sign_out(8506),
        VN2CN5_sign => VN_sign_out(8507),
        codeword => codeword(1417),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1418 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8513 downto 8508),
        Din0 => VN1418_in0,
        Din1 => VN1418_in1,
        Din2 => VN1418_in2,
        Din3 => VN1418_in3,
        Din4 => VN1418_in4,
        Din5 => VN1418_in5,
        VN2CN0_bit => VN_data_out(8508),
        VN2CN1_bit => VN_data_out(8509),
        VN2CN2_bit => VN_data_out(8510),
        VN2CN3_bit => VN_data_out(8511),
        VN2CN4_bit => VN_data_out(8512),
        VN2CN5_bit => VN_data_out(8513),
        VN2CN0_sign => VN_sign_out(8508),
        VN2CN1_sign => VN_sign_out(8509),
        VN2CN2_sign => VN_sign_out(8510),
        VN2CN3_sign => VN_sign_out(8511),
        VN2CN4_sign => VN_sign_out(8512),
        VN2CN5_sign => VN_sign_out(8513),
        codeword => codeword(1418),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1419 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8519 downto 8514),
        Din0 => VN1419_in0,
        Din1 => VN1419_in1,
        Din2 => VN1419_in2,
        Din3 => VN1419_in3,
        Din4 => VN1419_in4,
        Din5 => VN1419_in5,
        VN2CN0_bit => VN_data_out(8514),
        VN2CN1_bit => VN_data_out(8515),
        VN2CN2_bit => VN_data_out(8516),
        VN2CN3_bit => VN_data_out(8517),
        VN2CN4_bit => VN_data_out(8518),
        VN2CN5_bit => VN_data_out(8519),
        VN2CN0_sign => VN_sign_out(8514),
        VN2CN1_sign => VN_sign_out(8515),
        VN2CN2_sign => VN_sign_out(8516),
        VN2CN3_sign => VN_sign_out(8517),
        VN2CN4_sign => VN_sign_out(8518),
        VN2CN5_sign => VN_sign_out(8519),
        codeword => codeword(1419),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1420 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8525 downto 8520),
        Din0 => VN1420_in0,
        Din1 => VN1420_in1,
        Din2 => VN1420_in2,
        Din3 => VN1420_in3,
        Din4 => VN1420_in4,
        Din5 => VN1420_in5,
        VN2CN0_bit => VN_data_out(8520),
        VN2CN1_bit => VN_data_out(8521),
        VN2CN2_bit => VN_data_out(8522),
        VN2CN3_bit => VN_data_out(8523),
        VN2CN4_bit => VN_data_out(8524),
        VN2CN5_bit => VN_data_out(8525),
        VN2CN0_sign => VN_sign_out(8520),
        VN2CN1_sign => VN_sign_out(8521),
        VN2CN2_sign => VN_sign_out(8522),
        VN2CN3_sign => VN_sign_out(8523),
        VN2CN4_sign => VN_sign_out(8524),
        VN2CN5_sign => VN_sign_out(8525),
        codeword => codeword(1420),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1421 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8531 downto 8526),
        Din0 => VN1421_in0,
        Din1 => VN1421_in1,
        Din2 => VN1421_in2,
        Din3 => VN1421_in3,
        Din4 => VN1421_in4,
        Din5 => VN1421_in5,
        VN2CN0_bit => VN_data_out(8526),
        VN2CN1_bit => VN_data_out(8527),
        VN2CN2_bit => VN_data_out(8528),
        VN2CN3_bit => VN_data_out(8529),
        VN2CN4_bit => VN_data_out(8530),
        VN2CN5_bit => VN_data_out(8531),
        VN2CN0_sign => VN_sign_out(8526),
        VN2CN1_sign => VN_sign_out(8527),
        VN2CN2_sign => VN_sign_out(8528),
        VN2CN3_sign => VN_sign_out(8529),
        VN2CN4_sign => VN_sign_out(8530),
        VN2CN5_sign => VN_sign_out(8531),
        codeword => codeword(1421),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1422 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8537 downto 8532),
        Din0 => VN1422_in0,
        Din1 => VN1422_in1,
        Din2 => VN1422_in2,
        Din3 => VN1422_in3,
        Din4 => VN1422_in4,
        Din5 => VN1422_in5,
        VN2CN0_bit => VN_data_out(8532),
        VN2CN1_bit => VN_data_out(8533),
        VN2CN2_bit => VN_data_out(8534),
        VN2CN3_bit => VN_data_out(8535),
        VN2CN4_bit => VN_data_out(8536),
        VN2CN5_bit => VN_data_out(8537),
        VN2CN0_sign => VN_sign_out(8532),
        VN2CN1_sign => VN_sign_out(8533),
        VN2CN2_sign => VN_sign_out(8534),
        VN2CN3_sign => VN_sign_out(8535),
        VN2CN4_sign => VN_sign_out(8536),
        VN2CN5_sign => VN_sign_out(8537),
        codeword => codeword(1422),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1423 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8543 downto 8538),
        Din0 => VN1423_in0,
        Din1 => VN1423_in1,
        Din2 => VN1423_in2,
        Din3 => VN1423_in3,
        Din4 => VN1423_in4,
        Din5 => VN1423_in5,
        VN2CN0_bit => VN_data_out(8538),
        VN2CN1_bit => VN_data_out(8539),
        VN2CN2_bit => VN_data_out(8540),
        VN2CN3_bit => VN_data_out(8541),
        VN2CN4_bit => VN_data_out(8542),
        VN2CN5_bit => VN_data_out(8543),
        VN2CN0_sign => VN_sign_out(8538),
        VN2CN1_sign => VN_sign_out(8539),
        VN2CN2_sign => VN_sign_out(8540),
        VN2CN3_sign => VN_sign_out(8541),
        VN2CN4_sign => VN_sign_out(8542),
        VN2CN5_sign => VN_sign_out(8543),
        codeword => codeword(1423),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1424 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8549 downto 8544),
        Din0 => VN1424_in0,
        Din1 => VN1424_in1,
        Din2 => VN1424_in2,
        Din3 => VN1424_in3,
        Din4 => VN1424_in4,
        Din5 => VN1424_in5,
        VN2CN0_bit => VN_data_out(8544),
        VN2CN1_bit => VN_data_out(8545),
        VN2CN2_bit => VN_data_out(8546),
        VN2CN3_bit => VN_data_out(8547),
        VN2CN4_bit => VN_data_out(8548),
        VN2CN5_bit => VN_data_out(8549),
        VN2CN0_sign => VN_sign_out(8544),
        VN2CN1_sign => VN_sign_out(8545),
        VN2CN2_sign => VN_sign_out(8546),
        VN2CN3_sign => VN_sign_out(8547),
        VN2CN4_sign => VN_sign_out(8548),
        VN2CN5_sign => VN_sign_out(8549),
        codeword => codeword(1424),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1425 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8555 downto 8550),
        Din0 => VN1425_in0,
        Din1 => VN1425_in1,
        Din2 => VN1425_in2,
        Din3 => VN1425_in3,
        Din4 => VN1425_in4,
        Din5 => VN1425_in5,
        VN2CN0_bit => VN_data_out(8550),
        VN2CN1_bit => VN_data_out(8551),
        VN2CN2_bit => VN_data_out(8552),
        VN2CN3_bit => VN_data_out(8553),
        VN2CN4_bit => VN_data_out(8554),
        VN2CN5_bit => VN_data_out(8555),
        VN2CN0_sign => VN_sign_out(8550),
        VN2CN1_sign => VN_sign_out(8551),
        VN2CN2_sign => VN_sign_out(8552),
        VN2CN3_sign => VN_sign_out(8553),
        VN2CN4_sign => VN_sign_out(8554),
        VN2CN5_sign => VN_sign_out(8555),
        codeword => codeword(1425),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1426 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8561 downto 8556),
        Din0 => VN1426_in0,
        Din1 => VN1426_in1,
        Din2 => VN1426_in2,
        Din3 => VN1426_in3,
        Din4 => VN1426_in4,
        Din5 => VN1426_in5,
        VN2CN0_bit => VN_data_out(8556),
        VN2CN1_bit => VN_data_out(8557),
        VN2CN2_bit => VN_data_out(8558),
        VN2CN3_bit => VN_data_out(8559),
        VN2CN4_bit => VN_data_out(8560),
        VN2CN5_bit => VN_data_out(8561),
        VN2CN0_sign => VN_sign_out(8556),
        VN2CN1_sign => VN_sign_out(8557),
        VN2CN2_sign => VN_sign_out(8558),
        VN2CN3_sign => VN_sign_out(8559),
        VN2CN4_sign => VN_sign_out(8560),
        VN2CN5_sign => VN_sign_out(8561),
        codeword => codeword(1426),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1427 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8567 downto 8562),
        Din0 => VN1427_in0,
        Din1 => VN1427_in1,
        Din2 => VN1427_in2,
        Din3 => VN1427_in3,
        Din4 => VN1427_in4,
        Din5 => VN1427_in5,
        VN2CN0_bit => VN_data_out(8562),
        VN2CN1_bit => VN_data_out(8563),
        VN2CN2_bit => VN_data_out(8564),
        VN2CN3_bit => VN_data_out(8565),
        VN2CN4_bit => VN_data_out(8566),
        VN2CN5_bit => VN_data_out(8567),
        VN2CN0_sign => VN_sign_out(8562),
        VN2CN1_sign => VN_sign_out(8563),
        VN2CN2_sign => VN_sign_out(8564),
        VN2CN3_sign => VN_sign_out(8565),
        VN2CN4_sign => VN_sign_out(8566),
        VN2CN5_sign => VN_sign_out(8567),
        codeword => codeword(1427),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1428 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8573 downto 8568),
        Din0 => VN1428_in0,
        Din1 => VN1428_in1,
        Din2 => VN1428_in2,
        Din3 => VN1428_in3,
        Din4 => VN1428_in4,
        Din5 => VN1428_in5,
        VN2CN0_bit => VN_data_out(8568),
        VN2CN1_bit => VN_data_out(8569),
        VN2CN2_bit => VN_data_out(8570),
        VN2CN3_bit => VN_data_out(8571),
        VN2CN4_bit => VN_data_out(8572),
        VN2CN5_bit => VN_data_out(8573),
        VN2CN0_sign => VN_sign_out(8568),
        VN2CN1_sign => VN_sign_out(8569),
        VN2CN2_sign => VN_sign_out(8570),
        VN2CN3_sign => VN_sign_out(8571),
        VN2CN4_sign => VN_sign_out(8572),
        VN2CN5_sign => VN_sign_out(8573),
        codeword => codeword(1428),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1429 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8579 downto 8574),
        Din0 => VN1429_in0,
        Din1 => VN1429_in1,
        Din2 => VN1429_in2,
        Din3 => VN1429_in3,
        Din4 => VN1429_in4,
        Din5 => VN1429_in5,
        VN2CN0_bit => VN_data_out(8574),
        VN2CN1_bit => VN_data_out(8575),
        VN2CN2_bit => VN_data_out(8576),
        VN2CN3_bit => VN_data_out(8577),
        VN2CN4_bit => VN_data_out(8578),
        VN2CN5_bit => VN_data_out(8579),
        VN2CN0_sign => VN_sign_out(8574),
        VN2CN1_sign => VN_sign_out(8575),
        VN2CN2_sign => VN_sign_out(8576),
        VN2CN3_sign => VN_sign_out(8577),
        VN2CN4_sign => VN_sign_out(8578),
        VN2CN5_sign => VN_sign_out(8579),
        codeword => codeword(1429),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1430 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8585 downto 8580),
        Din0 => VN1430_in0,
        Din1 => VN1430_in1,
        Din2 => VN1430_in2,
        Din3 => VN1430_in3,
        Din4 => VN1430_in4,
        Din5 => VN1430_in5,
        VN2CN0_bit => VN_data_out(8580),
        VN2CN1_bit => VN_data_out(8581),
        VN2CN2_bit => VN_data_out(8582),
        VN2CN3_bit => VN_data_out(8583),
        VN2CN4_bit => VN_data_out(8584),
        VN2CN5_bit => VN_data_out(8585),
        VN2CN0_sign => VN_sign_out(8580),
        VN2CN1_sign => VN_sign_out(8581),
        VN2CN2_sign => VN_sign_out(8582),
        VN2CN3_sign => VN_sign_out(8583),
        VN2CN4_sign => VN_sign_out(8584),
        VN2CN5_sign => VN_sign_out(8585),
        codeword => codeword(1430),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1431 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8591 downto 8586),
        Din0 => VN1431_in0,
        Din1 => VN1431_in1,
        Din2 => VN1431_in2,
        Din3 => VN1431_in3,
        Din4 => VN1431_in4,
        Din5 => VN1431_in5,
        VN2CN0_bit => VN_data_out(8586),
        VN2CN1_bit => VN_data_out(8587),
        VN2CN2_bit => VN_data_out(8588),
        VN2CN3_bit => VN_data_out(8589),
        VN2CN4_bit => VN_data_out(8590),
        VN2CN5_bit => VN_data_out(8591),
        VN2CN0_sign => VN_sign_out(8586),
        VN2CN1_sign => VN_sign_out(8587),
        VN2CN2_sign => VN_sign_out(8588),
        VN2CN3_sign => VN_sign_out(8589),
        VN2CN4_sign => VN_sign_out(8590),
        VN2CN5_sign => VN_sign_out(8591),
        codeword => codeword(1431),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1432 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8597 downto 8592),
        Din0 => VN1432_in0,
        Din1 => VN1432_in1,
        Din2 => VN1432_in2,
        Din3 => VN1432_in3,
        Din4 => VN1432_in4,
        Din5 => VN1432_in5,
        VN2CN0_bit => VN_data_out(8592),
        VN2CN1_bit => VN_data_out(8593),
        VN2CN2_bit => VN_data_out(8594),
        VN2CN3_bit => VN_data_out(8595),
        VN2CN4_bit => VN_data_out(8596),
        VN2CN5_bit => VN_data_out(8597),
        VN2CN0_sign => VN_sign_out(8592),
        VN2CN1_sign => VN_sign_out(8593),
        VN2CN2_sign => VN_sign_out(8594),
        VN2CN3_sign => VN_sign_out(8595),
        VN2CN4_sign => VN_sign_out(8596),
        VN2CN5_sign => VN_sign_out(8597),
        codeword => codeword(1432),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1433 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8603 downto 8598),
        Din0 => VN1433_in0,
        Din1 => VN1433_in1,
        Din2 => VN1433_in2,
        Din3 => VN1433_in3,
        Din4 => VN1433_in4,
        Din5 => VN1433_in5,
        VN2CN0_bit => VN_data_out(8598),
        VN2CN1_bit => VN_data_out(8599),
        VN2CN2_bit => VN_data_out(8600),
        VN2CN3_bit => VN_data_out(8601),
        VN2CN4_bit => VN_data_out(8602),
        VN2CN5_bit => VN_data_out(8603),
        VN2CN0_sign => VN_sign_out(8598),
        VN2CN1_sign => VN_sign_out(8599),
        VN2CN2_sign => VN_sign_out(8600),
        VN2CN3_sign => VN_sign_out(8601),
        VN2CN4_sign => VN_sign_out(8602),
        VN2CN5_sign => VN_sign_out(8603),
        codeword => codeword(1433),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1434 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8609 downto 8604),
        Din0 => VN1434_in0,
        Din1 => VN1434_in1,
        Din2 => VN1434_in2,
        Din3 => VN1434_in3,
        Din4 => VN1434_in4,
        Din5 => VN1434_in5,
        VN2CN0_bit => VN_data_out(8604),
        VN2CN1_bit => VN_data_out(8605),
        VN2CN2_bit => VN_data_out(8606),
        VN2CN3_bit => VN_data_out(8607),
        VN2CN4_bit => VN_data_out(8608),
        VN2CN5_bit => VN_data_out(8609),
        VN2CN0_sign => VN_sign_out(8604),
        VN2CN1_sign => VN_sign_out(8605),
        VN2CN2_sign => VN_sign_out(8606),
        VN2CN3_sign => VN_sign_out(8607),
        VN2CN4_sign => VN_sign_out(8608),
        VN2CN5_sign => VN_sign_out(8609),
        codeword => codeword(1434),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1435 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8615 downto 8610),
        Din0 => VN1435_in0,
        Din1 => VN1435_in1,
        Din2 => VN1435_in2,
        Din3 => VN1435_in3,
        Din4 => VN1435_in4,
        Din5 => VN1435_in5,
        VN2CN0_bit => VN_data_out(8610),
        VN2CN1_bit => VN_data_out(8611),
        VN2CN2_bit => VN_data_out(8612),
        VN2CN3_bit => VN_data_out(8613),
        VN2CN4_bit => VN_data_out(8614),
        VN2CN5_bit => VN_data_out(8615),
        VN2CN0_sign => VN_sign_out(8610),
        VN2CN1_sign => VN_sign_out(8611),
        VN2CN2_sign => VN_sign_out(8612),
        VN2CN3_sign => VN_sign_out(8613),
        VN2CN4_sign => VN_sign_out(8614),
        VN2CN5_sign => VN_sign_out(8615),
        codeword => codeword(1435),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1436 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8621 downto 8616),
        Din0 => VN1436_in0,
        Din1 => VN1436_in1,
        Din2 => VN1436_in2,
        Din3 => VN1436_in3,
        Din4 => VN1436_in4,
        Din5 => VN1436_in5,
        VN2CN0_bit => VN_data_out(8616),
        VN2CN1_bit => VN_data_out(8617),
        VN2CN2_bit => VN_data_out(8618),
        VN2CN3_bit => VN_data_out(8619),
        VN2CN4_bit => VN_data_out(8620),
        VN2CN5_bit => VN_data_out(8621),
        VN2CN0_sign => VN_sign_out(8616),
        VN2CN1_sign => VN_sign_out(8617),
        VN2CN2_sign => VN_sign_out(8618),
        VN2CN3_sign => VN_sign_out(8619),
        VN2CN4_sign => VN_sign_out(8620),
        VN2CN5_sign => VN_sign_out(8621),
        codeword => codeword(1436),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1437 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8627 downto 8622),
        Din0 => VN1437_in0,
        Din1 => VN1437_in1,
        Din2 => VN1437_in2,
        Din3 => VN1437_in3,
        Din4 => VN1437_in4,
        Din5 => VN1437_in5,
        VN2CN0_bit => VN_data_out(8622),
        VN2CN1_bit => VN_data_out(8623),
        VN2CN2_bit => VN_data_out(8624),
        VN2CN3_bit => VN_data_out(8625),
        VN2CN4_bit => VN_data_out(8626),
        VN2CN5_bit => VN_data_out(8627),
        VN2CN0_sign => VN_sign_out(8622),
        VN2CN1_sign => VN_sign_out(8623),
        VN2CN2_sign => VN_sign_out(8624),
        VN2CN3_sign => VN_sign_out(8625),
        VN2CN4_sign => VN_sign_out(8626),
        VN2CN5_sign => VN_sign_out(8627),
        codeword => codeword(1437),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1438 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8633 downto 8628),
        Din0 => VN1438_in0,
        Din1 => VN1438_in1,
        Din2 => VN1438_in2,
        Din3 => VN1438_in3,
        Din4 => VN1438_in4,
        Din5 => VN1438_in5,
        VN2CN0_bit => VN_data_out(8628),
        VN2CN1_bit => VN_data_out(8629),
        VN2CN2_bit => VN_data_out(8630),
        VN2CN3_bit => VN_data_out(8631),
        VN2CN4_bit => VN_data_out(8632),
        VN2CN5_bit => VN_data_out(8633),
        VN2CN0_sign => VN_sign_out(8628),
        VN2CN1_sign => VN_sign_out(8629),
        VN2CN2_sign => VN_sign_out(8630),
        VN2CN3_sign => VN_sign_out(8631),
        VN2CN4_sign => VN_sign_out(8632),
        VN2CN5_sign => VN_sign_out(8633),
        codeword => codeword(1438),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1439 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8639 downto 8634),
        Din0 => VN1439_in0,
        Din1 => VN1439_in1,
        Din2 => VN1439_in2,
        Din3 => VN1439_in3,
        Din4 => VN1439_in4,
        Din5 => VN1439_in5,
        VN2CN0_bit => VN_data_out(8634),
        VN2CN1_bit => VN_data_out(8635),
        VN2CN2_bit => VN_data_out(8636),
        VN2CN3_bit => VN_data_out(8637),
        VN2CN4_bit => VN_data_out(8638),
        VN2CN5_bit => VN_data_out(8639),
        VN2CN0_sign => VN_sign_out(8634),
        VN2CN1_sign => VN_sign_out(8635),
        VN2CN2_sign => VN_sign_out(8636),
        VN2CN3_sign => VN_sign_out(8637),
        VN2CN4_sign => VN_sign_out(8638),
        VN2CN5_sign => VN_sign_out(8639),
        codeword => codeword(1439),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1440 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8645 downto 8640),
        Din0 => VN1440_in0,
        Din1 => VN1440_in1,
        Din2 => VN1440_in2,
        Din3 => VN1440_in3,
        Din4 => VN1440_in4,
        Din5 => VN1440_in5,
        VN2CN0_bit => VN_data_out(8640),
        VN2CN1_bit => VN_data_out(8641),
        VN2CN2_bit => VN_data_out(8642),
        VN2CN3_bit => VN_data_out(8643),
        VN2CN4_bit => VN_data_out(8644),
        VN2CN5_bit => VN_data_out(8645),
        VN2CN0_sign => VN_sign_out(8640),
        VN2CN1_sign => VN_sign_out(8641),
        VN2CN2_sign => VN_sign_out(8642),
        VN2CN3_sign => VN_sign_out(8643),
        VN2CN4_sign => VN_sign_out(8644),
        VN2CN5_sign => VN_sign_out(8645),
        codeword => codeword(1440),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1441 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8651 downto 8646),
        Din0 => VN1441_in0,
        Din1 => VN1441_in1,
        Din2 => VN1441_in2,
        Din3 => VN1441_in3,
        Din4 => VN1441_in4,
        Din5 => VN1441_in5,
        VN2CN0_bit => VN_data_out(8646),
        VN2CN1_bit => VN_data_out(8647),
        VN2CN2_bit => VN_data_out(8648),
        VN2CN3_bit => VN_data_out(8649),
        VN2CN4_bit => VN_data_out(8650),
        VN2CN5_bit => VN_data_out(8651),
        VN2CN0_sign => VN_sign_out(8646),
        VN2CN1_sign => VN_sign_out(8647),
        VN2CN2_sign => VN_sign_out(8648),
        VN2CN3_sign => VN_sign_out(8649),
        VN2CN4_sign => VN_sign_out(8650),
        VN2CN5_sign => VN_sign_out(8651),
        codeword => codeword(1441),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1442 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8657 downto 8652),
        Din0 => VN1442_in0,
        Din1 => VN1442_in1,
        Din2 => VN1442_in2,
        Din3 => VN1442_in3,
        Din4 => VN1442_in4,
        Din5 => VN1442_in5,
        VN2CN0_bit => VN_data_out(8652),
        VN2CN1_bit => VN_data_out(8653),
        VN2CN2_bit => VN_data_out(8654),
        VN2CN3_bit => VN_data_out(8655),
        VN2CN4_bit => VN_data_out(8656),
        VN2CN5_bit => VN_data_out(8657),
        VN2CN0_sign => VN_sign_out(8652),
        VN2CN1_sign => VN_sign_out(8653),
        VN2CN2_sign => VN_sign_out(8654),
        VN2CN3_sign => VN_sign_out(8655),
        VN2CN4_sign => VN_sign_out(8656),
        VN2CN5_sign => VN_sign_out(8657),
        codeword => codeword(1442),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1443 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8663 downto 8658),
        Din0 => VN1443_in0,
        Din1 => VN1443_in1,
        Din2 => VN1443_in2,
        Din3 => VN1443_in3,
        Din4 => VN1443_in4,
        Din5 => VN1443_in5,
        VN2CN0_bit => VN_data_out(8658),
        VN2CN1_bit => VN_data_out(8659),
        VN2CN2_bit => VN_data_out(8660),
        VN2CN3_bit => VN_data_out(8661),
        VN2CN4_bit => VN_data_out(8662),
        VN2CN5_bit => VN_data_out(8663),
        VN2CN0_sign => VN_sign_out(8658),
        VN2CN1_sign => VN_sign_out(8659),
        VN2CN2_sign => VN_sign_out(8660),
        VN2CN3_sign => VN_sign_out(8661),
        VN2CN4_sign => VN_sign_out(8662),
        VN2CN5_sign => VN_sign_out(8663),
        codeword => codeword(1443),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1444 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8669 downto 8664),
        Din0 => VN1444_in0,
        Din1 => VN1444_in1,
        Din2 => VN1444_in2,
        Din3 => VN1444_in3,
        Din4 => VN1444_in4,
        Din5 => VN1444_in5,
        VN2CN0_bit => VN_data_out(8664),
        VN2CN1_bit => VN_data_out(8665),
        VN2CN2_bit => VN_data_out(8666),
        VN2CN3_bit => VN_data_out(8667),
        VN2CN4_bit => VN_data_out(8668),
        VN2CN5_bit => VN_data_out(8669),
        VN2CN0_sign => VN_sign_out(8664),
        VN2CN1_sign => VN_sign_out(8665),
        VN2CN2_sign => VN_sign_out(8666),
        VN2CN3_sign => VN_sign_out(8667),
        VN2CN4_sign => VN_sign_out(8668),
        VN2CN5_sign => VN_sign_out(8669),
        codeword => codeword(1444),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1445 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8675 downto 8670),
        Din0 => VN1445_in0,
        Din1 => VN1445_in1,
        Din2 => VN1445_in2,
        Din3 => VN1445_in3,
        Din4 => VN1445_in4,
        Din5 => VN1445_in5,
        VN2CN0_bit => VN_data_out(8670),
        VN2CN1_bit => VN_data_out(8671),
        VN2CN2_bit => VN_data_out(8672),
        VN2CN3_bit => VN_data_out(8673),
        VN2CN4_bit => VN_data_out(8674),
        VN2CN5_bit => VN_data_out(8675),
        VN2CN0_sign => VN_sign_out(8670),
        VN2CN1_sign => VN_sign_out(8671),
        VN2CN2_sign => VN_sign_out(8672),
        VN2CN3_sign => VN_sign_out(8673),
        VN2CN4_sign => VN_sign_out(8674),
        VN2CN5_sign => VN_sign_out(8675),
        codeword => codeword(1445),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1446 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8681 downto 8676),
        Din0 => VN1446_in0,
        Din1 => VN1446_in1,
        Din2 => VN1446_in2,
        Din3 => VN1446_in3,
        Din4 => VN1446_in4,
        Din5 => VN1446_in5,
        VN2CN0_bit => VN_data_out(8676),
        VN2CN1_bit => VN_data_out(8677),
        VN2CN2_bit => VN_data_out(8678),
        VN2CN3_bit => VN_data_out(8679),
        VN2CN4_bit => VN_data_out(8680),
        VN2CN5_bit => VN_data_out(8681),
        VN2CN0_sign => VN_sign_out(8676),
        VN2CN1_sign => VN_sign_out(8677),
        VN2CN2_sign => VN_sign_out(8678),
        VN2CN3_sign => VN_sign_out(8679),
        VN2CN4_sign => VN_sign_out(8680),
        VN2CN5_sign => VN_sign_out(8681),
        codeword => codeword(1446),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1447 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8687 downto 8682),
        Din0 => VN1447_in0,
        Din1 => VN1447_in1,
        Din2 => VN1447_in2,
        Din3 => VN1447_in3,
        Din4 => VN1447_in4,
        Din5 => VN1447_in5,
        VN2CN0_bit => VN_data_out(8682),
        VN2CN1_bit => VN_data_out(8683),
        VN2CN2_bit => VN_data_out(8684),
        VN2CN3_bit => VN_data_out(8685),
        VN2CN4_bit => VN_data_out(8686),
        VN2CN5_bit => VN_data_out(8687),
        VN2CN0_sign => VN_sign_out(8682),
        VN2CN1_sign => VN_sign_out(8683),
        VN2CN2_sign => VN_sign_out(8684),
        VN2CN3_sign => VN_sign_out(8685),
        VN2CN4_sign => VN_sign_out(8686),
        VN2CN5_sign => VN_sign_out(8687),
        codeword => codeword(1447),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1448 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8693 downto 8688),
        Din0 => VN1448_in0,
        Din1 => VN1448_in1,
        Din2 => VN1448_in2,
        Din3 => VN1448_in3,
        Din4 => VN1448_in4,
        Din5 => VN1448_in5,
        VN2CN0_bit => VN_data_out(8688),
        VN2CN1_bit => VN_data_out(8689),
        VN2CN2_bit => VN_data_out(8690),
        VN2CN3_bit => VN_data_out(8691),
        VN2CN4_bit => VN_data_out(8692),
        VN2CN5_bit => VN_data_out(8693),
        VN2CN0_sign => VN_sign_out(8688),
        VN2CN1_sign => VN_sign_out(8689),
        VN2CN2_sign => VN_sign_out(8690),
        VN2CN3_sign => VN_sign_out(8691),
        VN2CN4_sign => VN_sign_out(8692),
        VN2CN5_sign => VN_sign_out(8693),
        codeword => codeword(1448),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1449 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8699 downto 8694),
        Din0 => VN1449_in0,
        Din1 => VN1449_in1,
        Din2 => VN1449_in2,
        Din3 => VN1449_in3,
        Din4 => VN1449_in4,
        Din5 => VN1449_in5,
        VN2CN0_bit => VN_data_out(8694),
        VN2CN1_bit => VN_data_out(8695),
        VN2CN2_bit => VN_data_out(8696),
        VN2CN3_bit => VN_data_out(8697),
        VN2CN4_bit => VN_data_out(8698),
        VN2CN5_bit => VN_data_out(8699),
        VN2CN0_sign => VN_sign_out(8694),
        VN2CN1_sign => VN_sign_out(8695),
        VN2CN2_sign => VN_sign_out(8696),
        VN2CN3_sign => VN_sign_out(8697),
        VN2CN4_sign => VN_sign_out(8698),
        VN2CN5_sign => VN_sign_out(8699),
        codeword => codeword(1449),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1450 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8705 downto 8700),
        Din0 => VN1450_in0,
        Din1 => VN1450_in1,
        Din2 => VN1450_in2,
        Din3 => VN1450_in3,
        Din4 => VN1450_in4,
        Din5 => VN1450_in5,
        VN2CN0_bit => VN_data_out(8700),
        VN2CN1_bit => VN_data_out(8701),
        VN2CN2_bit => VN_data_out(8702),
        VN2CN3_bit => VN_data_out(8703),
        VN2CN4_bit => VN_data_out(8704),
        VN2CN5_bit => VN_data_out(8705),
        VN2CN0_sign => VN_sign_out(8700),
        VN2CN1_sign => VN_sign_out(8701),
        VN2CN2_sign => VN_sign_out(8702),
        VN2CN3_sign => VN_sign_out(8703),
        VN2CN4_sign => VN_sign_out(8704),
        VN2CN5_sign => VN_sign_out(8705),
        codeword => codeword(1450),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1451 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8711 downto 8706),
        Din0 => VN1451_in0,
        Din1 => VN1451_in1,
        Din2 => VN1451_in2,
        Din3 => VN1451_in3,
        Din4 => VN1451_in4,
        Din5 => VN1451_in5,
        VN2CN0_bit => VN_data_out(8706),
        VN2CN1_bit => VN_data_out(8707),
        VN2CN2_bit => VN_data_out(8708),
        VN2CN3_bit => VN_data_out(8709),
        VN2CN4_bit => VN_data_out(8710),
        VN2CN5_bit => VN_data_out(8711),
        VN2CN0_sign => VN_sign_out(8706),
        VN2CN1_sign => VN_sign_out(8707),
        VN2CN2_sign => VN_sign_out(8708),
        VN2CN3_sign => VN_sign_out(8709),
        VN2CN4_sign => VN_sign_out(8710),
        VN2CN5_sign => VN_sign_out(8711),
        codeword => codeword(1451),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1452 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8717 downto 8712),
        Din0 => VN1452_in0,
        Din1 => VN1452_in1,
        Din2 => VN1452_in2,
        Din3 => VN1452_in3,
        Din4 => VN1452_in4,
        Din5 => VN1452_in5,
        VN2CN0_bit => VN_data_out(8712),
        VN2CN1_bit => VN_data_out(8713),
        VN2CN2_bit => VN_data_out(8714),
        VN2CN3_bit => VN_data_out(8715),
        VN2CN4_bit => VN_data_out(8716),
        VN2CN5_bit => VN_data_out(8717),
        VN2CN0_sign => VN_sign_out(8712),
        VN2CN1_sign => VN_sign_out(8713),
        VN2CN2_sign => VN_sign_out(8714),
        VN2CN3_sign => VN_sign_out(8715),
        VN2CN4_sign => VN_sign_out(8716),
        VN2CN5_sign => VN_sign_out(8717),
        codeword => codeword(1452),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1453 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8723 downto 8718),
        Din0 => VN1453_in0,
        Din1 => VN1453_in1,
        Din2 => VN1453_in2,
        Din3 => VN1453_in3,
        Din4 => VN1453_in4,
        Din5 => VN1453_in5,
        VN2CN0_bit => VN_data_out(8718),
        VN2CN1_bit => VN_data_out(8719),
        VN2CN2_bit => VN_data_out(8720),
        VN2CN3_bit => VN_data_out(8721),
        VN2CN4_bit => VN_data_out(8722),
        VN2CN5_bit => VN_data_out(8723),
        VN2CN0_sign => VN_sign_out(8718),
        VN2CN1_sign => VN_sign_out(8719),
        VN2CN2_sign => VN_sign_out(8720),
        VN2CN3_sign => VN_sign_out(8721),
        VN2CN4_sign => VN_sign_out(8722),
        VN2CN5_sign => VN_sign_out(8723),
        codeword => codeword(1453),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1454 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8729 downto 8724),
        Din0 => VN1454_in0,
        Din1 => VN1454_in1,
        Din2 => VN1454_in2,
        Din3 => VN1454_in3,
        Din4 => VN1454_in4,
        Din5 => VN1454_in5,
        VN2CN0_bit => VN_data_out(8724),
        VN2CN1_bit => VN_data_out(8725),
        VN2CN2_bit => VN_data_out(8726),
        VN2CN3_bit => VN_data_out(8727),
        VN2CN4_bit => VN_data_out(8728),
        VN2CN5_bit => VN_data_out(8729),
        VN2CN0_sign => VN_sign_out(8724),
        VN2CN1_sign => VN_sign_out(8725),
        VN2CN2_sign => VN_sign_out(8726),
        VN2CN3_sign => VN_sign_out(8727),
        VN2CN4_sign => VN_sign_out(8728),
        VN2CN5_sign => VN_sign_out(8729),
        codeword => codeword(1454),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1455 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8735 downto 8730),
        Din0 => VN1455_in0,
        Din1 => VN1455_in1,
        Din2 => VN1455_in2,
        Din3 => VN1455_in3,
        Din4 => VN1455_in4,
        Din5 => VN1455_in5,
        VN2CN0_bit => VN_data_out(8730),
        VN2CN1_bit => VN_data_out(8731),
        VN2CN2_bit => VN_data_out(8732),
        VN2CN3_bit => VN_data_out(8733),
        VN2CN4_bit => VN_data_out(8734),
        VN2CN5_bit => VN_data_out(8735),
        VN2CN0_sign => VN_sign_out(8730),
        VN2CN1_sign => VN_sign_out(8731),
        VN2CN2_sign => VN_sign_out(8732),
        VN2CN3_sign => VN_sign_out(8733),
        VN2CN4_sign => VN_sign_out(8734),
        VN2CN5_sign => VN_sign_out(8735),
        codeword => codeword(1455),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1456 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8741 downto 8736),
        Din0 => VN1456_in0,
        Din1 => VN1456_in1,
        Din2 => VN1456_in2,
        Din3 => VN1456_in3,
        Din4 => VN1456_in4,
        Din5 => VN1456_in5,
        VN2CN0_bit => VN_data_out(8736),
        VN2CN1_bit => VN_data_out(8737),
        VN2CN2_bit => VN_data_out(8738),
        VN2CN3_bit => VN_data_out(8739),
        VN2CN4_bit => VN_data_out(8740),
        VN2CN5_bit => VN_data_out(8741),
        VN2CN0_sign => VN_sign_out(8736),
        VN2CN1_sign => VN_sign_out(8737),
        VN2CN2_sign => VN_sign_out(8738),
        VN2CN3_sign => VN_sign_out(8739),
        VN2CN4_sign => VN_sign_out(8740),
        VN2CN5_sign => VN_sign_out(8741),
        codeword => codeword(1456),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1457 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8747 downto 8742),
        Din0 => VN1457_in0,
        Din1 => VN1457_in1,
        Din2 => VN1457_in2,
        Din3 => VN1457_in3,
        Din4 => VN1457_in4,
        Din5 => VN1457_in5,
        VN2CN0_bit => VN_data_out(8742),
        VN2CN1_bit => VN_data_out(8743),
        VN2CN2_bit => VN_data_out(8744),
        VN2CN3_bit => VN_data_out(8745),
        VN2CN4_bit => VN_data_out(8746),
        VN2CN5_bit => VN_data_out(8747),
        VN2CN0_sign => VN_sign_out(8742),
        VN2CN1_sign => VN_sign_out(8743),
        VN2CN2_sign => VN_sign_out(8744),
        VN2CN3_sign => VN_sign_out(8745),
        VN2CN4_sign => VN_sign_out(8746),
        VN2CN5_sign => VN_sign_out(8747),
        codeword => codeword(1457),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1458 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8753 downto 8748),
        Din0 => VN1458_in0,
        Din1 => VN1458_in1,
        Din2 => VN1458_in2,
        Din3 => VN1458_in3,
        Din4 => VN1458_in4,
        Din5 => VN1458_in5,
        VN2CN0_bit => VN_data_out(8748),
        VN2CN1_bit => VN_data_out(8749),
        VN2CN2_bit => VN_data_out(8750),
        VN2CN3_bit => VN_data_out(8751),
        VN2CN4_bit => VN_data_out(8752),
        VN2CN5_bit => VN_data_out(8753),
        VN2CN0_sign => VN_sign_out(8748),
        VN2CN1_sign => VN_sign_out(8749),
        VN2CN2_sign => VN_sign_out(8750),
        VN2CN3_sign => VN_sign_out(8751),
        VN2CN4_sign => VN_sign_out(8752),
        VN2CN5_sign => VN_sign_out(8753),
        codeword => codeword(1458),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1459 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8759 downto 8754),
        Din0 => VN1459_in0,
        Din1 => VN1459_in1,
        Din2 => VN1459_in2,
        Din3 => VN1459_in3,
        Din4 => VN1459_in4,
        Din5 => VN1459_in5,
        VN2CN0_bit => VN_data_out(8754),
        VN2CN1_bit => VN_data_out(8755),
        VN2CN2_bit => VN_data_out(8756),
        VN2CN3_bit => VN_data_out(8757),
        VN2CN4_bit => VN_data_out(8758),
        VN2CN5_bit => VN_data_out(8759),
        VN2CN0_sign => VN_sign_out(8754),
        VN2CN1_sign => VN_sign_out(8755),
        VN2CN2_sign => VN_sign_out(8756),
        VN2CN3_sign => VN_sign_out(8757),
        VN2CN4_sign => VN_sign_out(8758),
        VN2CN5_sign => VN_sign_out(8759),
        codeword => codeword(1459),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1460 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8765 downto 8760),
        Din0 => VN1460_in0,
        Din1 => VN1460_in1,
        Din2 => VN1460_in2,
        Din3 => VN1460_in3,
        Din4 => VN1460_in4,
        Din5 => VN1460_in5,
        VN2CN0_bit => VN_data_out(8760),
        VN2CN1_bit => VN_data_out(8761),
        VN2CN2_bit => VN_data_out(8762),
        VN2CN3_bit => VN_data_out(8763),
        VN2CN4_bit => VN_data_out(8764),
        VN2CN5_bit => VN_data_out(8765),
        VN2CN0_sign => VN_sign_out(8760),
        VN2CN1_sign => VN_sign_out(8761),
        VN2CN2_sign => VN_sign_out(8762),
        VN2CN3_sign => VN_sign_out(8763),
        VN2CN4_sign => VN_sign_out(8764),
        VN2CN5_sign => VN_sign_out(8765),
        codeword => codeword(1460),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1461 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8771 downto 8766),
        Din0 => VN1461_in0,
        Din1 => VN1461_in1,
        Din2 => VN1461_in2,
        Din3 => VN1461_in3,
        Din4 => VN1461_in4,
        Din5 => VN1461_in5,
        VN2CN0_bit => VN_data_out(8766),
        VN2CN1_bit => VN_data_out(8767),
        VN2CN2_bit => VN_data_out(8768),
        VN2CN3_bit => VN_data_out(8769),
        VN2CN4_bit => VN_data_out(8770),
        VN2CN5_bit => VN_data_out(8771),
        VN2CN0_sign => VN_sign_out(8766),
        VN2CN1_sign => VN_sign_out(8767),
        VN2CN2_sign => VN_sign_out(8768),
        VN2CN3_sign => VN_sign_out(8769),
        VN2CN4_sign => VN_sign_out(8770),
        VN2CN5_sign => VN_sign_out(8771),
        codeword => codeword(1461),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1462 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8777 downto 8772),
        Din0 => VN1462_in0,
        Din1 => VN1462_in1,
        Din2 => VN1462_in2,
        Din3 => VN1462_in3,
        Din4 => VN1462_in4,
        Din5 => VN1462_in5,
        VN2CN0_bit => VN_data_out(8772),
        VN2CN1_bit => VN_data_out(8773),
        VN2CN2_bit => VN_data_out(8774),
        VN2CN3_bit => VN_data_out(8775),
        VN2CN4_bit => VN_data_out(8776),
        VN2CN5_bit => VN_data_out(8777),
        VN2CN0_sign => VN_sign_out(8772),
        VN2CN1_sign => VN_sign_out(8773),
        VN2CN2_sign => VN_sign_out(8774),
        VN2CN3_sign => VN_sign_out(8775),
        VN2CN4_sign => VN_sign_out(8776),
        VN2CN5_sign => VN_sign_out(8777),
        codeword => codeword(1462),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1463 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8783 downto 8778),
        Din0 => VN1463_in0,
        Din1 => VN1463_in1,
        Din2 => VN1463_in2,
        Din3 => VN1463_in3,
        Din4 => VN1463_in4,
        Din5 => VN1463_in5,
        VN2CN0_bit => VN_data_out(8778),
        VN2CN1_bit => VN_data_out(8779),
        VN2CN2_bit => VN_data_out(8780),
        VN2CN3_bit => VN_data_out(8781),
        VN2CN4_bit => VN_data_out(8782),
        VN2CN5_bit => VN_data_out(8783),
        VN2CN0_sign => VN_sign_out(8778),
        VN2CN1_sign => VN_sign_out(8779),
        VN2CN2_sign => VN_sign_out(8780),
        VN2CN3_sign => VN_sign_out(8781),
        VN2CN4_sign => VN_sign_out(8782),
        VN2CN5_sign => VN_sign_out(8783),
        codeword => codeword(1463),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1464 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8789 downto 8784),
        Din0 => VN1464_in0,
        Din1 => VN1464_in1,
        Din2 => VN1464_in2,
        Din3 => VN1464_in3,
        Din4 => VN1464_in4,
        Din5 => VN1464_in5,
        VN2CN0_bit => VN_data_out(8784),
        VN2CN1_bit => VN_data_out(8785),
        VN2CN2_bit => VN_data_out(8786),
        VN2CN3_bit => VN_data_out(8787),
        VN2CN4_bit => VN_data_out(8788),
        VN2CN5_bit => VN_data_out(8789),
        VN2CN0_sign => VN_sign_out(8784),
        VN2CN1_sign => VN_sign_out(8785),
        VN2CN2_sign => VN_sign_out(8786),
        VN2CN3_sign => VN_sign_out(8787),
        VN2CN4_sign => VN_sign_out(8788),
        VN2CN5_sign => VN_sign_out(8789),
        codeword => codeword(1464),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1465 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8795 downto 8790),
        Din0 => VN1465_in0,
        Din1 => VN1465_in1,
        Din2 => VN1465_in2,
        Din3 => VN1465_in3,
        Din4 => VN1465_in4,
        Din5 => VN1465_in5,
        VN2CN0_bit => VN_data_out(8790),
        VN2CN1_bit => VN_data_out(8791),
        VN2CN2_bit => VN_data_out(8792),
        VN2CN3_bit => VN_data_out(8793),
        VN2CN4_bit => VN_data_out(8794),
        VN2CN5_bit => VN_data_out(8795),
        VN2CN0_sign => VN_sign_out(8790),
        VN2CN1_sign => VN_sign_out(8791),
        VN2CN2_sign => VN_sign_out(8792),
        VN2CN3_sign => VN_sign_out(8793),
        VN2CN4_sign => VN_sign_out(8794),
        VN2CN5_sign => VN_sign_out(8795),
        codeword => codeword(1465),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1466 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8801 downto 8796),
        Din0 => VN1466_in0,
        Din1 => VN1466_in1,
        Din2 => VN1466_in2,
        Din3 => VN1466_in3,
        Din4 => VN1466_in4,
        Din5 => VN1466_in5,
        VN2CN0_bit => VN_data_out(8796),
        VN2CN1_bit => VN_data_out(8797),
        VN2CN2_bit => VN_data_out(8798),
        VN2CN3_bit => VN_data_out(8799),
        VN2CN4_bit => VN_data_out(8800),
        VN2CN5_bit => VN_data_out(8801),
        VN2CN0_sign => VN_sign_out(8796),
        VN2CN1_sign => VN_sign_out(8797),
        VN2CN2_sign => VN_sign_out(8798),
        VN2CN3_sign => VN_sign_out(8799),
        VN2CN4_sign => VN_sign_out(8800),
        VN2CN5_sign => VN_sign_out(8801),
        codeword => codeword(1466),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1467 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8807 downto 8802),
        Din0 => VN1467_in0,
        Din1 => VN1467_in1,
        Din2 => VN1467_in2,
        Din3 => VN1467_in3,
        Din4 => VN1467_in4,
        Din5 => VN1467_in5,
        VN2CN0_bit => VN_data_out(8802),
        VN2CN1_bit => VN_data_out(8803),
        VN2CN2_bit => VN_data_out(8804),
        VN2CN3_bit => VN_data_out(8805),
        VN2CN4_bit => VN_data_out(8806),
        VN2CN5_bit => VN_data_out(8807),
        VN2CN0_sign => VN_sign_out(8802),
        VN2CN1_sign => VN_sign_out(8803),
        VN2CN2_sign => VN_sign_out(8804),
        VN2CN3_sign => VN_sign_out(8805),
        VN2CN4_sign => VN_sign_out(8806),
        VN2CN5_sign => VN_sign_out(8807),
        codeword => codeword(1467),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1468 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8813 downto 8808),
        Din0 => VN1468_in0,
        Din1 => VN1468_in1,
        Din2 => VN1468_in2,
        Din3 => VN1468_in3,
        Din4 => VN1468_in4,
        Din5 => VN1468_in5,
        VN2CN0_bit => VN_data_out(8808),
        VN2CN1_bit => VN_data_out(8809),
        VN2CN2_bit => VN_data_out(8810),
        VN2CN3_bit => VN_data_out(8811),
        VN2CN4_bit => VN_data_out(8812),
        VN2CN5_bit => VN_data_out(8813),
        VN2CN0_sign => VN_sign_out(8808),
        VN2CN1_sign => VN_sign_out(8809),
        VN2CN2_sign => VN_sign_out(8810),
        VN2CN3_sign => VN_sign_out(8811),
        VN2CN4_sign => VN_sign_out(8812),
        VN2CN5_sign => VN_sign_out(8813),
        codeword => codeword(1468),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1469 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8819 downto 8814),
        Din0 => VN1469_in0,
        Din1 => VN1469_in1,
        Din2 => VN1469_in2,
        Din3 => VN1469_in3,
        Din4 => VN1469_in4,
        Din5 => VN1469_in5,
        VN2CN0_bit => VN_data_out(8814),
        VN2CN1_bit => VN_data_out(8815),
        VN2CN2_bit => VN_data_out(8816),
        VN2CN3_bit => VN_data_out(8817),
        VN2CN4_bit => VN_data_out(8818),
        VN2CN5_bit => VN_data_out(8819),
        VN2CN0_sign => VN_sign_out(8814),
        VN2CN1_sign => VN_sign_out(8815),
        VN2CN2_sign => VN_sign_out(8816),
        VN2CN3_sign => VN_sign_out(8817),
        VN2CN4_sign => VN_sign_out(8818),
        VN2CN5_sign => VN_sign_out(8819),
        codeword => codeword(1469),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1470 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8825 downto 8820),
        Din0 => VN1470_in0,
        Din1 => VN1470_in1,
        Din2 => VN1470_in2,
        Din3 => VN1470_in3,
        Din4 => VN1470_in4,
        Din5 => VN1470_in5,
        VN2CN0_bit => VN_data_out(8820),
        VN2CN1_bit => VN_data_out(8821),
        VN2CN2_bit => VN_data_out(8822),
        VN2CN3_bit => VN_data_out(8823),
        VN2CN4_bit => VN_data_out(8824),
        VN2CN5_bit => VN_data_out(8825),
        VN2CN0_sign => VN_sign_out(8820),
        VN2CN1_sign => VN_sign_out(8821),
        VN2CN2_sign => VN_sign_out(8822),
        VN2CN3_sign => VN_sign_out(8823),
        VN2CN4_sign => VN_sign_out(8824),
        VN2CN5_sign => VN_sign_out(8825),
        codeword => codeword(1470),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1471 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8831 downto 8826),
        Din0 => VN1471_in0,
        Din1 => VN1471_in1,
        Din2 => VN1471_in2,
        Din3 => VN1471_in3,
        Din4 => VN1471_in4,
        Din5 => VN1471_in5,
        VN2CN0_bit => VN_data_out(8826),
        VN2CN1_bit => VN_data_out(8827),
        VN2CN2_bit => VN_data_out(8828),
        VN2CN3_bit => VN_data_out(8829),
        VN2CN4_bit => VN_data_out(8830),
        VN2CN5_bit => VN_data_out(8831),
        VN2CN0_sign => VN_sign_out(8826),
        VN2CN1_sign => VN_sign_out(8827),
        VN2CN2_sign => VN_sign_out(8828),
        VN2CN3_sign => VN_sign_out(8829),
        VN2CN4_sign => VN_sign_out(8830),
        VN2CN5_sign => VN_sign_out(8831),
        codeword => codeword(1471),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1472 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8837 downto 8832),
        Din0 => VN1472_in0,
        Din1 => VN1472_in1,
        Din2 => VN1472_in2,
        Din3 => VN1472_in3,
        Din4 => VN1472_in4,
        Din5 => VN1472_in5,
        VN2CN0_bit => VN_data_out(8832),
        VN2CN1_bit => VN_data_out(8833),
        VN2CN2_bit => VN_data_out(8834),
        VN2CN3_bit => VN_data_out(8835),
        VN2CN4_bit => VN_data_out(8836),
        VN2CN5_bit => VN_data_out(8837),
        VN2CN0_sign => VN_sign_out(8832),
        VN2CN1_sign => VN_sign_out(8833),
        VN2CN2_sign => VN_sign_out(8834),
        VN2CN3_sign => VN_sign_out(8835),
        VN2CN4_sign => VN_sign_out(8836),
        VN2CN5_sign => VN_sign_out(8837),
        codeword => codeword(1472),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1473 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8843 downto 8838),
        Din0 => VN1473_in0,
        Din1 => VN1473_in1,
        Din2 => VN1473_in2,
        Din3 => VN1473_in3,
        Din4 => VN1473_in4,
        Din5 => VN1473_in5,
        VN2CN0_bit => VN_data_out(8838),
        VN2CN1_bit => VN_data_out(8839),
        VN2CN2_bit => VN_data_out(8840),
        VN2CN3_bit => VN_data_out(8841),
        VN2CN4_bit => VN_data_out(8842),
        VN2CN5_bit => VN_data_out(8843),
        VN2CN0_sign => VN_sign_out(8838),
        VN2CN1_sign => VN_sign_out(8839),
        VN2CN2_sign => VN_sign_out(8840),
        VN2CN3_sign => VN_sign_out(8841),
        VN2CN4_sign => VN_sign_out(8842),
        VN2CN5_sign => VN_sign_out(8843),
        codeword => codeword(1473),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1474 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8849 downto 8844),
        Din0 => VN1474_in0,
        Din1 => VN1474_in1,
        Din2 => VN1474_in2,
        Din3 => VN1474_in3,
        Din4 => VN1474_in4,
        Din5 => VN1474_in5,
        VN2CN0_bit => VN_data_out(8844),
        VN2CN1_bit => VN_data_out(8845),
        VN2CN2_bit => VN_data_out(8846),
        VN2CN3_bit => VN_data_out(8847),
        VN2CN4_bit => VN_data_out(8848),
        VN2CN5_bit => VN_data_out(8849),
        VN2CN0_sign => VN_sign_out(8844),
        VN2CN1_sign => VN_sign_out(8845),
        VN2CN2_sign => VN_sign_out(8846),
        VN2CN3_sign => VN_sign_out(8847),
        VN2CN4_sign => VN_sign_out(8848),
        VN2CN5_sign => VN_sign_out(8849),
        codeword => codeword(1474),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1475 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8855 downto 8850),
        Din0 => VN1475_in0,
        Din1 => VN1475_in1,
        Din2 => VN1475_in2,
        Din3 => VN1475_in3,
        Din4 => VN1475_in4,
        Din5 => VN1475_in5,
        VN2CN0_bit => VN_data_out(8850),
        VN2CN1_bit => VN_data_out(8851),
        VN2CN2_bit => VN_data_out(8852),
        VN2CN3_bit => VN_data_out(8853),
        VN2CN4_bit => VN_data_out(8854),
        VN2CN5_bit => VN_data_out(8855),
        VN2CN0_sign => VN_sign_out(8850),
        VN2CN1_sign => VN_sign_out(8851),
        VN2CN2_sign => VN_sign_out(8852),
        VN2CN3_sign => VN_sign_out(8853),
        VN2CN4_sign => VN_sign_out(8854),
        VN2CN5_sign => VN_sign_out(8855),
        codeword => codeword(1475),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1476 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8861 downto 8856),
        Din0 => VN1476_in0,
        Din1 => VN1476_in1,
        Din2 => VN1476_in2,
        Din3 => VN1476_in3,
        Din4 => VN1476_in4,
        Din5 => VN1476_in5,
        VN2CN0_bit => VN_data_out(8856),
        VN2CN1_bit => VN_data_out(8857),
        VN2CN2_bit => VN_data_out(8858),
        VN2CN3_bit => VN_data_out(8859),
        VN2CN4_bit => VN_data_out(8860),
        VN2CN5_bit => VN_data_out(8861),
        VN2CN0_sign => VN_sign_out(8856),
        VN2CN1_sign => VN_sign_out(8857),
        VN2CN2_sign => VN_sign_out(8858),
        VN2CN3_sign => VN_sign_out(8859),
        VN2CN4_sign => VN_sign_out(8860),
        VN2CN5_sign => VN_sign_out(8861),
        codeword => codeword(1476),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1477 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8867 downto 8862),
        Din0 => VN1477_in0,
        Din1 => VN1477_in1,
        Din2 => VN1477_in2,
        Din3 => VN1477_in3,
        Din4 => VN1477_in4,
        Din5 => VN1477_in5,
        VN2CN0_bit => VN_data_out(8862),
        VN2CN1_bit => VN_data_out(8863),
        VN2CN2_bit => VN_data_out(8864),
        VN2CN3_bit => VN_data_out(8865),
        VN2CN4_bit => VN_data_out(8866),
        VN2CN5_bit => VN_data_out(8867),
        VN2CN0_sign => VN_sign_out(8862),
        VN2CN1_sign => VN_sign_out(8863),
        VN2CN2_sign => VN_sign_out(8864),
        VN2CN3_sign => VN_sign_out(8865),
        VN2CN4_sign => VN_sign_out(8866),
        VN2CN5_sign => VN_sign_out(8867),
        codeword => codeword(1477),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1478 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8873 downto 8868),
        Din0 => VN1478_in0,
        Din1 => VN1478_in1,
        Din2 => VN1478_in2,
        Din3 => VN1478_in3,
        Din4 => VN1478_in4,
        Din5 => VN1478_in5,
        VN2CN0_bit => VN_data_out(8868),
        VN2CN1_bit => VN_data_out(8869),
        VN2CN2_bit => VN_data_out(8870),
        VN2CN3_bit => VN_data_out(8871),
        VN2CN4_bit => VN_data_out(8872),
        VN2CN5_bit => VN_data_out(8873),
        VN2CN0_sign => VN_sign_out(8868),
        VN2CN1_sign => VN_sign_out(8869),
        VN2CN2_sign => VN_sign_out(8870),
        VN2CN3_sign => VN_sign_out(8871),
        VN2CN4_sign => VN_sign_out(8872),
        VN2CN5_sign => VN_sign_out(8873),
        codeword => codeword(1478),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1479 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8879 downto 8874),
        Din0 => VN1479_in0,
        Din1 => VN1479_in1,
        Din2 => VN1479_in2,
        Din3 => VN1479_in3,
        Din4 => VN1479_in4,
        Din5 => VN1479_in5,
        VN2CN0_bit => VN_data_out(8874),
        VN2CN1_bit => VN_data_out(8875),
        VN2CN2_bit => VN_data_out(8876),
        VN2CN3_bit => VN_data_out(8877),
        VN2CN4_bit => VN_data_out(8878),
        VN2CN5_bit => VN_data_out(8879),
        VN2CN0_sign => VN_sign_out(8874),
        VN2CN1_sign => VN_sign_out(8875),
        VN2CN2_sign => VN_sign_out(8876),
        VN2CN3_sign => VN_sign_out(8877),
        VN2CN4_sign => VN_sign_out(8878),
        VN2CN5_sign => VN_sign_out(8879),
        codeword => codeword(1479),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1480 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8885 downto 8880),
        Din0 => VN1480_in0,
        Din1 => VN1480_in1,
        Din2 => VN1480_in2,
        Din3 => VN1480_in3,
        Din4 => VN1480_in4,
        Din5 => VN1480_in5,
        VN2CN0_bit => VN_data_out(8880),
        VN2CN1_bit => VN_data_out(8881),
        VN2CN2_bit => VN_data_out(8882),
        VN2CN3_bit => VN_data_out(8883),
        VN2CN4_bit => VN_data_out(8884),
        VN2CN5_bit => VN_data_out(8885),
        VN2CN0_sign => VN_sign_out(8880),
        VN2CN1_sign => VN_sign_out(8881),
        VN2CN2_sign => VN_sign_out(8882),
        VN2CN3_sign => VN_sign_out(8883),
        VN2CN4_sign => VN_sign_out(8884),
        VN2CN5_sign => VN_sign_out(8885),
        codeword => codeword(1480),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1481 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8891 downto 8886),
        Din0 => VN1481_in0,
        Din1 => VN1481_in1,
        Din2 => VN1481_in2,
        Din3 => VN1481_in3,
        Din4 => VN1481_in4,
        Din5 => VN1481_in5,
        VN2CN0_bit => VN_data_out(8886),
        VN2CN1_bit => VN_data_out(8887),
        VN2CN2_bit => VN_data_out(8888),
        VN2CN3_bit => VN_data_out(8889),
        VN2CN4_bit => VN_data_out(8890),
        VN2CN5_bit => VN_data_out(8891),
        VN2CN0_sign => VN_sign_out(8886),
        VN2CN1_sign => VN_sign_out(8887),
        VN2CN2_sign => VN_sign_out(8888),
        VN2CN3_sign => VN_sign_out(8889),
        VN2CN4_sign => VN_sign_out(8890),
        VN2CN5_sign => VN_sign_out(8891),
        codeword => codeword(1481),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1482 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8897 downto 8892),
        Din0 => VN1482_in0,
        Din1 => VN1482_in1,
        Din2 => VN1482_in2,
        Din3 => VN1482_in3,
        Din4 => VN1482_in4,
        Din5 => VN1482_in5,
        VN2CN0_bit => VN_data_out(8892),
        VN2CN1_bit => VN_data_out(8893),
        VN2CN2_bit => VN_data_out(8894),
        VN2CN3_bit => VN_data_out(8895),
        VN2CN4_bit => VN_data_out(8896),
        VN2CN5_bit => VN_data_out(8897),
        VN2CN0_sign => VN_sign_out(8892),
        VN2CN1_sign => VN_sign_out(8893),
        VN2CN2_sign => VN_sign_out(8894),
        VN2CN3_sign => VN_sign_out(8895),
        VN2CN4_sign => VN_sign_out(8896),
        VN2CN5_sign => VN_sign_out(8897),
        codeword => codeword(1482),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1483 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8903 downto 8898),
        Din0 => VN1483_in0,
        Din1 => VN1483_in1,
        Din2 => VN1483_in2,
        Din3 => VN1483_in3,
        Din4 => VN1483_in4,
        Din5 => VN1483_in5,
        VN2CN0_bit => VN_data_out(8898),
        VN2CN1_bit => VN_data_out(8899),
        VN2CN2_bit => VN_data_out(8900),
        VN2CN3_bit => VN_data_out(8901),
        VN2CN4_bit => VN_data_out(8902),
        VN2CN5_bit => VN_data_out(8903),
        VN2CN0_sign => VN_sign_out(8898),
        VN2CN1_sign => VN_sign_out(8899),
        VN2CN2_sign => VN_sign_out(8900),
        VN2CN3_sign => VN_sign_out(8901),
        VN2CN4_sign => VN_sign_out(8902),
        VN2CN5_sign => VN_sign_out(8903),
        codeword => codeword(1483),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1484 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8909 downto 8904),
        Din0 => VN1484_in0,
        Din1 => VN1484_in1,
        Din2 => VN1484_in2,
        Din3 => VN1484_in3,
        Din4 => VN1484_in4,
        Din5 => VN1484_in5,
        VN2CN0_bit => VN_data_out(8904),
        VN2CN1_bit => VN_data_out(8905),
        VN2CN2_bit => VN_data_out(8906),
        VN2CN3_bit => VN_data_out(8907),
        VN2CN4_bit => VN_data_out(8908),
        VN2CN5_bit => VN_data_out(8909),
        VN2CN0_sign => VN_sign_out(8904),
        VN2CN1_sign => VN_sign_out(8905),
        VN2CN2_sign => VN_sign_out(8906),
        VN2CN3_sign => VN_sign_out(8907),
        VN2CN4_sign => VN_sign_out(8908),
        VN2CN5_sign => VN_sign_out(8909),
        codeword => codeword(1484),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1485 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8915 downto 8910),
        Din0 => VN1485_in0,
        Din1 => VN1485_in1,
        Din2 => VN1485_in2,
        Din3 => VN1485_in3,
        Din4 => VN1485_in4,
        Din5 => VN1485_in5,
        VN2CN0_bit => VN_data_out(8910),
        VN2CN1_bit => VN_data_out(8911),
        VN2CN2_bit => VN_data_out(8912),
        VN2CN3_bit => VN_data_out(8913),
        VN2CN4_bit => VN_data_out(8914),
        VN2CN5_bit => VN_data_out(8915),
        VN2CN0_sign => VN_sign_out(8910),
        VN2CN1_sign => VN_sign_out(8911),
        VN2CN2_sign => VN_sign_out(8912),
        VN2CN3_sign => VN_sign_out(8913),
        VN2CN4_sign => VN_sign_out(8914),
        VN2CN5_sign => VN_sign_out(8915),
        codeword => codeword(1485),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1486 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8921 downto 8916),
        Din0 => VN1486_in0,
        Din1 => VN1486_in1,
        Din2 => VN1486_in2,
        Din3 => VN1486_in3,
        Din4 => VN1486_in4,
        Din5 => VN1486_in5,
        VN2CN0_bit => VN_data_out(8916),
        VN2CN1_bit => VN_data_out(8917),
        VN2CN2_bit => VN_data_out(8918),
        VN2CN3_bit => VN_data_out(8919),
        VN2CN4_bit => VN_data_out(8920),
        VN2CN5_bit => VN_data_out(8921),
        VN2CN0_sign => VN_sign_out(8916),
        VN2CN1_sign => VN_sign_out(8917),
        VN2CN2_sign => VN_sign_out(8918),
        VN2CN3_sign => VN_sign_out(8919),
        VN2CN4_sign => VN_sign_out(8920),
        VN2CN5_sign => VN_sign_out(8921),
        codeword => codeword(1486),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1487 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8927 downto 8922),
        Din0 => VN1487_in0,
        Din1 => VN1487_in1,
        Din2 => VN1487_in2,
        Din3 => VN1487_in3,
        Din4 => VN1487_in4,
        Din5 => VN1487_in5,
        VN2CN0_bit => VN_data_out(8922),
        VN2CN1_bit => VN_data_out(8923),
        VN2CN2_bit => VN_data_out(8924),
        VN2CN3_bit => VN_data_out(8925),
        VN2CN4_bit => VN_data_out(8926),
        VN2CN5_bit => VN_data_out(8927),
        VN2CN0_sign => VN_sign_out(8922),
        VN2CN1_sign => VN_sign_out(8923),
        VN2CN2_sign => VN_sign_out(8924),
        VN2CN3_sign => VN_sign_out(8925),
        VN2CN4_sign => VN_sign_out(8926),
        VN2CN5_sign => VN_sign_out(8927),
        codeword => codeword(1487),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1488 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8933 downto 8928),
        Din0 => VN1488_in0,
        Din1 => VN1488_in1,
        Din2 => VN1488_in2,
        Din3 => VN1488_in3,
        Din4 => VN1488_in4,
        Din5 => VN1488_in5,
        VN2CN0_bit => VN_data_out(8928),
        VN2CN1_bit => VN_data_out(8929),
        VN2CN2_bit => VN_data_out(8930),
        VN2CN3_bit => VN_data_out(8931),
        VN2CN4_bit => VN_data_out(8932),
        VN2CN5_bit => VN_data_out(8933),
        VN2CN0_sign => VN_sign_out(8928),
        VN2CN1_sign => VN_sign_out(8929),
        VN2CN2_sign => VN_sign_out(8930),
        VN2CN3_sign => VN_sign_out(8931),
        VN2CN4_sign => VN_sign_out(8932),
        VN2CN5_sign => VN_sign_out(8933),
        codeword => codeword(1488),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1489 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8939 downto 8934),
        Din0 => VN1489_in0,
        Din1 => VN1489_in1,
        Din2 => VN1489_in2,
        Din3 => VN1489_in3,
        Din4 => VN1489_in4,
        Din5 => VN1489_in5,
        VN2CN0_bit => VN_data_out(8934),
        VN2CN1_bit => VN_data_out(8935),
        VN2CN2_bit => VN_data_out(8936),
        VN2CN3_bit => VN_data_out(8937),
        VN2CN4_bit => VN_data_out(8938),
        VN2CN5_bit => VN_data_out(8939),
        VN2CN0_sign => VN_sign_out(8934),
        VN2CN1_sign => VN_sign_out(8935),
        VN2CN2_sign => VN_sign_out(8936),
        VN2CN3_sign => VN_sign_out(8937),
        VN2CN4_sign => VN_sign_out(8938),
        VN2CN5_sign => VN_sign_out(8939),
        codeword => codeword(1489),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1490 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8945 downto 8940),
        Din0 => VN1490_in0,
        Din1 => VN1490_in1,
        Din2 => VN1490_in2,
        Din3 => VN1490_in3,
        Din4 => VN1490_in4,
        Din5 => VN1490_in5,
        VN2CN0_bit => VN_data_out(8940),
        VN2CN1_bit => VN_data_out(8941),
        VN2CN2_bit => VN_data_out(8942),
        VN2CN3_bit => VN_data_out(8943),
        VN2CN4_bit => VN_data_out(8944),
        VN2CN5_bit => VN_data_out(8945),
        VN2CN0_sign => VN_sign_out(8940),
        VN2CN1_sign => VN_sign_out(8941),
        VN2CN2_sign => VN_sign_out(8942),
        VN2CN3_sign => VN_sign_out(8943),
        VN2CN4_sign => VN_sign_out(8944),
        VN2CN5_sign => VN_sign_out(8945),
        codeword => codeword(1490),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1491 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8951 downto 8946),
        Din0 => VN1491_in0,
        Din1 => VN1491_in1,
        Din2 => VN1491_in2,
        Din3 => VN1491_in3,
        Din4 => VN1491_in4,
        Din5 => VN1491_in5,
        VN2CN0_bit => VN_data_out(8946),
        VN2CN1_bit => VN_data_out(8947),
        VN2CN2_bit => VN_data_out(8948),
        VN2CN3_bit => VN_data_out(8949),
        VN2CN4_bit => VN_data_out(8950),
        VN2CN5_bit => VN_data_out(8951),
        VN2CN0_sign => VN_sign_out(8946),
        VN2CN1_sign => VN_sign_out(8947),
        VN2CN2_sign => VN_sign_out(8948),
        VN2CN3_sign => VN_sign_out(8949),
        VN2CN4_sign => VN_sign_out(8950),
        VN2CN5_sign => VN_sign_out(8951),
        codeword => codeword(1491),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1492 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8957 downto 8952),
        Din0 => VN1492_in0,
        Din1 => VN1492_in1,
        Din2 => VN1492_in2,
        Din3 => VN1492_in3,
        Din4 => VN1492_in4,
        Din5 => VN1492_in5,
        VN2CN0_bit => VN_data_out(8952),
        VN2CN1_bit => VN_data_out(8953),
        VN2CN2_bit => VN_data_out(8954),
        VN2CN3_bit => VN_data_out(8955),
        VN2CN4_bit => VN_data_out(8956),
        VN2CN5_bit => VN_data_out(8957),
        VN2CN0_sign => VN_sign_out(8952),
        VN2CN1_sign => VN_sign_out(8953),
        VN2CN2_sign => VN_sign_out(8954),
        VN2CN3_sign => VN_sign_out(8955),
        VN2CN4_sign => VN_sign_out(8956),
        VN2CN5_sign => VN_sign_out(8957),
        codeword => codeword(1492),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1493 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8963 downto 8958),
        Din0 => VN1493_in0,
        Din1 => VN1493_in1,
        Din2 => VN1493_in2,
        Din3 => VN1493_in3,
        Din4 => VN1493_in4,
        Din5 => VN1493_in5,
        VN2CN0_bit => VN_data_out(8958),
        VN2CN1_bit => VN_data_out(8959),
        VN2CN2_bit => VN_data_out(8960),
        VN2CN3_bit => VN_data_out(8961),
        VN2CN4_bit => VN_data_out(8962),
        VN2CN5_bit => VN_data_out(8963),
        VN2CN0_sign => VN_sign_out(8958),
        VN2CN1_sign => VN_sign_out(8959),
        VN2CN2_sign => VN_sign_out(8960),
        VN2CN3_sign => VN_sign_out(8961),
        VN2CN4_sign => VN_sign_out(8962),
        VN2CN5_sign => VN_sign_out(8963),
        codeword => codeword(1493),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1494 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8969 downto 8964),
        Din0 => VN1494_in0,
        Din1 => VN1494_in1,
        Din2 => VN1494_in2,
        Din3 => VN1494_in3,
        Din4 => VN1494_in4,
        Din5 => VN1494_in5,
        VN2CN0_bit => VN_data_out(8964),
        VN2CN1_bit => VN_data_out(8965),
        VN2CN2_bit => VN_data_out(8966),
        VN2CN3_bit => VN_data_out(8967),
        VN2CN4_bit => VN_data_out(8968),
        VN2CN5_bit => VN_data_out(8969),
        VN2CN0_sign => VN_sign_out(8964),
        VN2CN1_sign => VN_sign_out(8965),
        VN2CN2_sign => VN_sign_out(8966),
        VN2CN3_sign => VN_sign_out(8967),
        VN2CN4_sign => VN_sign_out(8968),
        VN2CN5_sign => VN_sign_out(8969),
        codeword => codeword(1494),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1495 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8975 downto 8970),
        Din0 => VN1495_in0,
        Din1 => VN1495_in1,
        Din2 => VN1495_in2,
        Din3 => VN1495_in3,
        Din4 => VN1495_in4,
        Din5 => VN1495_in5,
        VN2CN0_bit => VN_data_out(8970),
        VN2CN1_bit => VN_data_out(8971),
        VN2CN2_bit => VN_data_out(8972),
        VN2CN3_bit => VN_data_out(8973),
        VN2CN4_bit => VN_data_out(8974),
        VN2CN5_bit => VN_data_out(8975),
        VN2CN0_sign => VN_sign_out(8970),
        VN2CN1_sign => VN_sign_out(8971),
        VN2CN2_sign => VN_sign_out(8972),
        VN2CN3_sign => VN_sign_out(8973),
        VN2CN4_sign => VN_sign_out(8974),
        VN2CN5_sign => VN_sign_out(8975),
        codeword => codeword(1495),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1496 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8981 downto 8976),
        Din0 => VN1496_in0,
        Din1 => VN1496_in1,
        Din2 => VN1496_in2,
        Din3 => VN1496_in3,
        Din4 => VN1496_in4,
        Din5 => VN1496_in5,
        VN2CN0_bit => VN_data_out(8976),
        VN2CN1_bit => VN_data_out(8977),
        VN2CN2_bit => VN_data_out(8978),
        VN2CN3_bit => VN_data_out(8979),
        VN2CN4_bit => VN_data_out(8980),
        VN2CN5_bit => VN_data_out(8981),
        VN2CN0_sign => VN_sign_out(8976),
        VN2CN1_sign => VN_sign_out(8977),
        VN2CN2_sign => VN_sign_out(8978),
        VN2CN3_sign => VN_sign_out(8979),
        VN2CN4_sign => VN_sign_out(8980),
        VN2CN5_sign => VN_sign_out(8981),
        codeword => codeword(1496),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1497 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8987 downto 8982),
        Din0 => VN1497_in0,
        Din1 => VN1497_in1,
        Din2 => VN1497_in2,
        Din3 => VN1497_in3,
        Din4 => VN1497_in4,
        Din5 => VN1497_in5,
        VN2CN0_bit => VN_data_out(8982),
        VN2CN1_bit => VN_data_out(8983),
        VN2CN2_bit => VN_data_out(8984),
        VN2CN3_bit => VN_data_out(8985),
        VN2CN4_bit => VN_data_out(8986),
        VN2CN5_bit => VN_data_out(8987),
        VN2CN0_sign => VN_sign_out(8982),
        VN2CN1_sign => VN_sign_out(8983),
        VN2CN2_sign => VN_sign_out(8984),
        VN2CN3_sign => VN_sign_out(8985),
        VN2CN4_sign => VN_sign_out(8986),
        VN2CN5_sign => VN_sign_out(8987),
        codeword => codeword(1497),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1498 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8993 downto 8988),
        Din0 => VN1498_in0,
        Din1 => VN1498_in1,
        Din2 => VN1498_in2,
        Din3 => VN1498_in3,
        Din4 => VN1498_in4,
        Din5 => VN1498_in5,
        VN2CN0_bit => VN_data_out(8988),
        VN2CN1_bit => VN_data_out(8989),
        VN2CN2_bit => VN_data_out(8990),
        VN2CN3_bit => VN_data_out(8991),
        VN2CN4_bit => VN_data_out(8992),
        VN2CN5_bit => VN_data_out(8993),
        VN2CN0_sign => VN_sign_out(8988),
        VN2CN1_sign => VN_sign_out(8989),
        VN2CN2_sign => VN_sign_out(8990),
        VN2CN3_sign => VN_sign_out(8991),
        VN2CN4_sign => VN_sign_out(8992),
        VN2CN5_sign => VN_sign_out(8993),
        codeword => codeword(1498),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1499 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(8999 downto 8994),
        Din0 => VN1499_in0,
        Din1 => VN1499_in1,
        Din2 => VN1499_in2,
        Din3 => VN1499_in3,
        Din4 => VN1499_in4,
        Din5 => VN1499_in5,
        VN2CN0_bit => VN_data_out(8994),
        VN2CN1_bit => VN_data_out(8995),
        VN2CN2_bit => VN_data_out(8996),
        VN2CN3_bit => VN_data_out(8997),
        VN2CN4_bit => VN_data_out(8998),
        VN2CN5_bit => VN_data_out(8999),
        VN2CN0_sign => VN_sign_out(8994),
        VN2CN1_sign => VN_sign_out(8995),
        VN2CN2_sign => VN_sign_out(8996),
        VN2CN3_sign => VN_sign_out(8997),
        VN2CN4_sign => VN_sign_out(8998),
        VN2CN5_sign => VN_sign_out(8999),
        codeword => codeword(1499),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1500 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9005 downto 9000),
        Din0 => VN1500_in0,
        Din1 => VN1500_in1,
        Din2 => VN1500_in2,
        Din3 => VN1500_in3,
        Din4 => VN1500_in4,
        Din5 => VN1500_in5,
        VN2CN0_bit => VN_data_out(9000),
        VN2CN1_bit => VN_data_out(9001),
        VN2CN2_bit => VN_data_out(9002),
        VN2CN3_bit => VN_data_out(9003),
        VN2CN4_bit => VN_data_out(9004),
        VN2CN5_bit => VN_data_out(9005),
        VN2CN0_sign => VN_sign_out(9000),
        VN2CN1_sign => VN_sign_out(9001),
        VN2CN2_sign => VN_sign_out(9002),
        VN2CN3_sign => VN_sign_out(9003),
        VN2CN4_sign => VN_sign_out(9004),
        VN2CN5_sign => VN_sign_out(9005),
        codeword => codeword(1500),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1501 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9011 downto 9006),
        Din0 => VN1501_in0,
        Din1 => VN1501_in1,
        Din2 => VN1501_in2,
        Din3 => VN1501_in3,
        Din4 => VN1501_in4,
        Din5 => VN1501_in5,
        VN2CN0_bit => VN_data_out(9006),
        VN2CN1_bit => VN_data_out(9007),
        VN2CN2_bit => VN_data_out(9008),
        VN2CN3_bit => VN_data_out(9009),
        VN2CN4_bit => VN_data_out(9010),
        VN2CN5_bit => VN_data_out(9011),
        VN2CN0_sign => VN_sign_out(9006),
        VN2CN1_sign => VN_sign_out(9007),
        VN2CN2_sign => VN_sign_out(9008),
        VN2CN3_sign => VN_sign_out(9009),
        VN2CN4_sign => VN_sign_out(9010),
        VN2CN5_sign => VN_sign_out(9011),
        codeword => codeword(1501),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1502 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9017 downto 9012),
        Din0 => VN1502_in0,
        Din1 => VN1502_in1,
        Din2 => VN1502_in2,
        Din3 => VN1502_in3,
        Din4 => VN1502_in4,
        Din5 => VN1502_in5,
        VN2CN0_bit => VN_data_out(9012),
        VN2CN1_bit => VN_data_out(9013),
        VN2CN2_bit => VN_data_out(9014),
        VN2CN3_bit => VN_data_out(9015),
        VN2CN4_bit => VN_data_out(9016),
        VN2CN5_bit => VN_data_out(9017),
        VN2CN0_sign => VN_sign_out(9012),
        VN2CN1_sign => VN_sign_out(9013),
        VN2CN2_sign => VN_sign_out(9014),
        VN2CN3_sign => VN_sign_out(9015),
        VN2CN4_sign => VN_sign_out(9016),
        VN2CN5_sign => VN_sign_out(9017),
        codeword => codeword(1502),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1503 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9023 downto 9018),
        Din0 => VN1503_in0,
        Din1 => VN1503_in1,
        Din2 => VN1503_in2,
        Din3 => VN1503_in3,
        Din4 => VN1503_in4,
        Din5 => VN1503_in5,
        VN2CN0_bit => VN_data_out(9018),
        VN2CN1_bit => VN_data_out(9019),
        VN2CN2_bit => VN_data_out(9020),
        VN2CN3_bit => VN_data_out(9021),
        VN2CN4_bit => VN_data_out(9022),
        VN2CN5_bit => VN_data_out(9023),
        VN2CN0_sign => VN_sign_out(9018),
        VN2CN1_sign => VN_sign_out(9019),
        VN2CN2_sign => VN_sign_out(9020),
        VN2CN3_sign => VN_sign_out(9021),
        VN2CN4_sign => VN_sign_out(9022),
        VN2CN5_sign => VN_sign_out(9023),
        codeword => codeword(1503),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1504 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9029 downto 9024),
        Din0 => VN1504_in0,
        Din1 => VN1504_in1,
        Din2 => VN1504_in2,
        Din3 => VN1504_in3,
        Din4 => VN1504_in4,
        Din5 => VN1504_in5,
        VN2CN0_bit => VN_data_out(9024),
        VN2CN1_bit => VN_data_out(9025),
        VN2CN2_bit => VN_data_out(9026),
        VN2CN3_bit => VN_data_out(9027),
        VN2CN4_bit => VN_data_out(9028),
        VN2CN5_bit => VN_data_out(9029),
        VN2CN0_sign => VN_sign_out(9024),
        VN2CN1_sign => VN_sign_out(9025),
        VN2CN2_sign => VN_sign_out(9026),
        VN2CN3_sign => VN_sign_out(9027),
        VN2CN4_sign => VN_sign_out(9028),
        VN2CN5_sign => VN_sign_out(9029),
        codeword => codeword(1504),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1505 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9035 downto 9030),
        Din0 => VN1505_in0,
        Din1 => VN1505_in1,
        Din2 => VN1505_in2,
        Din3 => VN1505_in3,
        Din4 => VN1505_in4,
        Din5 => VN1505_in5,
        VN2CN0_bit => VN_data_out(9030),
        VN2CN1_bit => VN_data_out(9031),
        VN2CN2_bit => VN_data_out(9032),
        VN2CN3_bit => VN_data_out(9033),
        VN2CN4_bit => VN_data_out(9034),
        VN2CN5_bit => VN_data_out(9035),
        VN2CN0_sign => VN_sign_out(9030),
        VN2CN1_sign => VN_sign_out(9031),
        VN2CN2_sign => VN_sign_out(9032),
        VN2CN3_sign => VN_sign_out(9033),
        VN2CN4_sign => VN_sign_out(9034),
        VN2CN5_sign => VN_sign_out(9035),
        codeword => codeword(1505),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1506 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9041 downto 9036),
        Din0 => VN1506_in0,
        Din1 => VN1506_in1,
        Din2 => VN1506_in2,
        Din3 => VN1506_in3,
        Din4 => VN1506_in4,
        Din5 => VN1506_in5,
        VN2CN0_bit => VN_data_out(9036),
        VN2CN1_bit => VN_data_out(9037),
        VN2CN2_bit => VN_data_out(9038),
        VN2CN3_bit => VN_data_out(9039),
        VN2CN4_bit => VN_data_out(9040),
        VN2CN5_bit => VN_data_out(9041),
        VN2CN0_sign => VN_sign_out(9036),
        VN2CN1_sign => VN_sign_out(9037),
        VN2CN2_sign => VN_sign_out(9038),
        VN2CN3_sign => VN_sign_out(9039),
        VN2CN4_sign => VN_sign_out(9040),
        VN2CN5_sign => VN_sign_out(9041),
        codeword => codeword(1506),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1507 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9047 downto 9042),
        Din0 => VN1507_in0,
        Din1 => VN1507_in1,
        Din2 => VN1507_in2,
        Din3 => VN1507_in3,
        Din4 => VN1507_in4,
        Din5 => VN1507_in5,
        VN2CN0_bit => VN_data_out(9042),
        VN2CN1_bit => VN_data_out(9043),
        VN2CN2_bit => VN_data_out(9044),
        VN2CN3_bit => VN_data_out(9045),
        VN2CN4_bit => VN_data_out(9046),
        VN2CN5_bit => VN_data_out(9047),
        VN2CN0_sign => VN_sign_out(9042),
        VN2CN1_sign => VN_sign_out(9043),
        VN2CN2_sign => VN_sign_out(9044),
        VN2CN3_sign => VN_sign_out(9045),
        VN2CN4_sign => VN_sign_out(9046),
        VN2CN5_sign => VN_sign_out(9047),
        codeword => codeword(1507),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1508 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9053 downto 9048),
        Din0 => VN1508_in0,
        Din1 => VN1508_in1,
        Din2 => VN1508_in2,
        Din3 => VN1508_in3,
        Din4 => VN1508_in4,
        Din5 => VN1508_in5,
        VN2CN0_bit => VN_data_out(9048),
        VN2CN1_bit => VN_data_out(9049),
        VN2CN2_bit => VN_data_out(9050),
        VN2CN3_bit => VN_data_out(9051),
        VN2CN4_bit => VN_data_out(9052),
        VN2CN5_bit => VN_data_out(9053),
        VN2CN0_sign => VN_sign_out(9048),
        VN2CN1_sign => VN_sign_out(9049),
        VN2CN2_sign => VN_sign_out(9050),
        VN2CN3_sign => VN_sign_out(9051),
        VN2CN4_sign => VN_sign_out(9052),
        VN2CN5_sign => VN_sign_out(9053),
        codeword => codeword(1508),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1509 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9059 downto 9054),
        Din0 => VN1509_in0,
        Din1 => VN1509_in1,
        Din2 => VN1509_in2,
        Din3 => VN1509_in3,
        Din4 => VN1509_in4,
        Din5 => VN1509_in5,
        VN2CN0_bit => VN_data_out(9054),
        VN2CN1_bit => VN_data_out(9055),
        VN2CN2_bit => VN_data_out(9056),
        VN2CN3_bit => VN_data_out(9057),
        VN2CN4_bit => VN_data_out(9058),
        VN2CN5_bit => VN_data_out(9059),
        VN2CN0_sign => VN_sign_out(9054),
        VN2CN1_sign => VN_sign_out(9055),
        VN2CN2_sign => VN_sign_out(9056),
        VN2CN3_sign => VN_sign_out(9057),
        VN2CN4_sign => VN_sign_out(9058),
        VN2CN5_sign => VN_sign_out(9059),
        codeword => codeword(1509),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1510 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9065 downto 9060),
        Din0 => VN1510_in0,
        Din1 => VN1510_in1,
        Din2 => VN1510_in2,
        Din3 => VN1510_in3,
        Din4 => VN1510_in4,
        Din5 => VN1510_in5,
        VN2CN0_bit => VN_data_out(9060),
        VN2CN1_bit => VN_data_out(9061),
        VN2CN2_bit => VN_data_out(9062),
        VN2CN3_bit => VN_data_out(9063),
        VN2CN4_bit => VN_data_out(9064),
        VN2CN5_bit => VN_data_out(9065),
        VN2CN0_sign => VN_sign_out(9060),
        VN2CN1_sign => VN_sign_out(9061),
        VN2CN2_sign => VN_sign_out(9062),
        VN2CN3_sign => VN_sign_out(9063),
        VN2CN4_sign => VN_sign_out(9064),
        VN2CN5_sign => VN_sign_out(9065),
        codeword => codeword(1510),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1511 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9071 downto 9066),
        Din0 => VN1511_in0,
        Din1 => VN1511_in1,
        Din2 => VN1511_in2,
        Din3 => VN1511_in3,
        Din4 => VN1511_in4,
        Din5 => VN1511_in5,
        VN2CN0_bit => VN_data_out(9066),
        VN2CN1_bit => VN_data_out(9067),
        VN2CN2_bit => VN_data_out(9068),
        VN2CN3_bit => VN_data_out(9069),
        VN2CN4_bit => VN_data_out(9070),
        VN2CN5_bit => VN_data_out(9071),
        VN2CN0_sign => VN_sign_out(9066),
        VN2CN1_sign => VN_sign_out(9067),
        VN2CN2_sign => VN_sign_out(9068),
        VN2CN3_sign => VN_sign_out(9069),
        VN2CN4_sign => VN_sign_out(9070),
        VN2CN5_sign => VN_sign_out(9071),
        codeword => codeword(1511),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1512 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9077 downto 9072),
        Din0 => VN1512_in0,
        Din1 => VN1512_in1,
        Din2 => VN1512_in2,
        Din3 => VN1512_in3,
        Din4 => VN1512_in4,
        Din5 => VN1512_in5,
        VN2CN0_bit => VN_data_out(9072),
        VN2CN1_bit => VN_data_out(9073),
        VN2CN2_bit => VN_data_out(9074),
        VN2CN3_bit => VN_data_out(9075),
        VN2CN4_bit => VN_data_out(9076),
        VN2CN5_bit => VN_data_out(9077),
        VN2CN0_sign => VN_sign_out(9072),
        VN2CN1_sign => VN_sign_out(9073),
        VN2CN2_sign => VN_sign_out(9074),
        VN2CN3_sign => VN_sign_out(9075),
        VN2CN4_sign => VN_sign_out(9076),
        VN2CN5_sign => VN_sign_out(9077),
        codeword => codeword(1512),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1513 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9083 downto 9078),
        Din0 => VN1513_in0,
        Din1 => VN1513_in1,
        Din2 => VN1513_in2,
        Din3 => VN1513_in3,
        Din4 => VN1513_in4,
        Din5 => VN1513_in5,
        VN2CN0_bit => VN_data_out(9078),
        VN2CN1_bit => VN_data_out(9079),
        VN2CN2_bit => VN_data_out(9080),
        VN2CN3_bit => VN_data_out(9081),
        VN2CN4_bit => VN_data_out(9082),
        VN2CN5_bit => VN_data_out(9083),
        VN2CN0_sign => VN_sign_out(9078),
        VN2CN1_sign => VN_sign_out(9079),
        VN2CN2_sign => VN_sign_out(9080),
        VN2CN3_sign => VN_sign_out(9081),
        VN2CN4_sign => VN_sign_out(9082),
        VN2CN5_sign => VN_sign_out(9083),
        codeword => codeword(1513),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1514 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9089 downto 9084),
        Din0 => VN1514_in0,
        Din1 => VN1514_in1,
        Din2 => VN1514_in2,
        Din3 => VN1514_in3,
        Din4 => VN1514_in4,
        Din5 => VN1514_in5,
        VN2CN0_bit => VN_data_out(9084),
        VN2CN1_bit => VN_data_out(9085),
        VN2CN2_bit => VN_data_out(9086),
        VN2CN3_bit => VN_data_out(9087),
        VN2CN4_bit => VN_data_out(9088),
        VN2CN5_bit => VN_data_out(9089),
        VN2CN0_sign => VN_sign_out(9084),
        VN2CN1_sign => VN_sign_out(9085),
        VN2CN2_sign => VN_sign_out(9086),
        VN2CN3_sign => VN_sign_out(9087),
        VN2CN4_sign => VN_sign_out(9088),
        VN2CN5_sign => VN_sign_out(9089),
        codeword => codeword(1514),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1515 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9095 downto 9090),
        Din0 => VN1515_in0,
        Din1 => VN1515_in1,
        Din2 => VN1515_in2,
        Din3 => VN1515_in3,
        Din4 => VN1515_in4,
        Din5 => VN1515_in5,
        VN2CN0_bit => VN_data_out(9090),
        VN2CN1_bit => VN_data_out(9091),
        VN2CN2_bit => VN_data_out(9092),
        VN2CN3_bit => VN_data_out(9093),
        VN2CN4_bit => VN_data_out(9094),
        VN2CN5_bit => VN_data_out(9095),
        VN2CN0_sign => VN_sign_out(9090),
        VN2CN1_sign => VN_sign_out(9091),
        VN2CN2_sign => VN_sign_out(9092),
        VN2CN3_sign => VN_sign_out(9093),
        VN2CN4_sign => VN_sign_out(9094),
        VN2CN5_sign => VN_sign_out(9095),
        codeword => codeword(1515),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1516 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9101 downto 9096),
        Din0 => VN1516_in0,
        Din1 => VN1516_in1,
        Din2 => VN1516_in2,
        Din3 => VN1516_in3,
        Din4 => VN1516_in4,
        Din5 => VN1516_in5,
        VN2CN0_bit => VN_data_out(9096),
        VN2CN1_bit => VN_data_out(9097),
        VN2CN2_bit => VN_data_out(9098),
        VN2CN3_bit => VN_data_out(9099),
        VN2CN4_bit => VN_data_out(9100),
        VN2CN5_bit => VN_data_out(9101),
        VN2CN0_sign => VN_sign_out(9096),
        VN2CN1_sign => VN_sign_out(9097),
        VN2CN2_sign => VN_sign_out(9098),
        VN2CN3_sign => VN_sign_out(9099),
        VN2CN4_sign => VN_sign_out(9100),
        VN2CN5_sign => VN_sign_out(9101),
        codeword => codeword(1516),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1517 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9107 downto 9102),
        Din0 => VN1517_in0,
        Din1 => VN1517_in1,
        Din2 => VN1517_in2,
        Din3 => VN1517_in3,
        Din4 => VN1517_in4,
        Din5 => VN1517_in5,
        VN2CN0_bit => VN_data_out(9102),
        VN2CN1_bit => VN_data_out(9103),
        VN2CN2_bit => VN_data_out(9104),
        VN2CN3_bit => VN_data_out(9105),
        VN2CN4_bit => VN_data_out(9106),
        VN2CN5_bit => VN_data_out(9107),
        VN2CN0_sign => VN_sign_out(9102),
        VN2CN1_sign => VN_sign_out(9103),
        VN2CN2_sign => VN_sign_out(9104),
        VN2CN3_sign => VN_sign_out(9105),
        VN2CN4_sign => VN_sign_out(9106),
        VN2CN5_sign => VN_sign_out(9107),
        codeword => codeword(1517),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1518 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9113 downto 9108),
        Din0 => VN1518_in0,
        Din1 => VN1518_in1,
        Din2 => VN1518_in2,
        Din3 => VN1518_in3,
        Din4 => VN1518_in4,
        Din5 => VN1518_in5,
        VN2CN0_bit => VN_data_out(9108),
        VN2CN1_bit => VN_data_out(9109),
        VN2CN2_bit => VN_data_out(9110),
        VN2CN3_bit => VN_data_out(9111),
        VN2CN4_bit => VN_data_out(9112),
        VN2CN5_bit => VN_data_out(9113),
        VN2CN0_sign => VN_sign_out(9108),
        VN2CN1_sign => VN_sign_out(9109),
        VN2CN2_sign => VN_sign_out(9110),
        VN2CN3_sign => VN_sign_out(9111),
        VN2CN4_sign => VN_sign_out(9112),
        VN2CN5_sign => VN_sign_out(9113),
        codeword => codeword(1518),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1519 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9119 downto 9114),
        Din0 => VN1519_in0,
        Din1 => VN1519_in1,
        Din2 => VN1519_in2,
        Din3 => VN1519_in3,
        Din4 => VN1519_in4,
        Din5 => VN1519_in5,
        VN2CN0_bit => VN_data_out(9114),
        VN2CN1_bit => VN_data_out(9115),
        VN2CN2_bit => VN_data_out(9116),
        VN2CN3_bit => VN_data_out(9117),
        VN2CN4_bit => VN_data_out(9118),
        VN2CN5_bit => VN_data_out(9119),
        VN2CN0_sign => VN_sign_out(9114),
        VN2CN1_sign => VN_sign_out(9115),
        VN2CN2_sign => VN_sign_out(9116),
        VN2CN3_sign => VN_sign_out(9117),
        VN2CN4_sign => VN_sign_out(9118),
        VN2CN5_sign => VN_sign_out(9119),
        codeword => codeword(1519),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1520 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9125 downto 9120),
        Din0 => VN1520_in0,
        Din1 => VN1520_in1,
        Din2 => VN1520_in2,
        Din3 => VN1520_in3,
        Din4 => VN1520_in4,
        Din5 => VN1520_in5,
        VN2CN0_bit => VN_data_out(9120),
        VN2CN1_bit => VN_data_out(9121),
        VN2CN2_bit => VN_data_out(9122),
        VN2CN3_bit => VN_data_out(9123),
        VN2CN4_bit => VN_data_out(9124),
        VN2CN5_bit => VN_data_out(9125),
        VN2CN0_sign => VN_sign_out(9120),
        VN2CN1_sign => VN_sign_out(9121),
        VN2CN2_sign => VN_sign_out(9122),
        VN2CN3_sign => VN_sign_out(9123),
        VN2CN4_sign => VN_sign_out(9124),
        VN2CN5_sign => VN_sign_out(9125),
        codeword => codeword(1520),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1521 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9131 downto 9126),
        Din0 => VN1521_in0,
        Din1 => VN1521_in1,
        Din2 => VN1521_in2,
        Din3 => VN1521_in3,
        Din4 => VN1521_in4,
        Din5 => VN1521_in5,
        VN2CN0_bit => VN_data_out(9126),
        VN2CN1_bit => VN_data_out(9127),
        VN2CN2_bit => VN_data_out(9128),
        VN2CN3_bit => VN_data_out(9129),
        VN2CN4_bit => VN_data_out(9130),
        VN2CN5_bit => VN_data_out(9131),
        VN2CN0_sign => VN_sign_out(9126),
        VN2CN1_sign => VN_sign_out(9127),
        VN2CN2_sign => VN_sign_out(9128),
        VN2CN3_sign => VN_sign_out(9129),
        VN2CN4_sign => VN_sign_out(9130),
        VN2CN5_sign => VN_sign_out(9131),
        codeword => codeword(1521),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1522 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9137 downto 9132),
        Din0 => VN1522_in0,
        Din1 => VN1522_in1,
        Din2 => VN1522_in2,
        Din3 => VN1522_in3,
        Din4 => VN1522_in4,
        Din5 => VN1522_in5,
        VN2CN0_bit => VN_data_out(9132),
        VN2CN1_bit => VN_data_out(9133),
        VN2CN2_bit => VN_data_out(9134),
        VN2CN3_bit => VN_data_out(9135),
        VN2CN4_bit => VN_data_out(9136),
        VN2CN5_bit => VN_data_out(9137),
        VN2CN0_sign => VN_sign_out(9132),
        VN2CN1_sign => VN_sign_out(9133),
        VN2CN2_sign => VN_sign_out(9134),
        VN2CN3_sign => VN_sign_out(9135),
        VN2CN4_sign => VN_sign_out(9136),
        VN2CN5_sign => VN_sign_out(9137),
        codeword => codeword(1522),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1523 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9143 downto 9138),
        Din0 => VN1523_in0,
        Din1 => VN1523_in1,
        Din2 => VN1523_in2,
        Din3 => VN1523_in3,
        Din4 => VN1523_in4,
        Din5 => VN1523_in5,
        VN2CN0_bit => VN_data_out(9138),
        VN2CN1_bit => VN_data_out(9139),
        VN2CN2_bit => VN_data_out(9140),
        VN2CN3_bit => VN_data_out(9141),
        VN2CN4_bit => VN_data_out(9142),
        VN2CN5_bit => VN_data_out(9143),
        VN2CN0_sign => VN_sign_out(9138),
        VN2CN1_sign => VN_sign_out(9139),
        VN2CN2_sign => VN_sign_out(9140),
        VN2CN3_sign => VN_sign_out(9141),
        VN2CN4_sign => VN_sign_out(9142),
        VN2CN5_sign => VN_sign_out(9143),
        codeword => codeword(1523),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1524 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9149 downto 9144),
        Din0 => VN1524_in0,
        Din1 => VN1524_in1,
        Din2 => VN1524_in2,
        Din3 => VN1524_in3,
        Din4 => VN1524_in4,
        Din5 => VN1524_in5,
        VN2CN0_bit => VN_data_out(9144),
        VN2CN1_bit => VN_data_out(9145),
        VN2CN2_bit => VN_data_out(9146),
        VN2CN3_bit => VN_data_out(9147),
        VN2CN4_bit => VN_data_out(9148),
        VN2CN5_bit => VN_data_out(9149),
        VN2CN0_sign => VN_sign_out(9144),
        VN2CN1_sign => VN_sign_out(9145),
        VN2CN2_sign => VN_sign_out(9146),
        VN2CN3_sign => VN_sign_out(9147),
        VN2CN4_sign => VN_sign_out(9148),
        VN2CN5_sign => VN_sign_out(9149),
        codeword => codeword(1524),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1525 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9155 downto 9150),
        Din0 => VN1525_in0,
        Din1 => VN1525_in1,
        Din2 => VN1525_in2,
        Din3 => VN1525_in3,
        Din4 => VN1525_in4,
        Din5 => VN1525_in5,
        VN2CN0_bit => VN_data_out(9150),
        VN2CN1_bit => VN_data_out(9151),
        VN2CN2_bit => VN_data_out(9152),
        VN2CN3_bit => VN_data_out(9153),
        VN2CN4_bit => VN_data_out(9154),
        VN2CN5_bit => VN_data_out(9155),
        VN2CN0_sign => VN_sign_out(9150),
        VN2CN1_sign => VN_sign_out(9151),
        VN2CN2_sign => VN_sign_out(9152),
        VN2CN3_sign => VN_sign_out(9153),
        VN2CN4_sign => VN_sign_out(9154),
        VN2CN5_sign => VN_sign_out(9155),
        codeword => codeword(1525),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1526 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9161 downto 9156),
        Din0 => VN1526_in0,
        Din1 => VN1526_in1,
        Din2 => VN1526_in2,
        Din3 => VN1526_in3,
        Din4 => VN1526_in4,
        Din5 => VN1526_in5,
        VN2CN0_bit => VN_data_out(9156),
        VN2CN1_bit => VN_data_out(9157),
        VN2CN2_bit => VN_data_out(9158),
        VN2CN3_bit => VN_data_out(9159),
        VN2CN4_bit => VN_data_out(9160),
        VN2CN5_bit => VN_data_out(9161),
        VN2CN0_sign => VN_sign_out(9156),
        VN2CN1_sign => VN_sign_out(9157),
        VN2CN2_sign => VN_sign_out(9158),
        VN2CN3_sign => VN_sign_out(9159),
        VN2CN4_sign => VN_sign_out(9160),
        VN2CN5_sign => VN_sign_out(9161),
        codeword => codeword(1526),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1527 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9167 downto 9162),
        Din0 => VN1527_in0,
        Din1 => VN1527_in1,
        Din2 => VN1527_in2,
        Din3 => VN1527_in3,
        Din4 => VN1527_in4,
        Din5 => VN1527_in5,
        VN2CN0_bit => VN_data_out(9162),
        VN2CN1_bit => VN_data_out(9163),
        VN2CN2_bit => VN_data_out(9164),
        VN2CN3_bit => VN_data_out(9165),
        VN2CN4_bit => VN_data_out(9166),
        VN2CN5_bit => VN_data_out(9167),
        VN2CN0_sign => VN_sign_out(9162),
        VN2CN1_sign => VN_sign_out(9163),
        VN2CN2_sign => VN_sign_out(9164),
        VN2CN3_sign => VN_sign_out(9165),
        VN2CN4_sign => VN_sign_out(9166),
        VN2CN5_sign => VN_sign_out(9167),
        codeword => codeword(1527),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1528 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9173 downto 9168),
        Din0 => VN1528_in0,
        Din1 => VN1528_in1,
        Din2 => VN1528_in2,
        Din3 => VN1528_in3,
        Din4 => VN1528_in4,
        Din5 => VN1528_in5,
        VN2CN0_bit => VN_data_out(9168),
        VN2CN1_bit => VN_data_out(9169),
        VN2CN2_bit => VN_data_out(9170),
        VN2CN3_bit => VN_data_out(9171),
        VN2CN4_bit => VN_data_out(9172),
        VN2CN5_bit => VN_data_out(9173),
        VN2CN0_sign => VN_sign_out(9168),
        VN2CN1_sign => VN_sign_out(9169),
        VN2CN2_sign => VN_sign_out(9170),
        VN2CN3_sign => VN_sign_out(9171),
        VN2CN4_sign => VN_sign_out(9172),
        VN2CN5_sign => VN_sign_out(9173),
        codeword => codeword(1528),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1529 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9179 downto 9174),
        Din0 => VN1529_in0,
        Din1 => VN1529_in1,
        Din2 => VN1529_in2,
        Din3 => VN1529_in3,
        Din4 => VN1529_in4,
        Din5 => VN1529_in5,
        VN2CN0_bit => VN_data_out(9174),
        VN2CN1_bit => VN_data_out(9175),
        VN2CN2_bit => VN_data_out(9176),
        VN2CN3_bit => VN_data_out(9177),
        VN2CN4_bit => VN_data_out(9178),
        VN2CN5_bit => VN_data_out(9179),
        VN2CN0_sign => VN_sign_out(9174),
        VN2CN1_sign => VN_sign_out(9175),
        VN2CN2_sign => VN_sign_out(9176),
        VN2CN3_sign => VN_sign_out(9177),
        VN2CN4_sign => VN_sign_out(9178),
        VN2CN5_sign => VN_sign_out(9179),
        codeword => codeword(1529),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1530 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9185 downto 9180),
        Din0 => VN1530_in0,
        Din1 => VN1530_in1,
        Din2 => VN1530_in2,
        Din3 => VN1530_in3,
        Din4 => VN1530_in4,
        Din5 => VN1530_in5,
        VN2CN0_bit => VN_data_out(9180),
        VN2CN1_bit => VN_data_out(9181),
        VN2CN2_bit => VN_data_out(9182),
        VN2CN3_bit => VN_data_out(9183),
        VN2CN4_bit => VN_data_out(9184),
        VN2CN5_bit => VN_data_out(9185),
        VN2CN0_sign => VN_sign_out(9180),
        VN2CN1_sign => VN_sign_out(9181),
        VN2CN2_sign => VN_sign_out(9182),
        VN2CN3_sign => VN_sign_out(9183),
        VN2CN4_sign => VN_sign_out(9184),
        VN2CN5_sign => VN_sign_out(9185),
        codeword => codeword(1530),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1531 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9191 downto 9186),
        Din0 => VN1531_in0,
        Din1 => VN1531_in1,
        Din2 => VN1531_in2,
        Din3 => VN1531_in3,
        Din4 => VN1531_in4,
        Din5 => VN1531_in5,
        VN2CN0_bit => VN_data_out(9186),
        VN2CN1_bit => VN_data_out(9187),
        VN2CN2_bit => VN_data_out(9188),
        VN2CN3_bit => VN_data_out(9189),
        VN2CN4_bit => VN_data_out(9190),
        VN2CN5_bit => VN_data_out(9191),
        VN2CN0_sign => VN_sign_out(9186),
        VN2CN1_sign => VN_sign_out(9187),
        VN2CN2_sign => VN_sign_out(9188),
        VN2CN3_sign => VN_sign_out(9189),
        VN2CN4_sign => VN_sign_out(9190),
        VN2CN5_sign => VN_sign_out(9191),
        codeword => codeword(1531),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1532 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9197 downto 9192),
        Din0 => VN1532_in0,
        Din1 => VN1532_in1,
        Din2 => VN1532_in2,
        Din3 => VN1532_in3,
        Din4 => VN1532_in4,
        Din5 => VN1532_in5,
        VN2CN0_bit => VN_data_out(9192),
        VN2CN1_bit => VN_data_out(9193),
        VN2CN2_bit => VN_data_out(9194),
        VN2CN3_bit => VN_data_out(9195),
        VN2CN4_bit => VN_data_out(9196),
        VN2CN5_bit => VN_data_out(9197),
        VN2CN0_sign => VN_sign_out(9192),
        VN2CN1_sign => VN_sign_out(9193),
        VN2CN2_sign => VN_sign_out(9194),
        VN2CN3_sign => VN_sign_out(9195),
        VN2CN4_sign => VN_sign_out(9196),
        VN2CN5_sign => VN_sign_out(9197),
        codeword => codeword(1532),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1533 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9203 downto 9198),
        Din0 => VN1533_in0,
        Din1 => VN1533_in1,
        Din2 => VN1533_in2,
        Din3 => VN1533_in3,
        Din4 => VN1533_in4,
        Din5 => VN1533_in5,
        VN2CN0_bit => VN_data_out(9198),
        VN2CN1_bit => VN_data_out(9199),
        VN2CN2_bit => VN_data_out(9200),
        VN2CN3_bit => VN_data_out(9201),
        VN2CN4_bit => VN_data_out(9202),
        VN2CN5_bit => VN_data_out(9203),
        VN2CN0_sign => VN_sign_out(9198),
        VN2CN1_sign => VN_sign_out(9199),
        VN2CN2_sign => VN_sign_out(9200),
        VN2CN3_sign => VN_sign_out(9201),
        VN2CN4_sign => VN_sign_out(9202),
        VN2CN5_sign => VN_sign_out(9203),
        codeword => codeword(1533),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1534 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9209 downto 9204),
        Din0 => VN1534_in0,
        Din1 => VN1534_in1,
        Din2 => VN1534_in2,
        Din3 => VN1534_in3,
        Din4 => VN1534_in4,
        Din5 => VN1534_in5,
        VN2CN0_bit => VN_data_out(9204),
        VN2CN1_bit => VN_data_out(9205),
        VN2CN2_bit => VN_data_out(9206),
        VN2CN3_bit => VN_data_out(9207),
        VN2CN4_bit => VN_data_out(9208),
        VN2CN5_bit => VN_data_out(9209),
        VN2CN0_sign => VN_sign_out(9204),
        VN2CN1_sign => VN_sign_out(9205),
        VN2CN2_sign => VN_sign_out(9206),
        VN2CN3_sign => VN_sign_out(9207),
        VN2CN4_sign => VN_sign_out(9208),
        VN2CN5_sign => VN_sign_out(9209),
        codeword => codeword(1534),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1535 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9215 downto 9210),
        Din0 => VN1535_in0,
        Din1 => VN1535_in1,
        Din2 => VN1535_in2,
        Din3 => VN1535_in3,
        Din4 => VN1535_in4,
        Din5 => VN1535_in5,
        VN2CN0_bit => VN_data_out(9210),
        VN2CN1_bit => VN_data_out(9211),
        VN2CN2_bit => VN_data_out(9212),
        VN2CN3_bit => VN_data_out(9213),
        VN2CN4_bit => VN_data_out(9214),
        VN2CN5_bit => VN_data_out(9215),
        VN2CN0_sign => VN_sign_out(9210),
        VN2CN1_sign => VN_sign_out(9211),
        VN2CN2_sign => VN_sign_out(9212),
        VN2CN3_sign => VN_sign_out(9213),
        VN2CN4_sign => VN_sign_out(9214),
        VN2CN5_sign => VN_sign_out(9215),
        codeword => codeword(1535),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1536 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9221 downto 9216),
        Din0 => VN1536_in0,
        Din1 => VN1536_in1,
        Din2 => VN1536_in2,
        Din3 => VN1536_in3,
        Din4 => VN1536_in4,
        Din5 => VN1536_in5,
        VN2CN0_bit => VN_data_out(9216),
        VN2CN1_bit => VN_data_out(9217),
        VN2CN2_bit => VN_data_out(9218),
        VN2CN3_bit => VN_data_out(9219),
        VN2CN4_bit => VN_data_out(9220),
        VN2CN5_bit => VN_data_out(9221),
        VN2CN0_sign => VN_sign_out(9216),
        VN2CN1_sign => VN_sign_out(9217),
        VN2CN2_sign => VN_sign_out(9218),
        VN2CN3_sign => VN_sign_out(9219),
        VN2CN4_sign => VN_sign_out(9220),
        VN2CN5_sign => VN_sign_out(9221),
        codeword => codeword(1536),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1537 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9227 downto 9222),
        Din0 => VN1537_in0,
        Din1 => VN1537_in1,
        Din2 => VN1537_in2,
        Din3 => VN1537_in3,
        Din4 => VN1537_in4,
        Din5 => VN1537_in5,
        VN2CN0_bit => VN_data_out(9222),
        VN2CN1_bit => VN_data_out(9223),
        VN2CN2_bit => VN_data_out(9224),
        VN2CN3_bit => VN_data_out(9225),
        VN2CN4_bit => VN_data_out(9226),
        VN2CN5_bit => VN_data_out(9227),
        VN2CN0_sign => VN_sign_out(9222),
        VN2CN1_sign => VN_sign_out(9223),
        VN2CN2_sign => VN_sign_out(9224),
        VN2CN3_sign => VN_sign_out(9225),
        VN2CN4_sign => VN_sign_out(9226),
        VN2CN5_sign => VN_sign_out(9227),
        codeword => codeword(1537),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1538 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9233 downto 9228),
        Din0 => VN1538_in0,
        Din1 => VN1538_in1,
        Din2 => VN1538_in2,
        Din3 => VN1538_in3,
        Din4 => VN1538_in4,
        Din5 => VN1538_in5,
        VN2CN0_bit => VN_data_out(9228),
        VN2CN1_bit => VN_data_out(9229),
        VN2CN2_bit => VN_data_out(9230),
        VN2CN3_bit => VN_data_out(9231),
        VN2CN4_bit => VN_data_out(9232),
        VN2CN5_bit => VN_data_out(9233),
        VN2CN0_sign => VN_sign_out(9228),
        VN2CN1_sign => VN_sign_out(9229),
        VN2CN2_sign => VN_sign_out(9230),
        VN2CN3_sign => VN_sign_out(9231),
        VN2CN4_sign => VN_sign_out(9232),
        VN2CN5_sign => VN_sign_out(9233),
        codeword => codeword(1538),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1539 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9239 downto 9234),
        Din0 => VN1539_in0,
        Din1 => VN1539_in1,
        Din2 => VN1539_in2,
        Din3 => VN1539_in3,
        Din4 => VN1539_in4,
        Din5 => VN1539_in5,
        VN2CN0_bit => VN_data_out(9234),
        VN2CN1_bit => VN_data_out(9235),
        VN2CN2_bit => VN_data_out(9236),
        VN2CN3_bit => VN_data_out(9237),
        VN2CN4_bit => VN_data_out(9238),
        VN2CN5_bit => VN_data_out(9239),
        VN2CN0_sign => VN_sign_out(9234),
        VN2CN1_sign => VN_sign_out(9235),
        VN2CN2_sign => VN_sign_out(9236),
        VN2CN3_sign => VN_sign_out(9237),
        VN2CN4_sign => VN_sign_out(9238),
        VN2CN5_sign => VN_sign_out(9239),
        codeword => codeword(1539),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1540 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9245 downto 9240),
        Din0 => VN1540_in0,
        Din1 => VN1540_in1,
        Din2 => VN1540_in2,
        Din3 => VN1540_in3,
        Din4 => VN1540_in4,
        Din5 => VN1540_in5,
        VN2CN0_bit => VN_data_out(9240),
        VN2CN1_bit => VN_data_out(9241),
        VN2CN2_bit => VN_data_out(9242),
        VN2CN3_bit => VN_data_out(9243),
        VN2CN4_bit => VN_data_out(9244),
        VN2CN5_bit => VN_data_out(9245),
        VN2CN0_sign => VN_sign_out(9240),
        VN2CN1_sign => VN_sign_out(9241),
        VN2CN2_sign => VN_sign_out(9242),
        VN2CN3_sign => VN_sign_out(9243),
        VN2CN4_sign => VN_sign_out(9244),
        VN2CN5_sign => VN_sign_out(9245),
        codeword => codeword(1540),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1541 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9251 downto 9246),
        Din0 => VN1541_in0,
        Din1 => VN1541_in1,
        Din2 => VN1541_in2,
        Din3 => VN1541_in3,
        Din4 => VN1541_in4,
        Din5 => VN1541_in5,
        VN2CN0_bit => VN_data_out(9246),
        VN2CN1_bit => VN_data_out(9247),
        VN2CN2_bit => VN_data_out(9248),
        VN2CN3_bit => VN_data_out(9249),
        VN2CN4_bit => VN_data_out(9250),
        VN2CN5_bit => VN_data_out(9251),
        VN2CN0_sign => VN_sign_out(9246),
        VN2CN1_sign => VN_sign_out(9247),
        VN2CN2_sign => VN_sign_out(9248),
        VN2CN3_sign => VN_sign_out(9249),
        VN2CN4_sign => VN_sign_out(9250),
        VN2CN5_sign => VN_sign_out(9251),
        codeword => codeword(1541),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1542 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9257 downto 9252),
        Din0 => VN1542_in0,
        Din1 => VN1542_in1,
        Din2 => VN1542_in2,
        Din3 => VN1542_in3,
        Din4 => VN1542_in4,
        Din5 => VN1542_in5,
        VN2CN0_bit => VN_data_out(9252),
        VN2CN1_bit => VN_data_out(9253),
        VN2CN2_bit => VN_data_out(9254),
        VN2CN3_bit => VN_data_out(9255),
        VN2CN4_bit => VN_data_out(9256),
        VN2CN5_bit => VN_data_out(9257),
        VN2CN0_sign => VN_sign_out(9252),
        VN2CN1_sign => VN_sign_out(9253),
        VN2CN2_sign => VN_sign_out(9254),
        VN2CN3_sign => VN_sign_out(9255),
        VN2CN4_sign => VN_sign_out(9256),
        VN2CN5_sign => VN_sign_out(9257),
        codeword => codeword(1542),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1543 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9263 downto 9258),
        Din0 => VN1543_in0,
        Din1 => VN1543_in1,
        Din2 => VN1543_in2,
        Din3 => VN1543_in3,
        Din4 => VN1543_in4,
        Din5 => VN1543_in5,
        VN2CN0_bit => VN_data_out(9258),
        VN2CN1_bit => VN_data_out(9259),
        VN2CN2_bit => VN_data_out(9260),
        VN2CN3_bit => VN_data_out(9261),
        VN2CN4_bit => VN_data_out(9262),
        VN2CN5_bit => VN_data_out(9263),
        VN2CN0_sign => VN_sign_out(9258),
        VN2CN1_sign => VN_sign_out(9259),
        VN2CN2_sign => VN_sign_out(9260),
        VN2CN3_sign => VN_sign_out(9261),
        VN2CN4_sign => VN_sign_out(9262),
        VN2CN5_sign => VN_sign_out(9263),
        codeword => codeword(1543),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1544 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9269 downto 9264),
        Din0 => VN1544_in0,
        Din1 => VN1544_in1,
        Din2 => VN1544_in2,
        Din3 => VN1544_in3,
        Din4 => VN1544_in4,
        Din5 => VN1544_in5,
        VN2CN0_bit => VN_data_out(9264),
        VN2CN1_bit => VN_data_out(9265),
        VN2CN2_bit => VN_data_out(9266),
        VN2CN3_bit => VN_data_out(9267),
        VN2CN4_bit => VN_data_out(9268),
        VN2CN5_bit => VN_data_out(9269),
        VN2CN0_sign => VN_sign_out(9264),
        VN2CN1_sign => VN_sign_out(9265),
        VN2CN2_sign => VN_sign_out(9266),
        VN2CN3_sign => VN_sign_out(9267),
        VN2CN4_sign => VN_sign_out(9268),
        VN2CN5_sign => VN_sign_out(9269),
        codeword => codeword(1544),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1545 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9275 downto 9270),
        Din0 => VN1545_in0,
        Din1 => VN1545_in1,
        Din2 => VN1545_in2,
        Din3 => VN1545_in3,
        Din4 => VN1545_in4,
        Din5 => VN1545_in5,
        VN2CN0_bit => VN_data_out(9270),
        VN2CN1_bit => VN_data_out(9271),
        VN2CN2_bit => VN_data_out(9272),
        VN2CN3_bit => VN_data_out(9273),
        VN2CN4_bit => VN_data_out(9274),
        VN2CN5_bit => VN_data_out(9275),
        VN2CN0_sign => VN_sign_out(9270),
        VN2CN1_sign => VN_sign_out(9271),
        VN2CN2_sign => VN_sign_out(9272),
        VN2CN3_sign => VN_sign_out(9273),
        VN2CN4_sign => VN_sign_out(9274),
        VN2CN5_sign => VN_sign_out(9275),
        codeword => codeword(1545),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1546 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9281 downto 9276),
        Din0 => VN1546_in0,
        Din1 => VN1546_in1,
        Din2 => VN1546_in2,
        Din3 => VN1546_in3,
        Din4 => VN1546_in4,
        Din5 => VN1546_in5,
        VN2CN0_bit => VN_data_out(9276),
        VN2CN1_bit => VN_data_out(9277),
        VN2CN2_bit => VN_data_out(9278),
        VN2CN3_bit => VN_data_out(9279),
        VN2CN4_bit => VN_data_out(9280),
        VN2CN5_bit => VN_data_out(9281),
        VN2CN0_sign => VN_sign_out(9276),
        VN2CN1_sign => VN_sign_out(9277),
        VN2CN2_sign => VN_sign_out(9278),
        VN2CN3_sign => VN_sign_out(9279),
        VN2CN4_sign => VN_sign_out(9280),
        VN2CN5_sign => VN_sign_out(9281),
        codeword => codeword(1546),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1547 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9287 downto 9282),
        Din0 => VN1547_in0,
        Din1 => VN1547_in1,
        Din2 => VN1547_in2,
        Din3 => VN1547_in3,
        Din4 => VN1547_in4,
        Din5 => VN1547_in5,
        VN2CN0_bit => VN_data_out(9282),
        VN2CN1_bit => VN_data_out(9283),
        VN2CN2_bit => VN_data_out(9284),
        VN2CN3_bit => VN_data_out(9285),
        VN2CN4_bit => VN_data_out(9286),
        VN2CN5_bit => VN_data_out(9287),
        VN2CN0_sign => VN_sign_out(9282),
        VN2CN1_sign => VN_sign_out(9283),
        VN2CN2_sign => VN_sign_out(9284),
        VN2CN3_sign => VN_sign_out(9285),
        VN2CN4_sign => VN_sign_out(9286),
        VN2CN5_sign => VN_sign_out(9287),
        codeword => codeword(1547),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1548 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9293 downto 9288),
        Din0 => VN1548_in0,
        Din1 => VN1548_in1,
        Din2 => VN1548_in2,
        Din3 => VN1548_in3,
        Din4 => VN1548_in4,
        Din5 => VN1548_in5,
        VN2CN0_bit => VN_data_out(9288),
        VN2CN1_bit => VN_data_out(9289),
        VN2CN2_bit => VN_data_out(9290),
        VN2CN3_bit => VN_data_out(9291),
        VN2CN4_bit => VN_data_out(9292),
        VN2CN5_bit => VN_data_out(9293),
        VN2CN0_sign => VN_sign_out(9288),
        VN2CN1_sign => VN_sign_out(9289),
        VN2CN2_sign => VN_sign_out(9290),
        VN2CN3_sign => VN_sign_out(9291),
        VN2CN4_sign => VN_sign_out(9292),
        VN2CN5_sign => VN_sign_out(9293),
        codeword => codeword(1548),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1549 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9299 downto 9294),
        Din0 => VN1549_in0,
        Din1 => VN1549_in1,
        Din2 => VN1549_in2,
        Din3 => VN1549_in3,
        Din4 => VN1549_in4,
        Din5 => VN1549_in5,
        VN2CN0_bit => VN_data_out(9294),
        VN2CN1_bit => VN_data_out(9295),
        VN2CN2_bit => VN_data_out(9296),
        VN2CN3_bit => VN_data_out(9297),
        VN2CN4_bit => VN_data_out(9298),
        VN2CN5_bit => VN_data_out(9299),
        VN2CN0_sign => VN_sign_out(9294),
        VN2CN1_sign => VN_sign_out(9295),
        VN2CN2_sign => VN_sign_out(9296),
        VN2CN3_sign => VN_sign_out(9297),
        VN2CN4_sign => VN_sign_out(9298),
        VN2CN5_sign => VN_sign_out(9299),
        codeword => codeword(1549),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1550 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9305 downto 9300),
        Din0 => VN1550_in0,
        Din1 => VN1550_in1,
        Din2 => VN1550_in2,
        Din3 => VN1550_in3,
        Din4 => VN1550_in4,
        Din5 => VN1550_in5,
        VN2CN0_bit => VN_data_out(9300),
        VN2CN1_bit => VN_data_out(9301),
        VN2CN2_bit => VN_data_out(9302),
        VN2CN3_bit => VN_data_out(9303),
        VN2CN4_bit => VN_data_out(9304),
        VN2CN5_bit => VN_data_out(9305),
        VN2CN0_sign => VN_sign_out(9300),
        VN2CN1_sign => VN_sign_out(9301),
        VN2CN2_sign => VN_sign_out(9302),
        VN2CN3_sign => VN_sign_out(9303),
        VN2CN4_sign => VN_sign_out(9304),
        VN2CN5_sign => VN_sign_out(9305),
        codeword => codeword(1550),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1551 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9311 downto 9306),
        Din0 => VN1551_in0,
        Din1 => VN1551_in1,
        Din2 => VN1551_in2,
        Din3 => VN1551_in3,
        Din4 => VN1551_in4,
        Din5 => VN1551_in5,
        VN2CN0_bit => VN_data_out(9306),
        VN2CN1_bit => VN_data_out(9307),
        VN2CN2_bit => VN_data_out(9308),
        VN2CN3_bit => VN_data_out(9309),
        VN2CN4_bit => VN_data_out(9310),
        VN2CN5_bit => VN_data_out(9311),
        VN2CN0_sign => VN_sign_out(9306),
        VN2CN1_sign => VN_sign_out(9307),
        VN2CN2_sign => VN_sign_out(9308),
        VN2CN3_sign => VN_sign_out(9309),
        VN2CN4_sign => VN_sign_out(9310),
        VN2CN5_sign => VN_sign_out(9311),
        codeword => codeword(1551),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1552 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9317 downto 9312),
        Din0 => VN1552_in0,
        Din1 => VN1552_in1,
        Din2 => VN1552_in2,
        Din3 => VN1552_in3,
        Din4 => VN1552_in4,
        Din5 => VN1552_in5,
        VN2CN0_bit => VN_data_out(9312),
        VN2CN1_bit => VN_data_out(9313),
        VN2CN2_bit => VN_data_out(9314),
        VN2CN3_bit => VN_data_out(9315),
        VN2CN4_bit => VN_data_out(9316),
        VN2CN5_bit => VN_data_out(9317),
        VN2CN0_sign => VN_sign_out(9312),
        VN2CN1_sign => VN_sign_out(9313),
        VN2CN2_sign => VN_sign_out(9314),
        VN2CN3_sign => VN_sign_out(9315),
        VN2CN4_sign => VN_sign_out(9316),
        VN2CN5_sign => VN_sign_out(9317),
        codeword => codeword(1552),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1553 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9323 downto 9318),
        Din0 => VN1553_in0,
        Din1 => VN1553_in1,
        Din2 => VN1553_in2,
        Din3 => VN1553_in3,
        Din4 => VN1553_in4,
        Din5 => VN1553_in5,
        VN2CN0_bit => VN_data_out(9318),
        VN2CN1_bit => VN_data_out(9319),
        VN2CN2_bit => VN_data_out(9320),
        VN2CN3_bit => VN_data_out(9321),
        VN2CN4_bit => VN_data_out(9322),
        VN2CN5_bit => VN_data_out(9323),
        VN2CN0_sign => VN_sign_out(9318),
        VN2CN1_sign => VN_sign_out(9319),
        VN2CN2_sign => VN_sign_out(9320),
        VN2CN3_sign => VN_sign_out(9321),
        VN2CN4_sign => VN_sign_out(9322),
        VN2CN5_sign => VN_sign_out(9323),
        codeword => codeword(1553),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1554 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9329 downto 9324),
        Din0 => VN1554_in0,
        Din1 => VN1554_in1,
        Din2 => VN1554_in2,
        Din3 => VN1554_in3,
        Din4 => VN1554_in4,
        Din5 => VN1554_in5,
        VN2CN0_bit => VN_data_out(9324),
        VN2CN1_bit => VN_data_out(9325),
        VN2CN2_bit => VN_data_out(9326),
        VN2CN3_bit => VN_data_out(9327),
        VN2CN4_bit => VN_data_out(9328),
        VN2CN5_bit => VN_data_out(9329),
        VN2CN0_sign => VN_sign_out(9324),
        VN2CN1_sign => VN_sign_out(9325),
        VN2CN2_sign => VN_sign_out(9326),
        VN2CN3_sign => VN_sign_out(9327),
        VN2CN4_sign => VN_sign_out(9328),
        VN2CN5_sign => VN_sign_out(9329),
        codeword => codeword(1554),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1555 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9335 downto 9330),
        Din0 => VN1555_in0,
        Din1 => VN1555_in1,
        Din2 => VN1555_in2,
        Din3 => VN1555_in3,
        Din4 => VN1555_in4,
        Din5 => VN1555_in5,
        VN2CN0_bit => VN_data_out(9330),
        VN2CN1_bit => VN_data_out(9331),
        VN2CN2_bit => VN_data_out(9332),
        VN2CN3_bit => VN_data_out(9333),
        VN2CN4_bit => VN_data_out(9334),
        VN2CN5_bit => VN_data_out(9335),
        VN2CN0_sign => VN_sign_out(9330),
        VN2CN1_sign => VN_sign_out(9331),
        VN2CN2_sign => VN_sign_out(9332),
        VN2CN3_sign => VN_sign_out(9333),
        VN2CN4_sign => VN_sign_out(9334),
        VN2CN5_sign => VN_sign_out(9335),
        codeword => codeword(1555),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1556 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9341 downto 9336),
        Din0 => VN1556_in0,
        Din1 => VN1556_in1,
        Din2 => VN1556_in2,
        Din3 => VN1556_in3,
        Din4 => VN1556_in4,
        Din5 => VN1556_in5,
        VN2CN0_bit => VN_data_out(9336),
        VN2CN1_bit => VN_data_out(9337),
        VN2CN2_bit => VN_data_out(9338),
        VN2CN3_bit => VN_data_out(9339),
        VN2CN4_bit => VN_data_out(9340),
        VN2CN5_bit => VN_data_out(9341),
        VN2CN0_sign => VN_sign_out(9336),
        VN2CN1_sign => VN_sign_out(9337),
        VN2CN2_sign => VN_sign_out(9338),
        VN2CN3_sign => VN_sign_out(9339),
        VN2CN4_sign => VN_sign_out(9340),
        VN2CN5_sign => VN_sign_out(9341),
        codeword => codeword(1556),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1557 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9347 downto 9342),
        Din0 => VN1557_in0,
        Din1 => VN1557_in1,
        Din2 => VN1557_in2,
        Din3 => VN1557_in3,
        Din4 => VN1557_in4,
        Din5 => VN1557_in5,
        VN2CN0_bit => VN_data_out(9342),
        VN2CN1_bit => VN_data_out(9343),
        VN2CN2_bit => VN_data_out(9344),
        VN2CN3_bit => VN_data_out(9345),
        VN2CN4_bit => VN_data_out(9346),
        VN2CN5_bit => VN_data_out(9347),
        VN2CN0_sign => VN_sign_out(9342),
        VN2CN1_sign => VN_sign_out(9343),
        VN2CN2_sign => VN_sign_out(9344),
        VN2CN3_sign => VN_sign_out(9345),
        VN2CN4_sign => VN_sign_out(9346),
        VN2CN5_sign => VN_sign_out(9347),
        codeword => codeword(1557),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1558 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9353 downto 9348),
        Din0 => VN1558_in0,
        Din1 => VN1558_in1,
        Din2 => VN1558_in2,
        Din3 => VN1558_in3,
        Din4 => VN1558_in4,
        Din5 => VN1558_in5,
        VN2CN0_bit => VN_data_out(9348),
        VN2CN1_bit => VN_data_out(9349),
        VN2CN2_bit => VN_data_out(9350),
        VN2CN3_bit => VN_data_out(9351),
        VN2CN4_bit => VN_data_out(9352),
        VN2CN5_bit => VN_data_out(9353),
        VN2CN0_sign => VN_sign_out(9348),
        VN2CN1_sign => VN_sign_out(9349),
        VN2CN2_sign => VN_sign_out(9350),
        VN2CN3_sign => VN_sign_out(9351),
        VN2CN4_sign => VN_sign_out(9352),
        VN2CN5_sign => VN_sign_out(9353),
        codeword => codeword(1558),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1559 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9359 downto 9354),
        Din0 => VN1559_in0,
        Din1 => VN1559_in1,
        Din2 => VN1559_in2,
        Din3 => VN1559_in3,
        Din4 => VN1559_in4,
        Din5 => VN1559_in5,
        VN2CN0_bit => VN_data_out(9354),
        VN2CN1_bit => VN_data_out(9355),
        VN2CN2_bit => VN_data_out(9356),
        VN2CN3_bit => VN_data_out(9357),
        VN2CN4_bit => VN_data_out(9358),
        VN2CN5_bit => VN_data_out(9359),
        VN2CN0_sign => VN_sign_out(9354),
        VN2CN1_sign => VN_sign_out(9355),
        VN2CN2_sign => VN_sign_out(9356),
        VN2CN3_sign => VN_sign_out(9357),
        VN2CN4_sign => VN_sign_out(9358),
        VN2CN5_sign => VN_sign_out(9359),
        codeword => codeword(1559),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1560 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9365 downto 9360),
        Din0 => VN1560_in0,
        Din1 => VN1560_in1,
        Din2 => VN1560_in2,
        Din3 => VN1560_in3,
        Din4 => VN1560_in4,
        Din5 => VN1560_in5,
        VN2CN0_bit => VN_data_out(9360),
        VN2CN1_bit => VN_data_out(9361),
        VN2CN2_bit => VN_data_out(9362),
        VN2CN3_bit => VN_data_out(9363),
        VN2CN4_bit => VN_data_out(9364),
        VN2CN5_bit => VN_data_out(9365),
        VN2CN0_sign => VN_sign_out(9360),
        VN2CN1_sign => VN_sign_out(9361),
        VN2CN2_sign => VN_sign_out(9362),
        VN2CN3_sign => VN_sign_out(9363),
        VN2CN4_sign => VN_sign_out(9364),
        VN2CN5_sign => VN_sign_out(9365),
        codeword => codeword(1560),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1561 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9371 downto 9366),
        Din0 => VN1561_in0,
        Din1 => VN1561_in1,
        Din2 => VN1561_in2,
        Din3 => VN1561_in3,
        Din4 => VN1561_in4,
        Din5 => VN1561_in5,
        VN2CN0_bit => VN_data_out(9366),
        VN2CN1_bit => VN_data_out(9367),
        VN2CN2_bit => VN_data_out(9368),
        VN2CN3_bit => VN_data_out(9369),
        VN2CN4_bit => VN_data_out(9370),
        VN2CN5_bit => VN_data_out(9371),
        VN2CN0_sign => VN_sign_out(9366),
        VN2CN1_sign => VN_sign_out(9367),
        VN2CN2_sign => VN_sign_out(9368),
        VN2CN3_sign => VN_sign_out(9369),
        VN2CN4_sign => VN_sign_out(9370),
        VN2CN5_sign => VN_sign_out(9371),
        codeword => codeword(1561),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1562 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9377 downto 9372),
        Din0 => VN1562_in0,
        Din1 => VN1562_in1,
        Din2 => VN1562_in2,
        Din3 => VN1562_in3,
        Din4 => VN1562_in4,
        Din5 => VN1562_in5,
        VN2CN0_bit => VN_data_out(9372),
        VN2CN1_bit => VN_data_out(9373),
        VN2CN2_bit => VN_data_out(9374),
        VN2CN3_bit => VN_data_out(9375),
        VN2CN4_bit => VN_data_out(9376),
        VN2CN5_bit => VN_data_out(9377),
        VN2CN0_sign => VN_sign_out(9372),
        VN2CN1_sign => VN_sign_out(9373),
        VN2CN2_sign => VN_sign_out(9374),
        VN2CN3_sign => VN_sign_out(9375),
        VN2CN4_sign => VN_sign_out(9376),
        VN2CN5_sign => VN_sign_out(9377),
        codeword => codeword(1562),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1563 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9383 downto 9378),
        Din0 => VN1563_in0,
        Din1 => VN1563_in1,
        Din2 => VN1563_in2,
        Din3 => VN1563_in3,
        Din4 => VN1563_in4,
        Din5 => VN1563_in5,
        VN2CN0_bit => VN_data_out(9378),
        VN2CN1_bit => VN_data_out(9379),
        VN2CN2_bit => VN_data_out(9380),
        VN2CN3_bit => VN_data_out(9381),
        VN2CN4_bit => VN_data_out(9382),
        VN2CN5_bit => VN_data_out(9383),
        VN2CN0_sign => VN_sign_out(9378),
        VN2CN1_sign => VN_sign_out(9379),
        VN2CN2_sign => VN_sign_out(9380),
        VN2CN3_sign => VN_sign_out(9381),
        VN2CN4_sign => VN_sign_out(9382),
        VN2CN5_sign => VN_sign_out(9383),
        codeword => codeword(1563),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1564 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9389 downto 9384),
        Din0 => VN1564_in0,
        Din1 => VN1564_in1,
        Din2 => VN1564_in2,
        Din3 => VN1564_in3,
        Din4 => VN1564_in4,
        Din5 => VN1564_in5,
        VN2CN0_bit => VN_data_out(9384),
        VN2CN1_bit => VN_data_out(9385),
        VN2CN2_bit => VN_data_out(9386),
        VN2CN3_bit => VN_data_out(9387),
        VN2CN4_bit => VN_data_out(9388),
        VN2CN5_bit => VN_data_out(9389),
        VN2CN0_sign => VN_sign_out(9384),
        VN2CN1_sign => VN_sign_out(9385),
        VN2CN2_sign => VN_sign_out(9386),
        VN2CN3_sign => VN_sign_out(9387),
        VN2CN4_sign => VN_sign_out(9388),
        VN2CN5_sign => VN_sign_out(9389),
        codeword => codeword(1564),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1565 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9395 downto 9390),
        Din0 => VN1565_in0,
        Din1 => VN1565_in1,
        Din2 => VN1565_in2,
        Din3 => VN1565_in3,
        Din4 => VN1565_in4,
        Din5 => VN1565_in5,
        VN2CN0_bit => VN_data_out(9390),
        VN2CN1_bit => VN_data_out(9391),
        VN2CN2_bit => VN_data_out(9392),
        VN2CN3_bit => VN_data_out(9393),
        VN2CN4_bit => VN_data_out(9394),
        VN2CN5_bit => VN_data_out(9395),
        VN2CN0_sign => VN_sign_out(9390),
        VN2CN1_sign => VN_sign_out(9391),
        VN2CN2_sign => VN_sign_out(9392),
        VN2CN3_sign => VN_sign_out(9393),
        VN2CN4_sign => VN_sign_out(9394),
        VN2CN5_sign => VN_sign_out(9395),
        codeword => codeword(1565),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1566 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9401 downto 9396),
        Din0 => VN1566_in0,
        Din1 => VN1566_in1,
        Din2 => VN1566_in2,
        Din3 => VN1566_in3,
        Din4 => VN1566_in4,
        Din5 => VN1566_in5,
        VN2CN0_bit => VN_data_out(9396),
        VN2CN1_bit => VN_data_out(9397),
        VN2CN2_bit => VN_data_out(9398),
        VN2CN3_bit => VN_data_out(9399),
        VN2CN4_bit => VN_data_out(9400),
        VN2CN5_bit => VN_data_out(9401),
        VN2CN0_sign => VN_sign_out(9396),
        VN2CN1_sign => VN_sign_out(9397),
        VN2CN2_sign => VN_sign_out(9398),
        VN2CN3_sign => VN_sign_out(9399),
        VN2CN4_sign => VN_sign_out(9400),
        VN2CN5_sign => VN_sign_out(9401),
        codeword => codeword(1566),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1567 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9407 downto 9402),
        Din0 => VN1567_in0,
        Din1 => VN1567_in1,
        Din2 => VN1567_in2,
        Din3 => VN1567_in3,
        Din4 => VN1567_in4,
        Din5 => VN1567_in5,
        VN2CN0_bit => VN_data_out(9402),
        VN2CN1_bit => VN_data_out(9403),
        VN2CN2_bit => VN_data_out(9404),
        VN2CN3_bit => VN_data_out(9405),
        VN2CN4_bit => VN_data_out(9406),
        VN2CN5_bit => VN_data_out(9407),
        VN2CN0_sign => VN_sign_out(9402),
        VN2CN1_sign => VN_sign_out(9403),
        VN2CN2_sign => VN_sign_out(9404),
        VN2CN3_sign => VN_sign_out(9405),
        VN2CN4_sign => VN_sign_out(9406),
        VN2CN5_sign => VN_sign_out(9407),
        codeword => codeword(1567),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1568 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9413 downto 9408),
        Din0 => VN1568_in0,
        Din1 => VN1568_in1,
        Din2 => VN1568_in2,
        Din3 => VN1568_in3,
        Din4 => VN1568_in4,
        Din5 => VN1568_in5,
        VN2CN0_bit => VN_data_out(9408),
        VN2CN1_bit => VN_data_out(9409),
        VN2CN2_bit => VN_data_out(9410),
        VN2CN3_bit => VN_data_out(9411),
        VN2CN4_bit => VN_data_out(9412),
        VN2CN5_bit => VN_data_out(9413),
        VN2CN0_sign => VN_sign_out(9408),
        VN2CN1_sign => VN_sign_out(9409),
        VN2CN2_sign => VN_sign_out(9410),
        VN2CN3_sign => VN_sign_out(9411),
        VN2CN4_sign => VN_sign_out(9412),
        VN2CN5_sign => VN_sign_out(9413),
        codeword => codeword(1568),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1569 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9419 downto 9414),
        Din0 => VN1569_in0,
        Din1 => VN1569_in1,
        Din2 => VN1569_in2,
        Din3 => VN1569_in3,
        Din4 => VN1569_in4,
        Din5 => VN1569_in5,
        VN2CN0_bit => VN_data_out(9414),
        VN2CN1_bit => VN_data_out(9415),
        VN2CN2_bit => VN_data_out(9416),
        VN2CN3_bit => VN_data_out(9417),
        VN2CN4_bit => VN_data_out(9418),
        VN2CN5_bit => VN_data_out(9419),
        VN2CN0_sign => VN_sign_out(9414),
        VN2CN1_sign => VN_sign_out(9415),
        VN2CN2_sign => VN_sign_out(9416),
        VN2CN3_sign => VN_sign_out(9417),
        VN2CN4_sign => VN_sign_out(9418),
        VN2CN5_sign => VN_sign_out(9419),
        codeword => codeword(1569),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1570 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9425 downto 9420),
        Din0 => VN1570_in0,
        Din1 => VN1570_in1,
        Din2 => VN1570_in2,
        Din3 => VN1570_in3,
        Din4 => VN1570_in4,
        Din5 => VN1570_in5,
        VN2CN0_bit => VN_data_out(9420),
        VN2CN1_bit => VN_data_out(9421),
        VN2CN2_bit => VN_data_out(9422),
        VN2CN3_bit => VN_data_out(9423),
        VN2CN4_bit => VN_data_out(9424),
        VN2CN5_bit => VN_data_out(9425),
        VN2CN0_sign => VN_sign_out(9420),
        VN2CN1_sign => VN_sign_out(9421),
        VN2CN2_sign => VN_sign_out(9422),
        VN2CN3_sign => VN_sign_out(9423),
        VN2CN4_sign => VN_sign_out(9424),
        VN2CN5_sign => VN_sign_out(9425),
        codeword => codeword(1570),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1571 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9431 downto 9426),
        Din0 => VN1571_in0,
        Din1 => VN1571_in1,
        Din2 => VN1571_in2,
        Din3 => VN1571_in3,
        Din4 => VN1571_in4,
        Din5 => VN1571_in5,
        VN2CN0_bit => VN_data_out(9426),
        VN2CN1_bit => VN_data_out(9427),
        VN2CN2_bit => VN_data_out(9428),
        VN2CN3_bit => VN_data_out(9429),
        VN2CN4_bit => VN_data_out(9430),
        VN2CN5_bit => VN_data_out(9431),
        VN2CN0_sign => VN_sign_out(9426),
        VN2CN1_sign => VN_sign_out(9427),
        VN2CN2_sign => VN_sign_out(9428),
        VN2CN3_sign => VN_sign_out(9429),
        VN2CN4_sign => VN_sign_out(9430),
        VN2CN5_sign => VN_sign_out(9431),
        codeword => codeword(1571),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1572 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9437 downto 9432),
        Din0 => VN1572_in0,
        Din1 => VN1572_in1,
        Din2 => VN1572_in2,
        Din3 => VN1572_in3,
        Din4 => VN1572_in4,
        Din5 => VN1572_in5,
        VN2CN0_bit => VN_data_out(9432),
        VN2CN1_bit => VN_data_out(9433),
        VN2CN2_bit => VN_data_out(9434),
        VN2CN3_bit => VN_data_out(9435),
        VN2CN4_bit => VN_data_out(9436),
        VN2CN5_bit => VN_data_out(9437),
        VN2CN0_sign => VN_sign_out(9432),
        VN2CN1_sign => VN_sign_out(9433),
        VN2CN2_sign => VN_sign_out(9434),
        VN2CN3_sign => VN_sign_out(9435),
        VN2CN4_sign => VN_sign_out(9436),
        VN2CN5_sign => VN_sign_out(9437),
        codeword => codeword(1572),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1573 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9443 downto 9438),
        Din0 => VN1573_in0,
        Din1 => VN1573_in1,
        Din2 => VN1573_in2,
        Din3 => VN1573_in3,
        Din4 => VN1573_in4,
        Din5 => VN1573_in5,
        VN2CN0_bit => VN_data_out(9438),
        VN2CN1_bit => VN_data_out(9439),
        VN2CN2_bit => VN_data_out(9440),
        VN2CN3_bit => VN_data_out(9441),
        VN2CN4_bit => VN_data_out(9442),
        VN2CN5_bit => VN_data_out(9443),
        VN2CN0_sign => VN_sign_out(9438),
        VN2CN1_sign => VN_sign_out(9439),
        VN2CN2_sign => VN_sign_out(9440),
        VN2CN3_sign => VN_sign_out(9441),
        VN2CN4_sign => VN_sign_out(9442),
        VN2CN5_sign => VN_sign_out(9443),
        codeword => codeword(1573),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1574 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9449 downto 9444),
        Din0 => VN1574_in0,
        Din1 => VN1574_in1,
        Din2 => VN1574_in2,
        Din3 => VN1574_in3,
        Din4 => VN1574_in4,
        Din5 => VN1574_in5,
        VN2CN0_bit => VN_data_out(9444),
        VN2CN1_bit => VN_data_out(9445),
        VN2CN2_bit => VN_data_out(9446),
        VN2CN3_bit => VN_data_out(9447),
        VN2CN4_bit => VN_data_out(9448),
        VN2CN5_bit => VN_data_out(9449),
        VN2CN0_sign => VN_sign_out(9444),
        VN2CN1_sign => VN_sign_out(9445),
        VN2CN2_sign => VN_sign_out(9446),
        VN2CN3_sign => VN_sign_out(9447),
        VN2CN4_sign => VN_sign_out(9448),
        VN2CN5_sign => VN_sign_out(9449),
        codeword => codeword(1574),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1575 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9455 downto 9450),
        Din0 => VN1575_in0,
        Din1 => VN1575_in1,
        Din2 => VN1575_in2,
        Din3 => VN1575_in3,
        Din4 => VN1575_in4,
        Din5 => VN1575_in5,
        VN2CN0_bit => VN_data_out(9450),
        VN2CN1_bit => VN_data_out(9451),
        VN2CN2_bit => VN_data_out(9452),
        VN2CN3_bit => VN_data_out(9453),
        VN2CN4_bit => VN_data_out(9454),
        VN2CN5_bit => VN_data_out(9455),
        VN2CN0_sign => VN_sign_out(9450),
        VN2CN1_sign => VN_sign_out(9451),
        VN2CN2_sign => VN_sign_out(9452),
        VN2CN3_sign => VN_sign_out(9453),
        VN2CN4_sign => VN_sign_out(9454),
        VN2CN5_sign => VN_sign_out(9455),
        codeword => codeword(1575),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1576 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9461 downto 9456),
        Din0 => VN1576_in0,
        Din1 => VN1576_in1,
        Din2 => VN1576_in2,
        Din3 => VN1576_in3,
        Din4 => VN1576_in4,
        Din5 => VN1576_in5,
        VN2CN0_bit => VN_data_out(9456),
        VN2CN1_bit => VN_data_out(9457),
        VN2CN2_bit => VN_data_out(9458),
        VN2CN3_bit => VN_data_out(9459),
        VN2CN4_bit => VN_data_out(9460),
        VN2CN5_bit => VN_data_out(9461),
        VN2CN0_sign => VN_sign_out(9456),
        VN2CN1_sign => VN_sign_out(9457),
        VN2CN2_sign => VN_sign_out(9458),
        VN2CN3_sign => VN_sign_out(9459),
        VN2CN4_sign => VN_sign_out(9460),
        VN2CN5_sign => VN_sign_out(9461),
        codeword => codeword(1576),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1577 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9467 downto 9462),
        Din0 => VN1577_in0,
        Din1 => VN1577_in1,
        Din2 => VN1577_in2,
        Din3 => VN1577_in3,
        Din4 => VN1577_in4,
        Din5 => VN1577_in5,
        VN2CN0_bit => VN_data_out(9462),
        VN2CN1_bit => VN_data_out(9463),
        VN2CN2_bit => VN_data_out(9464),
        VN2CN3_bit => VN_data_out(9465),
        VN2CN4_bit => VN_data_out(9466),
        VN2CN5_bit => VN_data_out(9467),
        VN2CN0_sign => VN_sign_out(9462),
        VN2CN1_sign => VN_sign_out(9463),
        VN2CN2_sign => VN_sign_out(9464),
        VN2CN3_sign => VN_sign_out(9465),
        VN2CN4_sign => VN_sign_out(9466),
        VN2CN5_sign => VN_sign_out(9467),
        codeword => codeword(1577),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1578 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9473 downto 9468),
        Din0 => VN1578_in0,
        Din1 => VN1578_in1,
        Din2 => VN1578_in2,
        Din3 => VN1578_in3,
        Din4 => VN1578_in4,
        Din5 => VN1578_in5,
        VN2CN0_bit => VN_data_out(9468),
        VN2CN1_bit => VN_data_out(9469),
        VN2CN2_bit => VN_data_out(9470),
        VN2CN3_bit => VN_data_out(9471),
        VN2CN4_bit => VN_data_out(9472),
        VN2CN5_bit => VN_data_out(9473),
        VN2CN0_sign => VN_sign_out(9468),
        VN2CN1_sign => VN_sign_out(9469),
        VN2CN2_sign => VN_sign_out(9470),
        VN2CN3_sign => VN_sign_out(9471),
        VN2CN4_sign => VN_sign_out(9472),
        VN2CN5_sign => VN_sign_out(9473),
        codeword => codeword(1578),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1579 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9479 downto 9474),
        Din0 => VN1579_in0,
        Din1 => VN1579_in1,
        Din2 => VN1579_in2,
        Din3 => VN1579_in3,
        Din4 => VN1579_in4,
        Din5 => VN1579_in5,
        VN2CN0_bit => VN_data_out(9474),
        VN2CN1_bit => VN_data_out(9475),
        VN2CN2_bit => VN_data_out(9476),
        VN2CN3_bit => VN_data_out(9477),
        VN2CN4_bit => VN_data_out(9478),
        VN2CN5_bit => VN_data_out(9479),
        VN2CN0_sign => VN_sign_out(9474),
        VN2CN1_sign => VN_sign_out(9475),
        VN2CN2_sign => VN_sign_out(9476),
        VN2CN3_sign => VN_sign_out(9477),
        VN2CN4_sign => VN_sign_out(9478),
        VN2CN5_sign => VN_sign_out(9479),
        codeword => codeword(1579),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1580 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9485 downto 9480),
        Din0 => VN1580_in0,
        Din1 => VN1580_in1,
        Din2 => VN1580_in2,
        Din3 => VN1580_in3,
        Din4 => VN1580_in4,
        Din5 => VN1580_in5,
        VN2CN0_bit => VN_data_out(9480),
        VN2CN1_bit => VN_data_out(9481),
        VN2CN2_bit => VN_data_out(9482),
        VN2CN3_bit => VN_data_out(9483),
        VN2CN4_bit => VN_data_out(9484),
        VN2CN5_bit => VN_data_out(9485),
        VN2CN0_sign => VN_sign_out(9480),
        VN2CN1_sign => VN_sign_out(9481),
        VN2CN2_sign => VN_sign_out(9482),
        VN2CN3_sign => VN_sign_out(9483),
        VN2CN4_sign => VN_sign_out(9484),
        VN2CN5_sign => VN_sign_out(9485),
        codeword => codeword(1580),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1581 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9491 downto 9486),
        Din0 => VN1581_in0,
        Din1 => VN1581_in1,
        Din2 => VN1581_in2,
        Din3 => VN1581_in3,
        Din4 => VN1581_in4,
        Din5 => VN1581_in5,
        VN2CN0_bit => VN_data_out(9486),
        VN2CN1_bit => VN_data_out(9487),
        VN2CN2_bit => VN_data_out(9488),
        VN2CN3_bit => VN_data_out(9489),
        VN2CN4_bit => VN_data_out(9490),
        VN2CN5_bit => VN_data_out(9491),
        VN2CN0_sign => VN_sign_out(9486),
        VN2CN1_sign => VN_sign_out(9487),
        VN2CN2_sign => VN_sign_out(9488),
        VN2CN3_sign => VN_sign_out(9489),
        VN2CN4_sign => VN_sign_out(9490),
        VN2CN5_sign => VN_sign_out(9491),
        codeword => codeword(1581),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1582 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9497 downto 9492),
        Din0 => VN1582_in0,
        Din1 => VN1582_in1,
        Din2 => VN1582_in2,
        Din3 => VN1582_in3,
        Din4 => VN1582_in4,
        Din5 => VN1582_in5,
        VN2CN0_bit => VN_data_out(9492),
        VN2CN1_bit => VN_data_out(9493),
        VN2CN2_bit => VN_data_out(9494),
        VN2CN3_bit => VN_data_out(9495),
        VN2CN4_bit => VN_data_out(9496),
        VN2CN5_bit => VN_data_out(9497),
        VN2CN0_sign => VN_sign_out(9492),
        VN2CN1_sign => VN_sign_out(9493),
        VN2CN2_sign => VN_sign_out(9494),
        VN2CN3_sign => VN_sign_out(9495),
        VN2CN4_sign => VN_sign_out(9496),
        VN2CN5_sign => VN_sign_out(9497),
        codeword => codeword(1582),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1583 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9503 downto 9498),
        Din0 => VN1583_in0,
        Din1 => VN1583_in1,
        Din2 => VN1583_in2,
        Din3 => VN1583_in3,
        Din4 => VN1583_in4,
        Din5 => VN1583_in5,
        VN2CN0_bit => VN_data_out(9498),
        VN2CN1_bit => VN_data_out(9499),
        VN2CN2_bit => VN_data_out(9500),
        VN2CN3_bit => VN_data_out(9501),
        VN2CN4_bit => VN_data_out(9502),
        VN2CN5_bit => VN_data_out(9503),
        VN2CN0_sign => VN_sign_out(9498),
        VN2CN1_sign => VN_sign_out(9499),
        VN2CN2_sign => VN_sign_out(9500),
        VN2CN3_sign => VN_sign_out(9501),
        VN2CN4_sign => VN_sign_out(9502),
        VN2CN5_sign => VN_sign_out(9503),
        codeword => codeword(1583),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1584 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9509 downto 9504),
        Din0 => VN1584_in0,
        Din1 => VN1584_in1,
        Din2 => VN1584_in2,
        Din3 => VN1584_in3,
        Din4 => VN1584_in4,
        Din5 => VN1584_in5,
        VN2CN0_bit => VN_data_out(9504),
        VN2CN1_bit => VN_data_out(9505),
        VN2CN2_bit => VN_data_out(9506),
        VN2CN3_bit => VN_data_out(9507),
        VN2CN4_bit => VN_data_out(9508),
        VN2CN5_bit => VN_data_out(9509),
        VN2CN0_sign => VN_sign_out(9504),
        VN2CN1_sign => VN_sign_out(9505),
        VN2CN2_sign => VN_sign_out(9506),
        VN2CN3_sign => VN_sign_out(9507),
        VN2CN4_sign => VN_sign_out(9508),
        VN2CN5_sign => VN_sign_out(9509),
        codeword => codeword(1584),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1585 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9515 downto 9510),
        Din0 => VN1585_in0,
        Din1 => VN1585_in1,
        Din2 => VN1585_in2,
        Din3 => VN1585_in3,
        Din4 => VN1585_in4,
        Din5 => VN1585_in5,
        VN2CN0_bit => VN_data_out(9510),
        VN2CN1_bit => VN_data_out(9511),
        VN2CN2_bit => VN_data_out(9512),
        VN2CN3_bit => VN_data_out(9513),
        VN2CN4_bit => VN_data_out(9514),
        VN2CN5_bit => VN_data_out(9515),
        VN2CN0_sign => VN_sign_out(9510),
        VN2CN1_sign => VN_sign_out(9511),
        VN2CN2_sign => VN_sign_out(9512),
        VN2CN3_sign => VN_sign_out(9513),
        VN2CN4_sign => VN_sign_out(9514),
        VN2CN5_sign => VN_sign_out(9515),
        codeword => codeword(1585),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1586 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9521 downto 9516),
        Din0 => VN1586_in0,
        Din1 => VN1586_in1,
        Din2 => VN1586_in2,
        Din3 => VN1586_in3,
        Din4 => VN1586_in4,
        Din5 => VN1586_in5,
        VN2CN0_bit => VN_data_out(9516),
        VN2CN1_bit => VN_data_out(9517),
        VN2CN2_bit => VN_data_out(9518),
        VN2CN3_bit => VN_data_out(9519),
        VN2CN4_bit => VN_data_out(9520),
        VN2CN5_bit => VN_data_out(9521),
        VN2CN0_sign => VN_sign_out(9516),
        VN2CN1_sign => VN_sign_out(9517),
        VN2CN2_sign => VN_sign_out(9518),
        VN2CN3_sign => VN_sign_out(9519),
        VN2CN4_sign => VN_sign_out(9520),
        VN2CN5_sign => VN_sign_out(9521),
        codeword => codeword(1586),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1587 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9527 downto 9522),
        Din0 => VN1587_in0,
        Din1 => VN1587_in1,
        Din2 => VN1587_in2,
        Din3 => VN1587_in3,
        Din4 => VN1587_in4,
        Din5 => VN1587_in5,
        VN2CN0_bit => VN_data_out(9522),
        VN2CN1_bit => VN_data_out(9523),
        VN2CN2_bit => VN_data_out(9524),
        VN2CN3_bit => VN_data_out(9525),
        VN2CN4_bit => VN_data_out(9526),
        VN2CN5_bit => VN_data_out(9527),
        VN2CN0_sign => VN_sign_out(9522),
        VN2CN1_sign => VN_sign_out(9523),
        VN2CN2_sign => VN_sign_out(9524),
        VN2CN3_sign => VN_sign_out(9525),
        VN2CN4_sign => VN_sign_out(9526),
        VN2CN5_sign => VN_sign_out(9527),
        codeword => codeword(1587),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1588 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9533 downto 9528),
        Din0 => VN1588_in0,
        Din1 => VN1588_in1,
        Din2 => VN1588_in2,
        Din3 => VN1588_in3,
        Din4 => VN1588_in4,
        Din5 => VN1588_in5,
        VN2CN0_bit => VN_data_out(9528),
        VN2CN1_bit => VN_data_out(9529),
        VN2CN2_bit => VN_data_out(9530),
        VN2CN3_bit => VN_data_out(9531),
        VN2CN4_bit => VN_data_out(9532),
        VN2CN5_bit => VN_data_out(9533),
        VN2CN0_sign => VN_sign_out(9528),
        VN2CN1_sign => VN_sign_out(9529),
        VN2CN2_sign => VN_sign_out(9530),
        VN2CN3_sign => VN_sign_out(9531),
        VN2CN4_sign => VN_sign_out(9532),
        VN2CN5_sign => VN_sign_out(9533),
        codeword => codeword(1588),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1589 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9539 downto 9534),
        Din0 => VN1589_in0,
        Din1 => VN1589_in1,
        Din2 => VN1589_in2,
        Din3 => VN1589_in3,
        Din4 => VN1589_in4,
        Din5 => VN1589_in5,
        VN2CN0_bit => VN_data_out(9534),
        VN2CN1_bit => VN_data_out(9535),
        VN2CN2_bit => VN_data_out(9536),
        VN2CN3_bit => VN_data_out(9537),
        VN2CN4_bit => VN_data_out(9538),
        VN2CN5_bit => VN_data_out(9539),
        VN2CN0_sign => VN_sign_out(9534),
        VN2CN1_sign => VN_sign_out(9535),
        VN2CN2_sign => VN_sign_out(9536),
        VN2CN3_sign => VN_sign_out(9537),
        VN2CN4_sign => VN_sign_out(9538),
        VN2CN5_sign => VN_sign_out(9539),
        codeword => codeword(1589),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1590 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9545 downto 9540),
        Din0 => VN1590_in0,
        Din1 => VN1590_in1,
        Din2 => VN1590_in2,
        Din3 => VN1590_in3,
        Din4 => VN1590_in4,
        Din5 => VN1590_in5,
        VN2CN0_bit => VN_data_out(9540),
        VN2CN1_bit => VN_data_out(9541),
        VN2CN2_bit => VN_data_out(9542),
        VN2CN3_bit => VN_data_out(9543),
        VN2CN4_bit => VN_data_out(9544),
        VN2CN5_bit => VN_data_out(9545),
        VN2CN0_sign => VN_sign_out(9540),
        VN2CN1_sign => VN_sign_out(9541),
        VN2CN2_sign => VN_sign_out(9542),
        VN2CN3_sign => VN_sign_out(9543),
        VN2CN4_sign => VN_sign_out(9544),
        VN2CN5_sign => VN_sign_out(9545),
        codeword => codeword(1590),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1591 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9551 downto 9546),
        Din0 => VN1591_in0,
        Din1 => VN1591_in1,
        Din2 => VN1591_in2,
        Din3 => VN1591_in3,
        Din4 => VN1591_in4,
        Din5 => VN1591_in5,
        VN2CN0_bit => VN_data_out(9546),
        VN2CN1_bit => VN_data_out(9547),
        VN2CN2_bit => VN_data_out(9548),
        VN2CN3_bit => VN_data_out(9549),
        VN2CN4_bit => VN_data_out(9550),
        VN2CN5_bit => VN_data_out(9551),
        VN2CN0_sign => VN_sign_out(9546),
        VN2CN1_sign => VN_sign_out(9547),
        VN2CN2_sign => VN_sign_out(9548),
        VN2CN3_sign => VN_sign_out(9549),
        VN2CN4_sign => VN_sign_out(9550),
        VN2CN5_sign => VN_sign_out(9551),
        codeword => codeword(1591),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1592 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9557 downto 9552),
        Din0 => VN1592_in0,
        Din1 => VN1592_in1,
        Din2 => VN1592_in2,
        Din3 => VN1592_in3,
        Din4 => VN1592_in4,
        Din5 => VN1592_in5,
        VN2CN0_bit => VN_data_out(9552),
        VN2CN1_bit => VN_data_out(9553),
        VN2CN2_bit => VN_data_out(9554),
        VN2CN3_bit => VN_data_out(9555),
        VN2CN4_bit => VN_data_out(9556),
        VN2CN5_bit => VN_data_out(9557),
        VN2CN0_sign => VN_sign_out(9552),
        VN2CN1_sign => VN_sign_out(9553),
        VN2CN2_sign => VN_sign_out(9554),
        VN2CN3_sign => VN_sign_out(9555),
        VN2CN4_sign => VN_sign_out(9556),
        VN2CN5_sign => VN_sign_out(9557),
        codeword => codeword(1592),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1593 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9563 downto 9558),
        Din0 => VN1593_in0,
        Din1 => VN1593_in1,
        Din2 => VN1593_in2,
        Din3 => VN1593_in3,
        Din4 => VN1593_in4,
        Din5 => VN1593_in5,
        VN2CN0_bit => VN_data_out(9558),
        VN2CN1_bit => VN_data_out(9559),
        VN2CN2_bit => VN_data_out(9560),
        VN2CN3_bit => VN_data_out(9561),
        VN2CN4_bit => VN_data_out(9562),
        VN2CN5_bit => VN_data_out(9563),
        VN2CN0_sign => VN_sign_out(9558),
        VN2CN1_sign => VN_sign_out(9559),
        VN2CN2_sign => VN_sign_out(9560),
        VN2CN3_sign => VN_sign_out(9561),
        VN2CN4_sign => VN_sign_out(9562),
        VN2CN5_sign => VN_sign_out(9563),
        codeword => codeword(1593),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1594 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9569 downto 9564),
        Din0 => VN1594_in0,
        Din1 => VN1594_in1,
        Din2 => VN1594_in2,
        Din3 => VN1594_in3,
        Din4 => VN1594_in4,
        Din5 => VN1594_in5,
        VN2CN0_bit => VN_data_out(9564),
        VN2CN1_bit => VN_data_out(9565),
        VN2CN2_bit => VN_data_out(9566),
        VN2CN3_bit => VN_data_out(9567),
        VN2CN4_bit => VN_data_out(9568),
        VN2CN5_bit => VN_data_out(9569),
        VN2CN0_sign => VN_sign_out(9564),
        VN2CN1_sign => VN_sign_out(9565),
        VN2CN2_sign => VN_sign_out(9566),
        VN2CN3_sign => VN_sign_out(9567),
        VN2CN4_sign => VN_sign_out(9568),
        VN2CN5_sign => VN_sign_out(9569),
        codeword => codeword(1594),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1595 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9575 downto 9570),
        Din0 => VN1595_in0,
        Din1 => VN1595_in1,
        Din2 => VN1595_in2,
        Din3 => VN1595_in3,
        Din4 => VN1595_in4,
        Din5 => VN1595_in5,
        VN2CN0_bit => VN_data_out(9570),
        VN2CN1_bit => VN_data_out(9571),
        VN2CN2_bit => VN_data_out(9572),
        VN2CN3_bit => VN_data_out(9573),
        VN2CN4_bit => VN_data_out(9574),
        VN2CN5_bit => VN_data_out(9575),
        VN2CN0_sign => VN_sign_out(9570),
        VN2CN1_sign => VN_sign_out(9571),
        VN2CN2_sign => VN_sign_out(9572),
        VN2CN3_sign => VN_sign_out(9573),
        VN2CN4_sign => VN_sign_out(9574),
        VN2CN5_sign => VN_sign_out(9575),
        codeword => codeword(1595),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1596 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9581 downto 9576),
        Din0 => VN1596_in0,
        Din1 => VN1596_in1,
        Din2 => VN1596_in2,
        Din3 => VN1596_in3,
        Din4 => VN1596_in4,
        Din5 => VN1596_in5,
        VN2CN0_bit => VN_data_out(9576),
        VN2CN1_bit => VN_data_out(9577),
        VN2CN2_bit => VN_data_out(9578),
        VN2CN3_bit => VN_data_out(9579),
        VN2CN4_bit => VN_data_out(9580),
        VN2CN5_bit => VN_data_out(9581),
        VN2CN0_sign => VN_sign_out(9576),
        VN2CN1_sign => VN_sign_out(9577),
        VN2CN2_sign => VN_sign_out(9578),
        VN2CN3_sign => VN_sign_out(9579),
        VN2CN4_sign => VN_sign_out(9580),
        VN2CN5_sign => VN_sign_out(9581),
        codeword => codeword(1596),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1597 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9587 downto 9582),
        Din0 => VN1597_in0,
        Din1 => VN1597_in1,
        Din2 => VN1597_in2,
        Din3 => VN1597_in3,
        Din4 => VN1597_in4,
        Din5 => VN1597_in5,
        VN2CN0_bit => VN_data_out(9582),
        VN2CN1_bit => VN_data_out(9583),
        VN2CN2_bit => VN_data_out(9584),
        VN2CN3_bit => VN_data_out(9585),
        VN2CN4_bit => VN_data_out(9586),
        VN2CN5_bit => VN_data_out(9587),
        VN2CN0_sign => VN_sign_out(9582),
        VN2CN1_sign => VN_sign_out(9583),
        VN2CN2_sign => VN_sign_out(9584),
        VN2CN3_sign => VN_sign_out(9585),
        VN2CN4_sign => VN_sign_out(9586),
        VN2CN5_sign => VN_sign_out(9587),
        codeword => codeword(1597),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1598 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9593 downto 9588),
        Din0 => VN1598_in0,
        Din1 => VN1598_in1,
        Din2 => VN1598_in2,
        Din3 => VN1598_in3,
        Din4 => VN1598_in4,
        Din5 => VN1598_in5,
        VN2CN0_bit => VN_data_out(9588),
        VN2CN1_bit => VN_data_out(9589),
        VN2CN2_bit => VN_data_out(9590),
        VN2CN3_bit => VN_data_out(9591),
        VN2CN4_bit => VN_data_out(9592),
        VN2CN5_bit => VN_data_out(9593),
        VN2CN0_sign => VN_sign_out(9588),
        VN2CN1_sign => VN_sign_out(9589),
        VN2CN2_sign => VN_sign_out(9590),
        VN2CN3_sign => VN_sign_out(9591),
        VN2CN4_sign => VN_sign_out(9592),
        VN2CN5_sign => VN_sign_out(9593),
        codeword => codeword(1598),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1599 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9599 downto 9594),
        Din0 => VN1599_in0,
        Din1 => VN1599_in1,
        Din2 => VN1599_in2,
        Din3 => VN1599_in3,
        Din4 => VN1599_in4,
        Din5 => VN1599_in5,
        VN2CN0_bit => VN_data_out(9594),
        VN2CN1_bit => VN_data_out(9595),
        VN2CN2_bit => VN_data_out(9596),
        VN2CN3_bit => VN_data_out(9597),
        VN2CN4_bit => VN_data_out(9598),
        VN2CN5_bit => VN_data_out(9599),
        VN2CN0_sign => VN_sign_out(9594),
        VN2CN1_sign => VN_sign_out(9595),
        VN2CN2_sign => VN_sign_out(9596),
        VN2CN3_sign => VN_sign_out(9597),
        VN2CN4_sign => VN_sign_out(9598),
        VN2CN5_sign => VN_sign_out(9599),
        codeword => codeword(1599),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1600 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9605 downto 9600),
        Din0 => VN1600_in0,
        Din1 => VN1600_in1,
        Din2 => VN1600_in2,
        Din3 => VN1600_in3,
        Din4 => VN1600_in4,
        Din5 => VN1600_in5,
        VN2CN0_bit => VN_data_out(9600),
        VN2CN1_bit => VN_data_out(9601),
        VN2CN2_bit => VN_data_out(9602),
        VN2CN3_bit => VN_data_out(9603),
        VN2CN4_bit => VN_data_out(9604),
        VN2CN5_bit => VN_data_out(9605),
        VN2CN0_sign => VN_sign_out(9600),
        VN2CN1_sign => VN_sign_out(9601),
        VN2CN2_sign => VN_sign_out(9602),
        VN2CN3_sign => VN_sign_out(9603),
        VN2CN4_sign => VN_sign_out(9604),
        VN2CN5_sign => VN_sign_out(9605),
        codeword => codeword(1600),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1601 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9611 downto 9606),
        Din0 => VN1601_in0,
        Din1 => VN1601_in1,
        Din2 => VN1601_in2,
        Din3 => VN1601_in3,
        Din4 => VN1601_in4,
        Din5 => VN1601_in5,
        VN2CN0_bit => VN_data_out(9606),
        VN2CN1_bit => VN_data_out(9607),
        VN2CN2_bit => VN_data_out(9608),
        VN2CN3_bit => VN_data_out(9609),
        VN2CN4_bit => VN_data_out(9610),
        VN2CN5_bit => VN_data_out(9611),
        VN2CN0_sign => VN_sign_out(9606),
        VN2CN1_sign => VN_sign_out(9607),
        VN2CN2_sign => VN_sign_out(9608),
        VN2CN3_sign => VN_sign_out(9609),
        VN2CN4_sign => VN_sign_out(9610),
        VN2CN5_sign => VN_sign_out(9611),
        codeword => codeword(1601),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1602 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9617 downto 9612),
        Din0 => VN1602_in0,
        Din1 => VN1602_in1,
        Din2 => VN1602_in2,
        Din3 => VN1602_in3,
        Din4 => VN1602_in4,
        Din5 => VN1602_in5,
        VN2CN0_bit => VN_data_out(9612),
        VN2CN1_bit => VN_data_out(9613),
        VN2CN2_bit => VN_data_out(9614),
        VN2CN3_bit => VN_data_out(9615),
        VN2CN4_bit => VN_data_out(9616),
        VN2CN5_bit => VN_data_out(9617),
        VN2CN0_sign => VN_sign_out(9612),
        VN2CN1_sign => VN_sign_out(9613),
        VN2CN2_sign => VN_sign_out(9614),
        VN2CN3_sign => VN_sign_out(9615),
        VN2CN4_sign => VN_sign_out(9616),
        VN2CN5_sign => VN_sign_out(9617),
        codeword => codeword(1602),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1603 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9623 downto 9618),
        Din0 => VN1603_in0,
        Din1 => VN1603_in1,
        Din2 => VN1603_in2,
        Din3 => VN1603_in3,
        Din4 => VN1603_in4,
        Din5 => VN1603_in5,
        VN2CN0_bit => VN_data_out(9618),
        VN2CN1_bit => VN_data_out(9619),
        VN2CN2_bit => VN_data_out(9620),
        VN2CN3_bit => VN_data_out(9621),
        VN2CN4_bit => VN_data_out(9622),
        VN2CN5_bit => VN_data_out(9623),
        VN2CN0_sign => VN_sign_out(9618),
        VN2CN1_sign => VN_sign_out(9619),
        VN2CN2_sign => VN_sign_out(9620),
        VN2CN3_sign => VN_sign_out(9621),
        VN2CN4_sign => VN_sign_out(9622),
        VN2CN5_sign => VN_sign_out(9623),
        codeword => codeword(1603),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1604 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9629 downto 9624),
        Din0 => VN1604_in0,
        Din1 => VN1604_in1,
        Din2 => VN1604_in2,
        Din3 => VN1604_in3,
        Din4 => VN1604_in4,
        Din5 => VN1604_in5,
        VN2CN0_bit => VN_data_out(9624),
        VN2CN1_bit => VN_data_out(9625),
        VN2CN2_bit => VN_data_out(9626),
        VN2CN3_bit => VN_data_out(9627),
        VN2CN4_bit => VN_data_out(9628),
        VN2CN5_bit => VN_data_out(9629),
        VN2CN0_sign => VN_sign_out(9624),
        VN2CN1_sign => VN_sign_out(9625),
        VN2CN2_sign => VN_sign_out(9626),
        VN2CN3_sign => VN_sign_out(9627),
        VN2CN4_sign => VN_sign_out(9628),
        VN2CN5_sign => VN_sign_out(9629),
        codeword => codeword(1604),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1605 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9635 downto 9630),
        Din0 => VN1605_in0,
        Din1 => VN1605_in1,
        Din2 => VN1605_in2,
        Din3 => VN1605_in3,
        Din4 => VN1605_in4,
        Din5 => VN1605_in5,
        VN2CN0_bit => VN_data_out(9630),
        VN2CN1_bit => VN_data_out(9631),
        VN2CN2_bit => VN_data_out(9632),
        VN2CN3_bit => VN_data_out(9633),
        VN2CN4_bit => VN_data_out(9634),
        VN2CN5_bit => VN_data_out(9635),
        VN2CN0_sign => VN_sign_out(9630),
        VN2CN1_sign => VN_sign_out(9631),
        VN2CN2_sign => VN_sign_out(9632),
        VN2CN3_sign => VN_sign_out(9633),
        VN2CN4_sign => VN_sign_out(9634),
        VN2CN5_sign => VN_sign_out(9635),
        codeword => codeword(1605),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1606 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9641 downto 9636),
        Din0 => VN1606_in0,
        Din1 => VN1606_in1,
        Din2 => VN1606_in2,
        Din3 => VN1606_in3,
        Din4 => VN1606_in4,
        Din5 => VN1606_in5,
        VN2CN0_bit => VN_data_out(9636),
        VN2CN1_bit => VN_data_out(9637),
        VN2CN2_bit => VN_data_out(9638),
        VN2CN3_bit => VN_data_out(9639),
        VN2CN4_bit => VN_data_out(9640),
        VN2CN5_bit => VN_data_out(9641),
        VN2CN0_sign => VN_sign_out(9636),
        VN2CN1_sign => VN_sign_out(9637),
        VN2CN2_sign => VN_sign_out(9638),
        VN2CN3_sign => VN_sign_out(9639),
        VN2CN4_sign => VN_sign_out(9640),
        VN2CN5_sign => VN_sign_out(9641),
        codeword => codeword(1606),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1607 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9647 downto 9642),
        Din0 => VN1607_in0,
        Din1 => VN1607_in1,
        Din2 => VN1607_in2,
        Din3 => VN1607_in3,
        Din4 => VN1607_in4,
        Din5 => VN1607_in5,
        VN2CN0_bit => VN_data_out(9642),
        VN2CN1_bit => VN_data_out(9643),
        VN2CN2_bit => VN_data_out(9644),
        VN2CN3_bit => VN_data_out(9645),
        VN2CN4_bit => VN_data_out(9646),
        VN2CN5_bit => VN_data_out(9647),
        VN2CN0_sign => VN_sign_out(9642),
        VN2CN1_sign => VN_sign_out(9643),
        VN2CN2_sign => VN_sign_out(9644),
        VN2CN3_sign => VN_sign_out(9645),
        VN2CN4_sign => VN_sign_out(9646),
        VN2CN5_sign => VN_sign_out(9647),
        codeword => codeword(1607),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1608 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9653 downto 9648),
        Din0 => VN1608_in0,
        Din1 => VN1608_in1,
        Din2 => VN1608_in2,
        Din3 => VN1608_in3,
        Din4 => VN1608_in4,
        Din5 => VN1608_in5,
        VN2CN0_bit => VN_data_out(9648),
        VN2CN1_bit => VN_data_out(9649),
        VN2CN2_bit => VN_data_out(9650),
        VN2CN3_bit => VN_data_out(9651),
        VN2CN4_bit => VN_data_out(9652),
        VN2CN5_bit => VN_data_out(9653),
        VN2CN0_sign => VN_sign_out(9648),
        VN2CN1_sign => VN_sign_out(9649),
        VN2CN2_sign => VN_sign_out(9650),
        VN2CN3_sign => VN_sign_out(9651),
        VN2CN4_sign => VN_sign_out(9652),
        VN2CN5_sign => VN_sign_out(9653),
        codeword => codeword(1608),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1609 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9659 downto 9654),
        Din0 => VN1609_in0,
        Din1 => VN1609_in1,
        Din2 => VN1609_in2,
        Din3 => VN1609_in3,
        Din4 => VN1609_in4,
        Din5 => VN1609_in5,
        VN2CN0_bit => VN_data_out(9654),
        VN2CN1_bit => VN_data_out(9655),
        VN2CN2_bit => VN_data_out(9656),
        VN2CN3_bit => VN_data_out(9657),
        VN2CN4_bit => VN_data_out(9658),
        VN2CN5_bit => VN_data_out(9659),
        VN2CN0_sign => VN_sign_out(9654),
        VN2CN1_sign => VN_sign_out(9655),
        VN2CN2_sign => VN_sign_out(9656),
        VN2CN3_sign => VN_sign_out(9657),
        VN2CN4_sign => VN_sign_out(9658),
        VN2CN5_sign => VN_sign_out(9659),
        codeword => codeword(1609),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1610 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9665 downto 9660),
        Din0 => VN1610_in0,
        Din1 => VN1610_in1,
        Din2 => VN1610_in2,
        Din3 => VN1610_in3,
        Din4 => VN1610_in4,
        Din5 => VN1610_in5,
        VN2CN0_bit => VN_data_out(9660),
        VN2CN1_bit => VN_data_out(9661),
        VN2CN2_bit => VN_data_out(9662),
        VN2CN3_bit => VN_data_out(9663),
        VN2CN4_bit => VN_data_out(9664),
        VN2CN5_bit => VN_data_out(9665),
        VN2CN0_sign => VN_sign_out(9660),
        VN2CN1_sign => VN_sign_out(9661),
        VN2CN2_sign => VN_sign_out(9662),
        VN2CN3_sign => VN_sign_out(9663),
        VN2CN4_sign => VN_sign_out(9664),
        VN2CN5_sign => VN_sign_out(9665),
        codeword => codeword(1610),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1611 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9671 downto 9666),
        Din0 => VN1611_in0,
        Din1 => VN1611_in1,
        Din2 => VN1611_in2,
        Din3 => VN1611_in3,
        Din4 => VN1611_in4,
        Din5 => VN1611_in5,
        VN2CN0_bit => VN_data_out(9666),
        VN2CN1_bit => VN_data_out(9667),
        VN2CN2_bit => VN_data_out(9668),
        VN2CN3_bit => VN_data_out(9669),
        VN2CN4_bit => VN_data_out(9670),
        VN2CN5_bit => VN_data_out(9671),
        VN2CN0_sign => VN_sign_out(9666),
        VN2CN1_sign => VN_sign_out(9667),
        VN2CN2_sign => VN_sign_out(9668),
        VN2CN3_sign => VN_sign_out(9669),
        VN2CN4_sign => VN_sign_out(9670),
        VN2CN5_sign => VN_sign_out(9671),
        codeword => codeword(1611),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1612 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9677 downto 9672),
        Din0 => VN1612_in0,
        Din1 => VN1612_in1,
        Din2 => VN1612_in2,
        Din3 => VN1612_in3,
        Din4 => VN1612_in4,
        Din5 => VN1612_in5,
        VN2CN0_bit => VN_data_out(9672),
        VN2CN1_bit => VN_data_out(9673),
        VN2CN2_bit => VN_data_out(9674),
        VN2CN3_bit => VN_data_out(9675),
        VN2CN4_bit => VN_data_out(9676),
        VN2CN5_bit => VN_data_out(9677),
        VN2CN0_sign => VN_sign_out(9672),
        VN2CN1_sign => VN_sign_out(9673),
        VN2CN2_sign => VN_sign_out(9674),
        VN2CN3_sign => VN_sign_out(9675),
        VN2CN4_sign => VN_sign_out(9676),
        VN2CN5_sign => VN_sign_out(9677),
        codeword => codeword(1612),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1613 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9683 downto 9678),
        Din0 => VN1613_in0,
        Din1 => VN1613_in1,
        Din2 => VN1613_in2,
        Din3 => VN1613_in3,
        Din4 => VN1613_in4,
        Din5 => VN1613_in5,
        VN2CN0_bit => VN_data_out(9678),
        VN2CN1_bit => VN_data_out(9679),
        VN2CN2_bit => VN_data_out(9680),
        VN2CN3_bit => VN_data_out(9681),
        VN2CN4_bit => VN_data_out(9682),
        VN2CN5_bit => VN_data_out(9683),
        VN2CN0_sign => VN_sign_out(9678),
        VN2CN1_sign => VN_sign_out(9679),
        VN2CN2_sign => VN_sign_out(9680),
        VN2CN3_sign => VN_sign_out(9681),
        VN2CN4_sign => VN_sign_out(9682),
        VN2CN5_sign => VN_sign_out(9683),
        codeword => codeword(1613),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1614 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9689 downto 9684),
        Din0 => VN1614_in0,
        Din1 => VN1614_in1,
        Din2 => VN1614_in2,
        Din3 => VN1614_in3,
        Din4 => VN1614_in4,
        Din5 => VN1614_in5,
        VN2CN0_bit => VN_data_out(9684),
        VN2CN1_bit => VN_data_out(9685),
        VN2CN2_bit => VN_data_out(9686),
        VN2CN3_bit => VN_data_out(9687),
        VN2CN4_bit => VN_data_out(9688),
        VN2CN5_bit => VN_data_out(9689),
        VN2CN0_sign => VN_sign_out(9684),
        VN2CN1_sign => VN_sign_out(9685),
        VN2CN2_sign => VN_sign_out(9686),
        VN2CN3_sign => VN_sign_out(9687),
        VN2CN4_sign => VN_sign_out(9688),
        VN2CN5_sign => VN_sign_out(9689),
        codeword => codeword(1614),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1615 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9695 downto 9690),
        Din0 => VN1615_in0,
        Din1 => VN1615_in1,
        Din2 => VN1615_in2,
        Din3 => VN1615_in3,
        Din4 => VN1615_in4,
        Din5 => VN1615_in5,
        VN2CN0_bit => VN_data_out(9690),
        VN2CN1_bit => VN_data_out(9691),
        VN2CN2_bit => VN_data_out(9692),
        VN2CN3_bit => VN_data_out(9693),
        VN2CN4_bit => VN_data_out(9694),
        VN2CN5_bit => VN_data_out(9695),
        VN2CN0_sign => VN_sign_out(9690),
        VN2CN1_sign => VN_sign_out(9691),
        VN2CN2_sign => VN_sign_out(9692),
        VN2CN3_sign => VN_sign_out(9693),
        VN2CN4_sign => VN_sign_out(9694),
        VN2CN5_sign => VN_sign_out(9695),
        codeword => codeword(1615),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1616 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9701 downto 9696),
        Din0 => VN1616_in0,
        Din1 => VN1616_in1,
        Din2 => VN1616_in2,
        Din3 => VN1616_in3,
        Din4 => VN1616_in4,
        Din5 => VN1616_in5,
        VN2CN0_bit => VN_data_out(9696),
        VN2CN1_bit => VN_data_out(9697),
        VN2CN2_bit => VN_data_out(9698),
        VN2CN3_bit => VN_data_out(9699),
        VN2CN4_bit => VN_data_out(9700),
        VN2CN5_bit => VN_data_out(9701),
        VN2CN0_sign => VN_sign_out(9696),
        VN2CN1_sign => VN_sign_out(9697),
        VN2CN2_sign => VN_sign_out(9698),
        VN2CN3_sign => VN_sign_out(9699),
        VN2CN4_sign => VN_sign_out(9700),
        VN2CN5_sign => VN_sign_out(9701),
        codeword => codeword(1616),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1617 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9707 downto 9702),
        Din0 => VN1617_in0,
        Din1 => VN1617_in1,
        Din2 => VN1617_in2,
        Din3 => VN1617_in3,
        Din4 => VN1617_in4,
        Din5 => VN1617_in5,
        VN2CN0_bit => VN_data_out(9702),
        VN2CN1_bit => VN_data_out(9703),
        VN2CN2_bit => VN_data_out(9704),
        VN2CN3_bit => VN_data_out(9705),
        VN2CN4_bit => VN_data_out(9706),
        VN2CN5_bit => VN_data_out(9707),
        VN2CN0_sign => VN_sign_out(9702),
        VN2CN1_sign => VN_sign_out(9703),
        VN2CN2_sign => VN_sign_out(9704),
        VN2CN3_sign => VN_sign_out(9705),
        VN2CN4_sign => VN_sign_out(9706),
        VN2CN5_sign => VN_sign_out(9707),
        codeword => codeword(1617),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1618 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9713 downto 9708),
        Din0 => VN1618_in0,
        Din1 => VN1618_in1,
        Din2 => VN1618_in2,
        Din3 => VN1618_in3,
        Din4 => VN1618_in4,
        Din5 => VN1618_in5,
        VN2CN0_bit => VN_data_out(9708),
        VN2CN1_bit => VN_data_out(9709),
        VN2CN2_bit => VN_data_out(9710),
        VN2CN3_bit => VN_data_out(9711),
        VN2CN4_bit => VN_data_out(9712),
        VN2CN5_bit => VN_data_out(9713),
        VN2CN0_sign => VN_sign_out(9708),
        VN2CN1_sign => VN_sign_out(9709),
        VN2CN2_sign => VN_sign_out(9710),
        VN2CN3_sign => VN_sign_out(9711),
        VN2CN4_sign => VN_sign_out(9712),
        VN2CN5_sign => VN_sign_out(9713),
        codeword => codeword(1618),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1619 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9719 downto 9714),
        Din0 => VN1619_in0,
        Din1 => VN1619_in1,
        Din2 => VN1619_in2,
        Din3 => VN1619_in3,
        Din4 => VN1619_in4,
        Din5 => VN1619_in5,
        VN2CN0_bit => VN_data_out(9714),
        VN2CN1_bit => VN_data_out(9715),
        VN2CN2_bit => VN_data_out(9716),
        VN2CN3_bit => VN_data_out(9717),
        VN2CN4_bit => VN_data_out(9718),
        VN2CN5_bit => VN_data_out(9719),
        VN2CN0_sign => VN_sign_out(9714),
        VN2CN1_sign => VN_sign_out(9715),
        VN2CN2_sign => VN_sign_out(9716),
        VN2CN3_sign => VN_sign_out(9717),
        VN2CN4_sign => VN_sign_out(9718),
        VN2CN5_sign => VN_sign_out(9719),
        codeword => codeword(1619),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1620 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9725 downto 9720),
        Din0 => VN1620_in0,
        Din1 => VN1620_in1,
        Din2 => VN1620_in2,
        Din3 => VN1620_in3,
        Din4 => VN1620_in4,
        Din5 => VN1620_in5,
        VN2CN0_bit => VN_data_out(9720),
        VN2CN1_bit => VN_data_out(9721),
        VN2CN2_bit => VN_data_out(9722),
        VN2CN3_bit => VN_data_out(9723),
        VN2CN4_bit => VN_data_out(9724),
        VN2CN5_bit => VN_data_out(9725),
        VN2CN0_sign => VN_sign_out(9720),
        VN2CN1_sign => VN_sign_out(9721),
        VN2CN2_sign => VN_sign_out(9722),
        VN2CN3_sign => VN_sign_out(9723),
        VN2CN4_sign => VN_sign_out(9724),
        VN2CN5_sign => VN_sign_out(9725),
        codeword => codeword(1620),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1621 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9731 downto 9726),
        Din0 => VN1621_in0,
        Din1 => VN1621_in1,
        Din2 => VN1621_in2,
        Din3 => VN1621_in3,
        Din4 => VN1621_in4,
        Din5 => VN1621_in5,
        VN2CN0_bit => VN_data_out(9726),
        VN2CN1_bit => VN_data_out(9727),
        VN2CN2_bit => VN_data_out(9728),
        VN2CN3_bit => VN_data_out(9729),
        VN2CN4_bit => VN_data_out(9730),
        VN2CN5_bit => VN_data_out(9731),
        VN2CN0_sign => VN_sign_out(9726),
        VN2CN1_sign => VN_sign_out(9727),
        VN2CN2_sign => VN_sign_out(9728),
        VN2CN3_sign => VN_sign_out(9729),
        VN2CN4_sign => VN_sign_out(9730),
        VN2CN5_sign => VN_sign_out(9731),
        codeword => codeword(1621),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1622 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9737 downto 9732),
        Din0 => VN1622_in0,
        Din1 => VN1622_in1,
        Din2 => VN1622_in2,
        Din3 => VN1622_in3,
        Din4 => VN1622_in4,
        Din5 => VN1622_in5,
        VN2CN0_bit => VN_data_out(9732),
        VN2CN1_bit => VN_data_out(9733),
        VN2CN2_bit => VN_data_out(9734),
        VN2CN3_bit => VN_data_out(9735),
        VN2CN4_bit => VN_data_out(9736),
        VN2CN5_bit => VN_data_out(9737),
        VN2CN0_sign => VN_sign_out(9732),
        VN2CN1_sign => VN_sign_out(9733),
        VN2CN2_sign => VN_sign_out(9734),
        VN2CN3_sign => VN_sign_out(9735),
        VN2CN4_sign => VN_sign_out(9736),
        VN2CN5_sign => VN_sign_out(9737),
        codeword => codeword(1622),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1623 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9743 downto 9738),
        Din0 => VN1623_in0,
        Din1 => VN1623_in1,
        Din2 => VN1623_in2,
        Din3 => VN1623_in3,
        Din4 => VN1623_in4,
        Din5 => VN1623_in5,
        VN2CN0_bit => VN_data_out(9738),
        VN2CN1_bit => VN_data_out(9739),
        VN2CN2_bit => VN_data_out(9740),
        VN2CN3_bit => VN_data_out(9741),
        VN2CN4_bit => VN_data_out(9742),
        VN2CN5_bit => VN_data_out(9743),
        VN2CN0_sign => VN_sign_out(9738),
        VN2CN1_sign => VN_sign_out(9739),
        VN2CN2_sign => VN_sign_out(9740),
        VN2CN3_sign => VN_sign_out(9741),
        VN2CN4_sign => VN_sign_out(9742),
        VN2CN5_sign => VN_sign_out(9743),
        codeword => codeword(1623),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1624 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9749 downto 9744),
        Din0 => VN1624_in0,
        Din1 => VN1624_in1,
        Din2 => VN1624_in2,
        Din3 => VN1624_in3,
        Din4 => VN1624_in4,
        Din5 => VN1624_in5,
        VN2CN0_bit => VN_data_out(9744),
        VN2CN1_bit => VN_data_out(9745),
        VN2CN2_bit => VN_data_out(9746),
        VN2CN3_bit => VN_data_out(9747),
        VN2CN4_bit => VN_data_out(9748),
        VN2CN5_bit => VN_data_out(9749),
        VN2CN0_sign => VN_sign_out(9744),
        VN2CN1_sign => VN_sign_out(9745),
        VN2CN2_sign => VN_sign_out(9746),
        VN2CN3_sign => VN_sign_out(9747),
        VN2CN4_sign => VN_sign_out(9748),
        VN2CN5_sign => VN_sign_out(9749),
        codeword => codeword(1624),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1625 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9755 downto 9750),
        Din0 => VN1625_in0,
        Din1 => VN1625_in1,
        Din2 => VN1625_in2,
        Din3 => VN1625_in3,
        Din4 => VN1625_in4,
        Din5 => VN1625_in5,
        VN2CN0_bit => VN_data_out(9750),
        VN2CN1_bit => VN_data_out(9751),
        VN2CN2_bit => VN_data_out(9752),
        VN2CN3_bit => VN_data_out(9753),
        VN2CN4_bit => VN_data_out(9754),
        VN2CN5_bit => VN_data_out(9755),
        VN2CN0_sign => VN_sign_out(9750),
        VN2CN1_sign => VN_sign_out(9751),
        VN2CN2_sign => VN_sign_out(9752),
        VN2CN3_sign => VN_sign_out(9753),
        VN2CN4_sign => VN_sign_out(9754),
        VN2CN5_sign => VN_sign_out(9755),
        codeword => codeword(1625),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1626 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9761 downto 9756),
        Din0 => VN1626_in0,
        Din1 => VN1626_in1,
        Din2 => VN1626_in2,
        Din3 => VN1626_in3,
        Din4 => VN1626_in4,
        Din5 => VN1626_in5,
        VN2CN0_bit => VN_data_out(9756),
        VN2CN1_bit => VN_data_out(9757),
        VN2CN2_bit => VN_data_out(9758),
        VN2CN3_bit => VN_data_out(9759),
        VN2CN4_bit => VN_data_out(9760),
        VN2CN5_bit => VN_data_out(9761),
        VN2CN0_sign => VN_sign_out(9756),
        VN2CN1_sign => VN_sign_out(9757),
        VN2CN2_sign => VN_sign_out(9758),
        VN2CN3_sign => VN_sign_out(9759),
        VN2CN4_sign => VN_sign_out(9760),
        VN2CN5_sign => VN_sign_out(9761),
        codeword => codeword(1626),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1627 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9767 downto 9762),
        Din0 => VN1627_in0,
        Din1 => VN1627_in1,
        Din2 => VN1627_in2,
        Din3 => VN1627_in3,
        Din4 => VN1627_in4,
        Din5 => VN1627_in5,
        VN2CN0_bit => VN_data_out(9762),
        VN2CN1_bit => VN_data_out(9763),
        VN2CN2_bit => VN_data_out(9764),
        VN2CN3_bit => VN_data_out(9765),
        VN2CN4_bit => VN_data_out(9766),
        VN2CN5_bit => VN_data_out(9767),
        VN2CN0_sign => VN_sign_out(9762),
        VN2CN1_sign => VN_sign_out(9763),
        VN2CN2_sign => VN_sign_out(9764),
        VN2CN3_sign => VN_sign_out(9765),
        VN2CN4_sign => VN_sign_out(9766),
        VN2CN5_sign => VN_sign_out(9767),
        codeword => codeword(1627),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1628 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9773 downto 9768),
        Din0 => VN1628_in0,
        Din1 => VN1628_in1,
        Din2 => VN1628_in2,
        Din3 => VN1628_in3,
        Din4 => VN1628_in4,
        Din5 => VN1628_in5,
        VN2CN0_bit => VN_data_out(9768),
        VN2CN1_bit => VN_data_out(9769),
        VN2CN2_bit => VN_data_out(9770),
        VN2CN3_bit => VN_data_out(9771),
        VN2CN4_bit => VN_data_out(9772),
        VN2CN5_bit => VN_data_out(9773),
        VN2CN0_sign => VN_sign_out(9768),
        VN2CN1_sign => VN_sign_out(9769),
        VN2CN2_sign => VN_sign_out(9770),
        VN2CN3_sign => VN_sign_out(9771),
        VN2CN4_sign => VN_sign_out(9772),
        VN2CN5_sign => VN_sign_out(9773),
        codeword => codeword(1628),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1629 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9779 downto 9774),
        Din0 => VN1629_in0,
        Din1 => VN1629_in1,
        Din2 => VN1629_in2,
        Din3 => VN1629_in3,
        Din4 => VN1629_in4,
        Din5 => VN1629_in5,
        VN2CN0_bit => VN_data_out(9774),
        VN2CN1_bit => VN_data_out(9775),
        VN2CN2_bit => VN_data_out(9776),
        VN2CN3_bit => VN_data_out(9777),
        VN2CN4_bit => VN_data_out(9778),
        VN2CN5_bit => VN_data_out(9779),
        VN2CN0_sign => VN_sign_out(9774),
        VN2CN1_sign => VN_sign_out(9775),
        VN2CN2_sign => VN_sign_out(9776),
        VN2CN3_sign => VN_sign_out(9777),
        VN2CN4_sign => VN_sign_out(9778),
        VN2CN5_sign => VN_sign_out(9779),
        codeword => codeword(1629),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1630 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9785 downto 9780),
        Din0 => VN1630_in0,
        Din1 => VN1630_in1,
        Din2 => VN1630_in2,
        Din3 => VN1630_in3,
        Din4 => VN1630_in4,
        Din5 => VN1630_in5,
        VN2CN0_bit => VN_data_out(9780),
        VN2CN1_bit => VN_data_out(9781),
        VN2CN2_bit => VN_data_out(9782),
        VN2CN3_bit => VN_data_out(9783),
        VN2CN4_bit => VN_data_out(9784),
        VN2CN5_bit => VN_data_out(9785),
        VN2CN0_sign => VN_sign_out(9780),
        VN2CN1_sign => VN_sign_out(9781),
        VN2CN2_sign => VN_sign_out(9782),
        VN2CN3_sign => VN_sign_out(9783),
        VN2CN4_sign => VN_sign_out(9784),
        VN2CN5_sign => VN_sign_out(9785),
        codeword => codeword(1630),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1631 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9791 downto 9786),
        Din0 => VN1631_in0,
        Din1 => VN1631_in1,
        Din2 => VN1631_in2,
        Din3 => VN1631_in3,
        Din4 => VN1631_in4,
        Din5 => VN1631_in5,
        VN2CN0_bit => VN_data_out(9786),
        VN2CN1_bit => VN_data_out(9787),
        VN2CN2_bit => VN_data_out(9788),
        VN2CN3_bit => VN_data_out(9789),
        VN2CN4_bit => VN_data_out(9790),
        VN2CN5_bit => VN_data_out(9791),
        VN2CN0_sign => VN_sign_out(9786),
        VN2CN1_sign => VN_sign_out(9787),
        VN2CN2_sign => VN_sign_out(9788),
        VN2CN3_sign => VN_sign_out(9789),
        VN2CN4_sign => VN_sign_out(9790),
        VN2CN5_sign => VN_sign_out(9791),
        codeword => codeword(1631),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1632 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9797 downto 9792),
        Din0 => VN1632_in0,
        Din1 => VN1632_in1,
        Din2 => VN1632_in2,
        Din3 => VN1632_in3,
        Din4 => VN1632_in4,
        Din5 => VN1632_in5,
        VN2CN0_bit => VN_data_out(9792),
        VN2CN1_bit => VN_data_out(9793),
        VN2CN2_bit => VN_data_out(9794),
        VN2CN3_bit => VN_data_out(9795),
        VN2CN4_bit => VN_data_out(9796),
        VN2CN5_bit => VN_data_out(9797),
        VN2CN0_sign => VN_sign_out(9792),
        VN2CN1_sign => VN_sign_out(9793),
        VN2CN2_sign => VN_sign_out(9794),
        VN2CN3_sign => VN_sign_out(9795),
        VN2CN4_sign => VN_sign_out(9796),
        VN2CN5_sign => VN_sign_out(9797),
        codeword => codeword(1632),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1633 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9803 downto 9798),
        Din0 => VN1633_in0,
        Din1 => VN1633_in1,
        Din2 => VN1633_in2,
        Din3 => VN1633_in3,
        Din4 => VN1633_in4,
        Din5 => VN1633_in5,
        VN2CN0_bit => VN_data_out(9798),
        VN2CN1_bit => VN_data_out(9799),
        VN2CN2_bit => VN_data_out(9800),
        VN2CN3_bit => VN_data_out(9801),
        VN2CN4_bit => VN_data_out(9802),
        VN2CN5_bit => VN_data_out(9803),
        VN2CN0_sign => VN_sign_out(9798),
        VN2CN1_sign => VN_sign_out(9799),
        VN2CN2_sign => VN_sign_out(9800),
        VN2CN3_sign => VN_sign_out(9801),
        VN2CN4_sign => VN_sign_out(9802),
        VN2CN5_sign => VN_sign_out(9803),
        codeword => codeword(1633),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1634 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9809 downto 9804),
        Din0 => VN1634_in0,
        Din1 => VN1634_in1,
        Din2 => VN1634_in2,
        Din3 => VN1634_in3,
        Din4 => VN1634_in4,
        Din5 => VN1634_in5,
        VN2CN0_bit => VN_data_out(9804),
        VN2CN1_bit => VN_data_out(9805),
        VN2CN2_bit => VN_data_out(9806),
        VN2CN3_bit => VN_data_out(9807),
        VN2CN4_bit => VN_data_out(9808),
        VN2CN5_bit => VN_data_out(9809),
        VN2CN0_sign => VN_sign_out(9804),
        VN2CN1_sign => VN_sign_out(9805),
        VN2CN2_sign => VN_sign_out(9806),
        VN2CN3_sign => VN_sign_out(9807),
        VN2CN4_sign => VN_sign_out(9808),
        VN2CN5_sign => VN_sign_out(9809),
        codeword => codeword(1634),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1635 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9815 downto 9810),
        Din0 => VN1635_in0,
        Din1 => VN1635_in1,
        Din2 => VN1635_in2,
        Din3 => VN1635_in3,
        Din4 => VN1635_in4,
        Din5 => VN1635_in5,
        VN2CN0_bit => VN_data_out(9810),
        VN2CN1_bit => VN_data_out(9811),
        VN2CN2_bit => VN_data_out(9812),
        VN2CN3_bit => VN_data_out(9813),
        VN2CN4_bit => VN_data_out(9814),
        VN2CN5_bit => VN_data_out(9815),
        VN2CN0_sign => VN_sign_out(9810),
        VN2CN1_sign => VN_sign_out(9811),
        VN2CN2_sign => VN_sign_out(9812),
        VN2CN3_sign => VN_sign_out(9813),
        VN2CN4_sign => VN_sign_out(9814),
        VN2CN5_sign => VN_sign_out(9815),
        codeword => codeword(1635),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1636 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9821 downto 9816),
        Din0 => VN1636_in0,
        Din1 => VN1636_in1,
        Din2 => VN1636_in2,
        Din3 => VN1636_in3,
        Din4 => VN1636_in4,
        Din5 => VN1636_in5,
        VN2CN0_bit => VN_data_out(9816),
        VN2CN1_bit => VN_data_out(9817),
        VN2CN2_bit => VN_data_out(9818),
        VN2CN3_bit => VN_data_out(9819),
        VN2CN4_bit => VN_data_out(9820),
        VN2CN5_bit => VN_data_out(9821),
        VN2CN0_sign => VN_sign_out(9816),
        VN2CN1_sign => VN_sign_out(9817),
        VN2CN2_sign => VN_sign_out(9818),
        VN2CN3_sign => VN_sign_out(9819),
        VN2CN4_sign => VN_sign_out(9820),
        VN2CN5_sign => VN_sign_out(9821),
        codeword => codeword(1636),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1637 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9827 downto 9822),
        Din0 => VN1637_in0,
        Din1 => VN1637_in1,
        Din2 => VN1637_in2,
        Din3 => VN1637_in3,
        Din4 => VN1637_in4,
        Din5 => VN1637_in5,
        VN2CN0_bit => VN_data_out(9822),
        VN2CN1_bit => VN_data_out(9823),
        VN2CN2_bit => VN_data_out(9824),
        VN2CN3_bit => VN_data_out(9825),
        VN2CN4_bit => VN_data_out(9826),
        VN2CN5_bit => VN_data_out(9827),
        VN2CN0_sign => VN_sign_out(9822),
        VN2CN1_sign => VN_sign_out(9823),
        VN2CN2_sign => VN_sign_out(9824),
        VN2CN3_sign => VN_sign_out(9825),
        VN2CN4_sign => VN_sign_out(9826),
        VN2CN5_sign => VN_sign_out(9827),
        codeword => codeword(1637),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1638 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9833 downto 9828),
        Din0 => VN1638_in0,
        Din1 => VN1638_in1,
        Din2 => VN1638_in2,
        Din3 => VN1638_in3,
        Din4 => VN1638_in4,
        Din5 => VN1638_in5,
        VN2CN0_bit => VN_data_out(9828),
        VN2CN1_bit => VN_data_out(9829),
        VN2CN2_bit => VN_data_out(9830),
        VN2CN3_bit => VN_data_out(9831),
        VN2CN4_bit => VN_data_out(9832),
        VN2CN5_bit => VN_data_out(9833),
        VN2CN0_sign => VN_sign_out(9828),
        VN2CN1_sign => VN_sign_out(9829),
        VN2CN2_sign => VN_sign_out(9830),
        VN2CN3_sign => VN_sign_out(9831),
        VN2CN4_sign => VN_sign_out(9832),
        VN2CN5_sign => VN_sign_out(9833),
        codeword => codeword(1638),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1639 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9839 downto 9834),
        Din0 => VN1639_in0,
        Din1 => VN1639_in1,
        Din2 => VN1639_in2,
        Din3 => VN1639_in3,
        Din4 => VN1639_in4,
        Din5 => VN1639_in5,
        VN2CN0_bit => VN_data_out(9834),
        VN2CN1_bit => VN_data_out(9835),
        VN2CN2_bit => VN_data_out(9836),
        VN2CN3_bit => VN_data_out(9837),
        VN2CN4_bit => VN_data_out(9838),
        VN2CN5_bit => VN_data_out(9839),
        VN2CN0_sign => VN_sign_out(9834),
        VN2CN1_sign => VN_sign_out(9835),
        VN2CN2_sign => VN_sign_out(9836),
        VN2CN3_sign => VN_sign_out(9837),
        VN2CN4_sign => VN_sign_out(9838),
        VN2CN5_sign => VN_sign_out(9839),
        codeword => codeword(1639),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1640 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9845 downto 9840),
        Din0 => VN1640_in0,
        Din1 => VN1640_in1,
        Din2 => VN1640_in2,
        Din3 => VN1640_in3,
        Din4 => VN1640_in4,
        Din5 => VN1640_in5,
        VN2CN0_bit => VN_data_out(9840),
        VN2CN1_bit => VN_data_out(9841),
        VN2CN2_bit => VN_data_out(9842),
        VN2CN3_bit => VN_data_out(9843),
        VN2CN4_bit => VN_data_out(9844),
        VN2CN5_bit => VN_data_out(9845),
        VN2CN0_sign => VN_sign_out(9840),
        VN2CN1_sign => VN_sign_out(9841),
        VN2CN2_sign => VN_sign_out(9842),
        VN2CN3_sign => VN_sign_out(9843),
        VN2CN4_sign => VN_sign_out(9844),
        VN2CN5_sign => VN_sign_out(9845),
        codeword => codeword(1640),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1641 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9851 downto 9846),
        Din0 => VN1641_in0,
        Din1 => VN1641_in1,
        Din2 => VN1641_in2,
        Din3 => VN1641_in3,
        Din4 => VN1641_in4,
        Din5 => VN1641_in5,
        VN2CN0_bit => VN_data_out(9846),
        VN2CN1_bit => VN_data_out(9847),
        VN2CN2_bit => VN_data_out(9848),
        VN2CN3_bit => VN_data_out(9849),
        VN2CN4_bit => VN_data_out(9850),
        VN2CN5_bit => VN_data_out(9851),
        VN2CN0_sign => VN_sign_out(9846),
        VN2CN1_sign => VN_sign_out(9847),
        VN2CN2_sign => VN_sign_out(9848),
        VN2CN3_sign => VN_sign_out(9849),
        VN2CN4_sign => VN_sign_out(9850),
        VN2CN5_sign => VN_sign_out(9851),
        codeword => codeword(1641),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1642 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9857 downto 9852),
        Din0 => VN1642_in0,
        Din1 => VN1642_in1,
        Din2 => VN1642_in2,
        Din3 => VN1642_in3,
        Din4 => VN1642_in4,
        Din5 => VN1642_in5,
        VN2CN0_bit => VN_data_out(9852),
        VN2CN1_bit => VN_data_out(9853),
        VN2CN2_bit => VN_data_out(9854),
        VN2CN3_bit => VN_data_out(9855),
        VN2CN4_bit => VN_data_out(9856),
        VN2CN5_bit => VN_data_out(9857),
        VN2CN0_sign => VN_sign_out(9852),
        VN2CN1_sign => VN_sign_out(9853),
        VN2CN2_sign => VN_sign_out(9854),
        VN2CN3_sign => VN_sign_out(9855),
        VN2CN4_sign => VN_sign_out(9856),
        VN2CN5_sign => VN_sign_out(9857),
        codeword => codeword(1642),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1643 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9863 downto 9858),
        Din0 => VN1643_in0,
        Din1 => VN1643_in1,
        Din2 => VN1643_in2,
        Din3 => VN1643_in3,
        Din4 => VN1643_in4,
        Din5 => VN1643_in5,
        VN2CN0_bit => VN_data_out(9858),
        VN2CN1_bit => VN_data_out(9859),
        VN2CN2_bit => VN_data_out(9860),
        VN2CN3_bit => VN_data_out(9861),
        VN2CN4_bit => VN_data_out(9862),
        VN2CN5_bit => VN_data_out(9863),
        VN2CN0_sign => VN_sign_out(9858),
        VN2CN1_sign => VN_sign_out(9859),
        VN2CN2_sign => VN_sign_out(9860),
        VN2CN3_sign => VN_sign_out(9861),
        VN2CN4_sign => VN_sign_out(9862),
        VN2CN5_sign => VN_sign_out(9863),
        codeword => codeword(1643),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1644 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9869 downto 9864),
        Din0 => VN1644_in0,
        Din1 => VN1644_in1,
        Din2 => VN1644_in2,
        Din3 => VN1644_in3,
        Din4 => VN1644_in4,
        Din5 => VN1644_in5,
        VN2CN0_bit => VN_data_out(9864),
        VN2CN1_bit => VN_data_out(9865),
        VN2CN2_bit => VN_data_out(9866),
        VN2CN3_bit => VN_data_out(9867),
        VN2CN4_bit => VN_data_out(9868),
        VN2CN5_bit => VN_data_out(9869),
        VN2CN0_sign => VN_sign_out(9864),
        VN2CN1_sign => VN_sign_out(9865),
        VN2CN2_sign => VN_sign_out(9866),
        VN2CN3_sign => VN_sign_out(9867),
        VN2CN4_sign => VN_sign_out(9868),
        VN2CN5_sign => VN_sign_out(9869),
        codeword => codeword(1644),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1645 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9875 downto 9870),
        Din0 => VN1645_in0,
        Din1 => VN1645_in1,
        Din2 => VN1645_in2,
        Din3 => VN1645_in3,
        Din4 => VN1645_in4,
        Din5 => VN1645_in5,
        VN2CN0_bit => VN_data_out(9870),
        VN2CN1_bit => VN_data_out(9871),
        VN2CN2_bit => VN_data_out(9872),
        VN2CN3_bit => VN_data_out(9873),
        VN2CN4_bit => VN_data_out(9874),
        VN2CN5_bit => VN_data_out(9875),
        VN2CN0_sign => VN_sign_out(9870),
        VN2CN1_sign => VN_sign_out(9871),
        VN2CN2_sign => VN_sign_out(9872),
        VN2CN3_sign => VN_sign_out(9873),
        VN2CN4_sign => VN_sign_out(9874),
        VN2CN5_sign => VN_sign_out(9875),
        codeword => codeword(1645),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1646 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9881 downto 9876),
        Din0 => VN1646_in0,
        Din1 => VN1646_in1,
        Din2 => VN1646_in2,
        Din3 => VN1646_in3,
        Din4 => VN1646_in4,
        Din5 => VN1646_in5,
        VN2CN0_bit => VN_data_out(9876),
        VN2CN1_bit => VN_data_out(9877),
        VN2CN2_bit => VN_data_out(9878),
        VN2CN3_bit => VN_data_out(9879),
        VN2CN4_bit => VN_data_out(9880),
        VN2CN5_bit => VN_data_out(9881),
        VN2CN0_sign => VN_sign_out(9876),
        VN2CN1_sign => VN_sign_out(9877),
        VN2CN2_sign => VN_sign_out(9878),
        VN2CN3_sign => VN_sign_out(9879),
        VN2CN4_sign => VN_sign_out(9880),
        VN2CN5_sign => VN_sign_out(9881),
        codeword => codeword(1646),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1647 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9887 downto 9882),
        Din0 => VN1647_in0,
        Din1 => VN1647_in1,
        Din2 => VN1647_in2,
        Din3 => VN1647_in3,
        Din4 => VN1647_in4,
        Din5 => VN1647_in5,
        VN2CN0_bit => VN_data_out(9882),
        VN2CN1_bit => VN_data_out(9883),
        VN2CN2_bit => VN_data_out(9884),
        VN2CN3_bit => VN_data_out(9885),
        VN2CN4_bit => VN_data_out(9886),
        VN2CN5_bit => VN_data_out(9887),
        VN2CN0_sign => VN_sign_out(9882),
        VN2CN1_sign => VN_sign_out(9883),
        VN2CN2_sign => VN_sign_out(9884),
        VN2CN3_sign => VN_sign_out(9885),
        VN2CN4_sign => VN_sign_out(9886),
        VN2CN5_sign => VN_sign_out(9887),
        codeword => codeword(1647),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1648 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9893 downto 9888),
        Din0 => VN1648_in0,
        Din1 => VN1648_in1,
        Din2 => VN1648_in2,
        Din3 => VN1648_in3,
        Din4 => VN1648_in4,
        Din5 => VN1648_in5,
        VN2CN0_bit => VN_data_out(9888),
        VN2CN1_bit => VN_data_out(9889),
        VN2CN2_bit => VN_data_out(9890),
        VN2CN3_bit => VN_data_out(9891),
        VN2CN4_bit => VN_data_out(9892),
        VN2CN5_bit => VN_data_out(9893),
        VN2CN0_sign => VN_sign_out(9888),
        VN2CN1_sign => VN_sign_out(9889),
        VN2CN2_sign => VN_sign_out(9890),
        VN2CN3_sign => VN_sign_out(9891),
        VN2CN4_sign => VN_sign_out(9892),
        VN2CN5_sign => VN_sign_out(9893),
        codeword => codeword(1648),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1649 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9899 downto 9894),
        Din0 => VN1649_in0,
        Din1 => VN1649_in1,
        Din2 => VN1649_in2,
        Din3 => VN1649_in3,
        Din4 => VN1649_in4,
        Din5 => VN1649_in5,
        VN2CN0_bit => VN_data_out(9894),
        VN2CN1_bit => VN_data_out(9895),
        VN2CN2_bit => VN_data_out(9896),
        VN2CN3_bit => VN_data_out(9897),
        VN2CN4_bit => VN_data_out(9898),
        VN2CN5_bit => VN_data_out(9899),
        VN2CN0_sign => VN_sign_out(9894),
        VN2CN1_sign => VN_sign_out(9895),
        VN2CN2_sign => VN_sign_out(9896),
        VN2CN3_sign => VN_sign_out(9897),
        VN2CN4_sign => VN_sign_out(9898),
        VN2CN5_sign => VN_sign_out(9899),
        codeword => codeword(1649),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1650 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9905 downto 9900),
        Din0 => VN1650_in0,
        Din1 => VN1650_in1,
        Din2 => VN1650_in2,
        Din3 => VN1650_in3,
        Din4 => VN1650_in4,
        Din5 => VN1650_in5,
        VN2CN0_bit => VN_data_out(9900),
        VN2CN1_bit => VN_data_out(9901),
        VN2CN2_bit => VN_data_out(9902),
        VN2CN3_bit => VN_data_out(9903),
        VN2CN4_bit => VN_data_out(9904),
        VN2CN5_bit => VN_data_out(9905),
        VN2CN0_sign => VN_sign_out(9900),
        VN2CN1_sign => VN_sign_out(9901),
        VN2CN2_sign => VN_sign_out(9902),
        VN2CN3_sign => VN_sign_out(9903),
        VN2CN4_sign => VN_sign_out(9904),
        VN2CN5_sign => VN_sign_out(9905),
        codeword => codeword(1650),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1651 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9911 downto 9906),
        Din0 => VN1651_in0,
        Din1 => VN1651_in1,
        Din2 => VN1651_in2,
        Din3 => VN1651_in3,
        Din4 => VN1651_in4,
        Din5 => VN1651_in5,
        VN2CN0_bit => VN_data_out(9906),
        VN2CN1_bit => VN_data_out(9907),
        VN2CN2_bit => VN_data_out(9908),
        VN2CN3_bit => VN_data_out(9909),
        VN2CN4_bit => VN_data_out(9910),
        VN2CN5_bit => VN_data_out(9911),
        VN2CN0_sign => VN_sign_out(9906),
        VN2CN1_sign => VN_sign_out(9907),
        VN2CN2_sign => VN_sign_out(9908),
        VN2CN3_sign => VN_sign_out(9909),
        VN2CN4_sign => VN_sign_out(9910),
        VN2CN5_sign => VN_sign_out(9911),
        codeword => codeword(1651),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1652 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9917 downto 9912),
        Din0 => VN1652_in0,
        Din1 => VN1652_in1,
        Din2 => VN1652_in2,
        Din3 => VN1652_in3,
        Din4 => VN1652_in4,
        Din5 => VN1652_in5,
        VN2CN0_bit => VN_data_out(9912),
        VN2CN1_bit => VN_data_out(9913),
        VN2CN2_bit => VN_data_out(9914),
        VN2CN3_bit => VN_data_out(9915),
        VN2CN4_bit => VN_data_out(9916),
        VN2CN5_bit => VN_data_out(9917),
        VN2CN0_sign => VN_sign_out(9912),
        VN2CN1_sign => VN_sign_out(9913),
        VN2CN2_sign => VN_sign_out(9914),
        VN2CN3_sign => VN_sign_out(9915),
        VN2CN4_sign => VN_sign_out(9916),
        VN2CN5_sign => VN_sign_out(9917),
        codeword => codeword(1652),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1653 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9923 downto 9918),
        Din0 => VN1653_in0,
        Din1 => VN1653_in1,
        Din2 => VN1653_in2,
        Din3 => VN1653_in3,
        Din4 => VN1653_in4,
        Din5 => VN1653_in5,
        VN2CN0_bit => VN_data_out(9918),
        VN2CN1_bit => VN_data_out(9919),
        VN2CN2_bit => VN_data_out(9920),
        VN2CN3_bit => VN_data_out(9921),
        VN2CN4_bit => VN_data_out(9922),
        VN2CN5_bit => VN_data_out(9923),
        VN2CN0_sign => VN_sign_out(9918),
        VN2CN1_sign => VN_sign_out(9919),
        VN2CN2_sign => VN_sign_out(9920),
        VN2CN3_sign => VN_sign_out(9921),
        VN2CN4_sign => VN_sign_out(9922),
        VN2CN5_sign => VN_sign_out(9923),
        codeword => codeword(1653),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1654 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9929 downto 9924),
        Din0 => VN1654_in0,
        Din1 => VN1654_in1,
        Din2 => VN1654_in2,
        Din3 => VN1654_in3,
        Din4 => VN1654_in4,
        Din5 => VN1654_in5,
        VN2CN0_bit => VN_data_out(9924),
        VN2CN1_bit => VN_data_out(9925),
        VN2CN2_bit => VN_data_out(9926),
        VN2CN3_bit => VN_data_out(9927),
        VN2CN4_bit => VN_data_out(9928),
        VN2CN5_bit => VN_data_out(9929),
        VN2CN0_sign => VN_sign_out(9924),
        VN2CN1_sign => VN_sign_out(9925),
        VN2CN2_sign => VN_sign_out(9926),
        VN2CN3_sign => VN_sign_out(9927),
        VN2CN4_sign => VN_sign_out(9928),
        VN2CN5_sign => VN_sign_out(9929),
        codeword => codeword(1654),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1655 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9935 downto 9930),
        Din0 => VN1655_in0,
        Din1 => VN1655_in1,
        Din2 => VN1655_in2,
        Din3 => VN1655_in3,
        Din4 => VN1655_in4,
        Din5 => VN1655_in5,
        VN2CN0_bit => VN_data_out(9930),
        VN2CN1_bit => VN_data_out(9931),
        VN2CN2_bit => VN_data_out(9932),
        VN2CN3_bit => VN_data_out(9933),
        VN2CN4_bit => VN_data_out(9934),
        VN2CN5_bit => VN_data_out(9935),
        VN2CN0_sign => VN_sign_out(9930),
        VN2CN1_sign => VN_sign_out(9931),
        VN2CN2_sign => VN_sign_out(9932),
        VN2CN3_sign => VN_sign_out(9933),
        VN2CN4_sign => VN_sign_out(9934),
        VN2CN5_sign => VN_sign_out(9935),
        codeword => codeword(1655),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1656 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9941 downto 9936),
        Din0 => VN1656_in0,
        Din1 => VN1656_in1,
        Din2 => VN1656_in2,
        Din3 => VN1656_in3,
        Din4 => VN1656_in4,
        Din5 => VN1656_in5,
        VN2CN0_bit => VN_data_out(9936),
        VN2CN1_bit => VN_data_out(9937),
        VN2CN2_bit => VN_data_out(9938),
        VN2CN3_bit => VN_data_out(9939),
        VN2CN4_bit => VN_data_out(9940),
        VN2CN5_bit => VN_data_out(9941),
        VN2CN0_sign => VN_sign_out(9936),
        VN2CN1_sign => VN_sign_out(9937),
        VN2CN2_sign => VN_sign_out(9938),
        VN2CN3_sign => VN_sign_out(9939),
        VN2CN4_sign => VN_sign_out(9940),
        VN2CN5_sign => VN_sign_out(9941),
        codeword => codeword(1656),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1657 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9947 downto 9942),
        Din0 => VN1657_in0,
        Din1 => VN1657_in1,
        Din2 => VN1657_in2,
        Din3 => VN1657_in3,
        Din4 => VN1657_in4,
        Din5 => VN1657_in5,
        VN2CN0_bit => VN_data_out(9942),
        VN2CN1_bit => VN_data_out(9943),
        VN2CN2_bit => VN_data_out(9944),
        VN2CN3_bit => VN_data_out(9945),
        VN2CN4_bit => VN_data_out(9946),
        VN2CN5_bit => VN_data_out(9947),
        VN2CN0_sign => VN_sign_out(9942),
        VN2CN1_sign => VN_sign_out(9943),
        VN2CN2_sign => VN_sign_out(9944),
        VN2CN3_sign => VN_sign_out(9945),
        VN2CN4_sign => VN_sign_out(9946),
        VN2CN5_sign => VN_sign_out(9947),
        codeword => codeword(1657),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1658 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9953 downto 9948),
        Din0 => VN1658_in0,
        Din1 => VN1658_in1,
        Din2 => VN1658_in2,
        Din3 => VN1658_in3,
        Din4 => VN1658_in4,
        Din5 => VN1658_in5,
        VN2CN0_bit => VN_data_out(9948),
        VN2CN1_bit => VN_data_out(9949),
        VN2CN2_bit => VN_data_out(9950),
        VN2CN3_bit => VN_data_out(9951),
        VN2CN4_bit => VN_data_out(9952),
        VN2CN5_bit => VN_data_out(9953),
        VN2CN0_sign => VN_sign_out(9948),
        VN2CN1_sign => VN_sign_out(9949),
        VN2CN2_sign => VN_sign_out(9950),
        VN2CN3_sign => VN_sign_out(9951),
        VN2CN4_sign => VN_sign_out(9952),
        VN2CN5_sign => VN_sign_out(9953),
        codeword => codeword(1658),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1659 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9959 downto 9954),
        Din0 => VN1659_in0,
        Din1 => VN1659_in1,
        Din2 => VN1659_in2,
        Din3 => VN1659_in3,
        Din4 => VN1659_in4,
        Din5 => VN1659_in5,
        VN2CN0_bit => VN_data_out(9954),
        VN2CN1_bit => VN_data_out(9955),
        VN2CN2_bit => VN_data_out(9956),
        VN2CN3_bit => VN_data_out(9957),
        VN2CN4_bit => VN_data_out(9958),
        VN2CN5_bit => VN_data_out(9959),
        VN2CN0_sign => VN_sign_out(9954),
        VN2CN1_sign => VN_sign_out(9955),
        VN2CN2_sign => VN_sign_out(9956),
        VN2CN3_sign => VN_sign_out(9957),
        VN2CN4_sign => VN_sign_out(9958),
        VN2CN5_sign => VN_sign_out(9959),
        codeword => codeword(1659),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1660 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9965 downto 9960),
        Din0 => VN1660_in0,
        Din1 => VN1660_in1,
        Din2 => VN1660_in2,
        Din3 => VN1660_in3,
        Din4 => VN1660_in4,
        Din5 => VN1660_in5,
        VN2CN0_bit => VN_data_out(9960),
        VN2CN1_bit => VN_data_out(9961),
        VN2CN2_bit => VN_data_out(9962),
        VN2CN3_bit => VN_data_out(9963),
        VN2CN4_bit => VN_data_out(9964),
        VN2CN5_bit => VN_data_out(9965),
        VN2CN0_sign => VN_sign_out(9960),
        VN2CN1_sign => VN_sign_out(9961),
        VN2CN2_sign => VN_sign_out(9962),
        VN2CN3_sign => VN_sign_out(9963),
        VN2CN4_sign => VN_sign_out(9964),
        VN2CN5_sign => VN_sign_out(9965),
        codeword => codeword(1660),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1661 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9971 downto 9966),
        Din0 => VN1661_in0,
        Din1 => VN1661_in1,
        Din2 => VN1661_in2,
        Din3 => VN1661_in3,
        Din4 => VN1661_in4,
        Din5 => VN1661_in5,
        VN2CN0_bit => VN_data_out(9966),
        VN2CN1_bit => VN_data_out(9967),
        VN2CN2_bit => VN_data_out(9968),
        VN2CN3_bit => VN_data_out(9969),
        VN2CN4_bit => VN_data_out(9970),
        VN2CN5_bit => VN_data_out(9971),
        VN2CN0_sign => VN_sign_out(9966),
        VN2CN1_sign => VN_sign_out(9967),
        VN2CN2_sign => VN_sign_out(9968),
        VN2CN3_sign => VN_sign_out(9969),
        VN2CN4_sign => VN_sign_out(9970),
        VN2CN5_sign => VN_sign_out(9971),
        codeword => codeword(1661),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1662 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9977 downto 9972),
        Din0 => VN1662_in0,
        Din1 => VN1662_in1,
        Din2 => VN1662_in2,
        Din3 => VN1662_in3,
        Din4 => VN1662_in4,
        Din5 => VN1662_in5,
        VN2CN0_bit => VN_data_out(9972),
        VN2CN1_bit => VN_data_out(9973),
        VN2CN2_bit => VN_data_out(9974),
        VN2CN3_bit => VN_data_out(9975),
        VN2CN4_bit => VN_data_out(9976),
        VN2CN5_bit => VN_data_out(9977),
        VN2CN0_sign => VN_sign_out(9972),
        VN2CN1_sign => VN_sign_out(9973),
        VN2CN2_sign => VN_sign_out(9974),
        VN2CN3_sign => VN_sign_out(9975),
        VN2CN4_sign => VN_sign_out(9976),
        VN2CN5_sign => VN_sign_out(9977),
        codeword => codeword(1662),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1663 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9983 downto 9978),
        Din0 => VN1663_in0,
        Din1 => VN1663_in1,
        Din2 => VN1663_in2,
        Din3 => VN1663_in3,
        Din4 => VN1663_in4,
        Din5 => VN1663_in5,
        VN2CN0_bit => VN_data_out(9978),
        VN2CN1_bit => VN_data_out(9979),
        VN2CN2_bit => VN_data_out(9980),
        VN2CN3_bit => VN_data_out(9981),
        VN2CN4_bit => VN_data_out(9982),
        VN2CN5_bit => VN_data_out(9983),
        VN2CN0_sign => VN_sign_out(9978),
        VN2CN1_sign => VN_sign_out(9979),
        VN2CN2_sign => VN_sign_out(9980),
        VN2CN3_sign => VN_sign_out(9981),
        VN2CN4_sign => VN_sign_out(9982),
        VN2CN5_sign => VN_sign_out(9983),
        codeword => codeword(1663),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1664 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9989 downto 9984),
        Din0 => VN1664_in0,
        Din1 => VN1664_in1,
        Din2 => VN1664_in2,
        Din3 => VN1664_in3,
        Din4 => VN1664_in4,
        Din5 => VN1664_in5,
        VN2CN0_bit => VN_data_out(9984),
        VN2CN1_bit => VN_data_out(9985),
        VN2CN2_bit => VN_data_out(9986),
        VN2CN3_bit => VN_data_out(9987),
        VN2CN4_bit => VN_data_out(9988),
        VN2CN5_bit => VN_data_out(9989),
        VN2CN0_sign => VN_sign_out(9984),
        VN2CN1_sign => VN_sign_out(9985),
        VN2CN2_sign => VN_sign_out(9986),
        VN2CN3_sign => VN_sign_out(9987),
        VN2CN4_sign => VN_sign_out(9988),
        VN2CN5_sign => VN_sign_out(9989),
        codeword => codeword(1664),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1665 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(9995 downto 9990),
        Din0 => VN1665_in0,
        Din1 => VN1665_in1,
        Din2 => VN1665_in2,
        Din3 => VN1665_in3,
        Din4 => VN1665_in4,
        Din5 => VN1665_in5,
        VN2CN0_bit => VN_data_out(9990),
        VN2CN1_bit => VN_data_out(9991),
        VN2CN2_bit => VN_data_out(9992),
        VN2CN3_bit => VN_data_out(9993),
        VN2CN4_bit => VN_data_out(9994),
        VN2CN5_bit => VN_data_out(9995),
        VN2CN0_sign => VN_sign_out(9990),
        VN2CN1_sign => VN_sign_out(9991),
        VN2CN2_sign => VN_sign_out(9992),
        VN2CN3_sign => VN_sign_out(9993),
        VN2CN4_sign => VN_sign_out(9994),
        VN2CN5_sign => VN_sign_out(9995),
        codeword => codeword(1665),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1666 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10001 downto 9996),
        Din0 => VN1666_in0,
        Din1 => VN1666_in1,
        Din2 => VN1666_in2,
        Din3 => VN1666_in3,
        Din4 => VN1666_in4,
        Din5 => VN1666_in5,
        VN2CN0_bit => VN_data_out(9996),
        VN2CN1_bit => VN_data_out(9997),
        VN2CN2_bit => VN_data_out(9998),
        VN2CN3_bit => VN_data_out(9999),
        VN2CN4_bit => VN_data_out(10000),
        VN2CN5_bit => VN_data_out(10001),
        VN2CN0_sign => VN_sign_out(9996),
        VN2CN1_sign => VN_sign_out(9997),
        VN2CN2_sign => VN_sign_out(9998),
        VN2CN3_sign => VN_sign_out(9999),
        VN2CN4_sign => VN_sign_out(10000),
        VN2CN5_sign => VN_sign_out(10001),
        codeword => codeword(1666),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1667 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10007 downto 10002),
        Din0 => VN1667_in0,
        Din1 => VN1667_in1,
        Din2 => VN1667_in2,
        Din3 => VN1667_in3,
        Din4 => VN1667_in4,
        Din5 => VN1667_in5,
        VN2CN0_bit => VN_data_out(10002),
        VN2CN1_bit => VN_data_out(10003),
        VN2CN2_bit => VN_data_out(10004),
        VN2CN3_bit => VN_data_out(10005),
        VN2CN4_bit => VN_data_out(10006),
        VN2CN5_bit => VN_data_out(10007),
        VN2CN0_sign => VN_sign_out(10002),
        VN2CN1_sign => VN_sign_out(10003),
        VN2CN2_sign => VN_sign_out(10004),
        VN2CN3_sign => VN_sign_out(10005),
        VN2CN4_sign => VN_sign_out(10006),
        VN2CN5_sign => VN_sign_out(10007),
        codeword => codeword(1667),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1668 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10013 downto 10008),
        Din0 => VN1668_in0,
        Din1 => VN1668_in1,
        Din2 => VN1668_in2,
        Din3 => VN1668_in3,
        Din4 => VN1668_in4,
        Din5 => VN1668_in5,
        VN2CN0_bit => VN_data_out(10008),
        VN2CN1_bit => VN_data_out(10009),
        VN2CN2_bit => VN_data_out(10010),
        VN2CN3_bit => VN_data_out(10011),
        VN2CN4_bit => VN_data_out(10012),
        VN2CN5_bit => VN_data_out(10013),
        VN2CN0_sign => VN_sign_out(10008),
        VN2CN1_sign => VN_sign_out(10009),
        VN2CN2_sign => VN_sign_out(10010),
        VN2CN3_sign => VN_sign_out(10011),
        VN2CN4_sign => VN_sign_out(10012),
        VN2CN5_sign => VN_sign_out(10013),
        codeword => codeword(1668),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1669 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10019 downto 10014),
        Din0 => VN1669_in0,
        Din1 => VN1669_in1,
        Din2 => VN1669_in2,
        Din3 => VN1669_in3,
        Din4 => VN1669_in4,
        Din5 => VN1669_in5,
        VN2CN0_bit => VN_data_out(10014),
        VN2CN1_bit => VN_data_out(10015),
        VN2CN2_bit => VN_data_out(10016),
        VN2CN3_bit => VN_data_out(10017),
        VN2CN4_bit => VN_data_out(10018),
        VN2CN5_bit => VN_data_out(10019),
        VN2CN0_sign => VN_sign_out(10014),
        VN2CN1_sign => VN_sign_out(10015),
        VN2CN2_sign => VN_sign_out(10016),
        VN2CN3_sign => VN_sign_out(10017),
        VN2CN4_sign => VN_sign_out(10018),
        VN2CN5_sign => VN_sign_out(10019),
        codeword => codeword(1669),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1670 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10025 downto 10020),
        Din0 => VN1670_in0,
        Din1 => VN1670_in1,
        Din2 => VN1670_in2,
        Din3 => VN1670_in3,
        Din4 => VN1670_in4,
        Din5 => VN1670_in5,
        VN2CN0_bit => VN_data_out(10020),
        VN2CN1_bit => VN_data_out(10021),
        VN2CN2_bit => VN_data_out(10022),
        VN2CN3_bit => VN_data_out(10023),
        VN2CN4_bit => VN_data_out(10024),
        VN2CN5_bit => VN_data_out(10025),
        VN2CN0_sign => VN_sign_out(10020),
        VN2CN1_sign => VN_sign_out(10021),
        VN2CN2_sign => VN_sign_out(10022),
        VN2CN3_sign => VN_sign_out(10023),
        VN2CN4_sign => VN_sign_out(10024),
        VN2CN5_sign => VN_sign_out(10025),
        codeword => codeword(1670),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1671 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10031 downto 10026),
        Din0 => VN1671_in0,
        Din1 => VN1671_in1,
        Din2 => VN1671_in2,
        Din3 => VN1671_in3,
        Din4 => VN1671_in4,
        Din5 => VN1671_in5,
        VN2CN0_bit => VN_data_out(10026),
        VN2CN1_bit => VN_data_out(10027),
        VN2CN2_bit => VN_data_out(10028),
        VN2CN3_bit => VN_data_out(10029),
        VN2CN4_bit => VN_data_out(10030),
        VN2CN5_bit => VN_data_out(10031),
        VN2CN0_sign => VN_sign_out(10026),
        VN2CN1_sign => VN_sign_out(10027),
        VN2CN2_sign => VN_sign_out(10028),
        VN2CN3_sign => VN_sign_out(10029),
        VN2CN4_sign => VN_sign_out(10030),
        VN2CN5_sign => VN_sign_out(10031),
        codeword => codeword(1671),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1672 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10037 downto 10032),
        Din0 => VN1672_in0,
        Din1 => VN1672_in1,
        Din2 => VN1672_in2,
        Din3 => VN1672_in3,
        Din4 => VN1672_in4,
        Din5 => VN1672_in5,
        VN2CN0_bit => VN_data_out(10032),
        VN2CN1_bit => VN_data_out(10033),
        VN2CN2_bit => VN_data_out(10034),
        VN2CN3_bit => VN_data_out(10035),
        VN2CN4_bit => VN_data_out(10036),
        VN2CN5_bit => VN_data_out(10037),
        VN2CN0_sign => VN_sign_out(10032),
        VN2CN1_sign => VN_sign_out(10033),
        VN2CN2_sign => VN_sign_out(10034),
        VN2CN3_sign => VN_sign_out(10035),
        VN2CN4_sign => VN_sign_out(10036),
        VN2CN5_sign => VN_sign_out(10037),
        codeword => codeword(1672),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1673 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10043 downto 10038),
        Din0 => VN1673_in0,
        Din1 => VN1673_in1,
        Din2 => VN1673_in2,
        Din3 => VN1673_in3,
        Din4 => VN1673_in4,
        Din5 => VN1673_in5,
        VN2CN0_bit => VN_data_out(10038),
        VN2CN1_bit => VN_data_out(10039),
        VN2CN2_bit => VN_data_out(10040),
        VN2CN3_bit => VN_data_out(10041),
        VN2CN4_bit => VN_data_out(10042),
        VN2CN5_bit => VN_data_out(10043),
        VN2CN0_sign => VN_sign_out(10038),
        VN2CN1_sign => VN_sign_out(10039),
        VN2CN2_sign => VN_sign_out(10040),
        VN2CN3_sign => VN_sign_out(10041),
        VN2CN4_sign => VN_sign_out(10042),
        VN2CN5_sign => VN_sign_out(10043),
        codeword => codeword(1673),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1674 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10049 downto 10044),
        Din0 => VN1674_in0,
        Din1 => VN1674_in1,
        Din2 => VN1674_in2,
        Din3 => VN1674_in3,
        Din4 => VN1674_in4,
        Din5 => VN1674_in5,
        VN2CN0_bit => VN_data_out(10044),
        VN2CN1_bit => VN_data_out(10045),
        VN2CN2_bit => VN_data_out(10046),
        VN2CN3_bit => VN_data_out(10047),
        VN2CN4_bit => VN_data_out(10048),
        VN2CN5_bit => VN_data_out(10049),
        VN2CN0_sign => VN_sign_out(10044),
        VN2CN1_sign => VN_sign_out(10045),
        VN2CN2_sign => VN_sign_out(10046),
        VN2CN3_sign => VN_sign_out(10047),
        VN2CN4_sign => VN_sign_out(10048),
        VN2CN5_sign => VN_sign_out(10049),
        codeword => codeword(1674),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1675 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10055 downto 10050),
        Din0 => VN1675_in0,
        Din1 => VN1675_in1,
        Din2 => VN1675_in2,
        Din3 => VN1675_in3,
        Din4 => VN1675_in4,
        Din5 => VN1675_in5,
        VN2CN0_bit => VN_data_out(10050),
        VN2CN1_bit => VN_data_out(10051),
        VN2CN2_bit => VN_data_out(10052),
        VN2CN3_bit => VN_data_out(10053),
        VN2CN4_bit => VN_data_out(10054),
        VN2CN5_bit => VN_data_out(10055),
        VN2CN0_sign => VN_sign_out(10050),
        VN2CN1_sign => VN_sign_out(10051),
        VN2CN2_sign => VN_sign_out(10052),
        VN2CN3_sign => VN_sign_out(10053),
        VN2CN4_sign => VN_sign_out(10054),
        VN2CN5_sign => VN_sign_out(10055),
        codeword => codeword(1675),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1676 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10061 downto 10056),
        Din0 => VN1676_in0,
        Din1 => VN1676_in1,
        Din2 => VN1676_in2,
        Din3 => VN1676_in3,
        Din4 => VN1676_in4,
        Din5 => VN1676_in5,
        VN2CN0_bit => VN_data_out(10056),
        VN2CN1_bit => VN_data_out(10057),
        VN2CN2_bit => VN_data_out(10058),
        VN2CN3_bit => VN_data_out(10059),
        VN2CN4_bit => VN_data_out(10060),
        VN2CN5_bit => VN_data_out(10061),
        VN2CN0_sign => VN_sign_out(10056),
        VN2CN1_sign => VN_sign_out(10057),
        VN2CN2_sign => VN_sign_out(10058),
        VN2CN3_sign => VN_sign_out(10059),
        VN2CN4_sign => VN_sign_out(10060),
        VN2CN5_sign => VN_sign_out(10061),
        codeword => codeword(1676),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1677 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10067 downto 10062),
        Din0 => VN1677_in0,
        Din1 => VN1677_in1,
        Din2 => VN1677_in2,
        Din3 => VN1677_in3,
        Din4 => VN1677_in4,
        Din5 => VN1677_in5,
        VN2CN0_bit => VN_data_out(10062),
        VN2CN1_bit => VN_data_out(10063),
        VN2CN2_bit => VN_data_out(10064),
        VN2CN3_bit => VN_data_out(10065),
        VN2CN4_bit => VN_data_out(10066),
        VN2CN5_bit => VN_data_out(10067),
        VN2CN0_sign => VN_sign_out(10062),
        VN2CN1_sign => VN_sign_out(10063),
        VN2CN2_sign => VN_sign_out(10064),
        VN2CN3_sign => VN_sign_out(10065),
        VN2CN4_sign => VN_sign_out(10066),
        VN2CN5_sign => VN_sign_out(10067),
        codeword => codeword(1677),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1678 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10073 downto 10068),
        Din0 => VN1678_in0,
        Din1 => VN1678_in1,
        Din2 => VN1678_in2,
        Din3 => VN1678_in3,
        Din4 => VN1678_in4,
        Din5 => VN1678_in5,
        VN2CN0_bit => VN_data_out(10068),
        VN2CN1_bit => VN_data_out(10069),
        VN2CN2_bit => VN_data_out(10070),
        VN2CN3_bit => VN_data_out(10071),
        VN2CN4_bit => VN_data_out(10072),
        VN2CN5_bit => VN_data_out(10073),
        VN2CN0_sign => VN_sign_out(10068),
        VN2CN1_sign => VN_sign_out(10069),
        VN2CN2_sign => VN_sign_out(10070),
        VN2CN3_sign => VN_sign_out(10071),
        VN2CN4_sign => VN_sign_out(10072),
        VN2CN5_sign => VN_sign_out(10073),
        codeword => codeword(1678),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1679 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10079 downto 10074),
        Din0 => VN1679_in0,
        Din1 => VN1679_in1,
        Din2 => VN1679_in2,
        Din3 => VN1679_in3,
        Din4 => VN1679_in4,
        Din5 => VN1679_in5,
        VN2CN0_bit => VN_data_out(10074),
        VN2CN1_bit => VN_data_out(10075),
        VN2CN2_bit => VN_data_out(10076),
        VN2CN3_bit => VN_data_out(10077),
        VN2CN4_bit => VN_data_out(10078),
        VN2CN5_bit => VN_data_out(10079),
        VN2CN0_sign => VN_sign_out(10074),
        VN2CN1_sign => VN_sign_out(10075),
        VN2CN2_sign => VN_sign_out(10076),
        VN2CN3_sign => VN_sign_out(10077),
        VN2CN4_sign => VN_sign_out(10078),
        VN2CN5_sign => VN_sign_out(10079),
        codeword => codeword(1679),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1680 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10085 downto 10080),
        Din0 => VN1680_in0,
        Din1 => VN1680_in1,
        Din2 => VN1680_in2,
        Din3 => VN1680_in3,
        Din4 => VN1680_in4,
        Din5 => VN1680_in5,
        VN2CN0_bit => VN_data_out(10080),
        VN2CN1_bit => VN_data_out(10081),
        VN2CN2_bit => VN_data_out(10082),
        VN2CN3_bit => VN_data_out(10083),
        VN2CN4_bit => VN_data_out(10084),
        VN2CN5_bit => VN_data_out(10085),
        VN2CN0_sign => VN_sign_out(10080),
        VN2CN1_sign => VN_sign_out(10081),
        VN2CN2_sign => VN_sign_out(10082),
        VN2CN3_sign => VN_sign_out(10083),
        VN2CN4_sign => VN_sign_out(10084),
        VN2CN5_sign => VN_sign_out(10085),
        codeword => codeword(1680),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1681 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10091 downto 10086),
        Din0 => VN1681_in0,
        Din1 => VN1681_in1,
        Din2 => VN1681_in2,
        Din3 => VN1681_in3,
        Din4 => VN1681_in4,
        Din5 => VN1681_in5,
        VN2CN0_bit => VN_data_out(10086),
        VN2CN1_bit => VN_data_out(10087),
        VN2CN2_bit => VN_data_out(10088),
        VN2CN3_bit => VN_data_out(10089),
        VN2CN4_bit => VN_data_out(10090),
        VN2CN5_bit => VN_data_out(10091),
        VN2CN0_sign => VN_sign_out(10086),
        VN2CN1_sign => VN_sign_out(10087),
        VN2CN2_sign => VN_sign_out(10088),
        VN2CN3_sign => VN_sign_out(10089),
        VN2CN4_sign => VN_sign_out(10090),
        VN2CN5_sign => VN_sign_out(10091),
        codeword => codeword(1681),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1682 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10097 downto 10092),
        Din0 => VN1682_in0,
        Din1 => VN1682_in1,
        Din2 => VN1682_in2,
        Din3 => VN1682_in3,
        Din4 => VN1682_in4,
        Din5 => VN1682_in5,
        VN2CN0_bit => VN_data_out(10092),
        VN2CN1_bit => VN_data_out(10093),
        VN2CN2_bit => VN_data_out(10094),
        VN2CN3_bit => VN_data_out(10095),
        VN2CN4_bit => VN_data_out(10096),
        VN2CN5_bit => VN_data_out(10097),
        VN2CN0_sign => VN_sign_out(10092),
        VN2CN1_sign => VN_sign_out(10093),
        VN2CN2_sign => VN_sign_out(10094),
        VN2CN3_sign => VN_sign_out(10095),
        VN2CN4_sign => VN_sign_out(10096),
        VN2CN5_sign => VN_sign_out(10097),
        codeword => codeword(1682),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1683 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10103 downto 10098),
        Din0 => VN1683_in0,
        Din1 => VN1683_in1,
        Din2 => VN1683_in2,
        Din3 => VN1683_in3,
        Din4 => VN1683_in4,
        Din5 => VN1683_in5,
        VN2CN0_bit => VN_data_out(10098),
        VN2CN1_bit => VN_data_out(10099),
        VN2CN2_bit => VN_data_out(10100),
        VN2CN3_bit => VN_data_out(10101),
        VN2CN4_bit => VN_data_out(10102),
        VN2CN5_bit => VN_data_out(10103),
        VN2CN0_sign => VN_sign_out(10098),
        VN2CN1_sign => VN_sign_out(10099),
        VN2CN2_sign => VN_sign_out(10100),
        VN2CN3_sign => VN_sign_out(10101),
        VN2CN4_sign => VN_sign_out(10102),
        VN2CN5_sign => VN_sign_out(10103),
        codeword => codeword(1683),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1684 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10109 downto 10104),
        Din0 => VN1684_in0,
        Din1 => VN1684_in1,
        Din2 => VN1684_in2,
        Din3 => VN1684_in3,
        Din4 => VN1684_in4,
        Din5 => VN1684_in5,
        VN2CN0_bit => VN_data_out(10104),
        VN2CN1_bit => VN_data_out(10105),
        VN2CN2_bit => VN_data_out(10106),
        VN2CN3_bit => VN_data_out(10107),
        VN2CN4_bit => VN_data_out(10108),
        VN2CN5_bit => VN_data_out(10109),
        VN2CN0_sign => VN_sign_out(10104),
        VN2CN1_sign => VN_sign_out(10105),
        VN2CN2_sign => VN_sign_out(10106),
        VN2CN3_sign => VN_sign_out(10107),
        VN2CN4_sign => VN_sign_out(10108),
        VN2CN5_sign => VN_sign_out(10109),
        codeword => codeword(1684),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1685 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10115 downto 10110),
        Din0 => VN1685_in0,
        Din1 => VN1685_in1,
        Din2 => VN1685_in2,
        Din3 => VN1685_in3,
        Din4 => VN1685_in4,
        Din5 => VN1685_in5,
        VN2CN0_bit => VN_data_out(10110),
        VN2CN1_bit => VN_data_out(10111),
        VN2CN2_bit => VN_data_out(10112),
        VN2CN3_bit => VN_data_out(10113),
        VN2CN4_bit => VN_data_out(10114),
        VN2CN5_bit => VN_data_out(10115),
        VN2CN0_sign => VN_sign_out(10110),
        VN2CN1_sign => VN_sign_out(10111),
        VN2CN2_sign => VN_sign_out(10112),
        VN2CN3_sign => VN_sign_out(10113),
        VN2CN4_sign => VN_sign_out(10114),
        VN2CN5_sign => VN_sign_out(10115),
        codeword => codeword(1685),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1686 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10121 downto 10116),
        Din0 => VN1686_in0,
        Din1 => VN1686_in1,
        Din2 => VN1686_in2,
        Din3 => VN1686_in3,
        Din4 => VN1686_in4,
        Din5 => VN1686_in5,
        VN2CN0_bit => VN_data_out(10116),
        VN2CN1_bit => VN_data_out(10117),
        VN2CN2_bit => VN_data_out(10118),
        VN2CN3_bit => VN_data_out(10119),
        VN2CN4_bit => VN_data_out(10120),
        VN2CN5_bit => VN_data_out(10121),
        VN2CN0_sign => VN_sign_out(10116),
        VN2CN1_sign => VN_sign_out(10117),
        VN2CN2_sign => VN_sign_out(10118),
        VN2CN3_sign => VN_sign_out(10119),
        VN2CN4_sign => VN_sign_out(10120),
        VN2CN5_sign => VN_sign_out(10121),
        codeword => codeword(1686),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1687 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10127 downto 10122),
        Din0 => VN1687_in0,
        Din1 => VN1687_in1,
        Din2 => VN1687_in2,
        Din3 => VN1687_in3,
        Din4 => VN1687_in4,
        Din5 => VN1687_in5,
        VN2CN0_bit => VN_data_out(10122),
        VN2CN1_bit => VN_data_out(10123),
        VN2CN2_bit => VN_data_out(10124),
        VN2CN3_bit => VN_data_out(10125),
        VN2CN4_bit => VN_data_out(10126),
        VN2CN5_bit => VN_data_out(10127),
        VN2CN0_sign => VN_sign_out(10122),
        VN2CN1_sign => VN_sign_out(10123),
        VN2CN2_sign => VN_sign_out(10124),
        VN2CN3_sign => VN_sign_out(10125),
        VN2CN4_sign => VN_sign_out(10126),
        VN2CN5_sign => VN_sign_out(10127),
        codeword => codeword(1687),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1688 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10133 downto 10128),
        Din0 => VN1688_in0,
        Din1 => VN1688_in1,
        Din2 => VN1688_in2,
        Din3 => VN1688_in3,
        Din4 => VN1688_in4,
        Din5 => VN1688_in5,
        VN2CN0_bit => VN_data_out(10128),
        VN2CN1_bit => VN_data_out(10129),
        VN2CN2_bit => VN_data_out(10130),
        VN2CN3_bit => VN_data_out(10131),
        VN2CN4_bit => VN_data_out(10132),
        VN2CN5_bit => VN_data_out(10133),
        VN2CN0_sign => VN_sign_out(10128),
        VN2CN1_sign => VN_sign_out(10129),
        VN2CN2_sign => VN_sign_out(10130),
        VN2CN3_sign => VN_sign_out(10131),
        VN2CN4_sign => VN_sign_out(10132),
        VN2CN5_sign => VN_sign_out(10133),
        codeword => codeword(1688),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1689 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10139 downto 10134),
        Din0 => VN1689_in0,
        Din1 => VN1689_in1,
        Din2 => VN1689_in2,
        Din3 => VN1689_in3,
        Din4 => VN1689_in4,
        Din5 => VN1689_in5,
        VN2CN0_bit => VN_data_out(10134),
        VN2CN1_bit => VN_data_out(10135),
        VN2CN2_bit => VN_data_out(10136),
        VN2CN3_bit => VN_data_out(10137),
        VN2CN4_bit => VN_data_out(10138),
        VN2CN5_bit => VN_data_out(10139),
        VN2CN0_sign => VN_sign_out(10134),
        VN2CN1_sign => VN_sign_out(10135),
        VN2CN2_sign => VN_sign_out(10136),
        VN2CN3_sign => VN_sign_out(10137),
        VN2CN4_sign => VN_sign_out(10138),
        VN2CN5_sign => VN_sign_out(10139),
        codeword => codeword(1689),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1690 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10145 downto 10140),
        Din0 => VN1690_in0,
        Din1 => VN1690_in1,
        Din2 => VN1690_in2,
        Din3 => VN1690_in3,
        Din4 => VN1690_in4,
        Din5 => VN1690_in5,
        VN2CN0_bit => VN_data_out(10140),
        VN2CN1_bit => VN_data_out(10141),
        VN2CN2_bit => VN_data_out(10142),
        VN2CN3_bit => VN_data_out(10143),
        VN2CN4_bit => VN_data_out(10144),
        VN2CN5_bit => VN_data_out(10145),
        VN2CN0_sign => VN_sign_out(10140),
        VN2CN1_sign => VN_sign_out(10141),
        VN2CN2_sign => VN_sign_out(10142),
        VN2CN3_sign => VN_sign_out(10143),
        VN2CN4_sign => VN_sign_out(10144),
        VN2CN5_sign => VN_sign_out(10145),
        codeword => codeword(1690),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1691 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10151 downto 10146),
        Din0 => VN1691_in0,
        Din1 => VN1691_in1,
        Din2 => VN1691_in2,
        Din3 => VN1691_in3,
        Din4 => VN1691_in4,
        Din5 => VN1691_in5,
        VN2CN0_bit => VN_data_out(10146),
        VN2CN1_bit => VN_data_out(10147),
        VN2CN2_bit => VN_data_out(10148),
        VN2CN3_bit => VN_data_out(10149),
        VN2CN4_bit => VN_data_out(10150),
        VN2CN5_bit => VN_data_out(10151),
        VN2CN0_sign => VN_sign_out(10146),
        VN2CN1_sign => VN_sign_out(10147),
        VN2CN2_sign => VN_sign_out(10148),
        VN2CN3_sign => VN_sign_out(10149),
        VN2CN4_sign => VN_sign_out(10150),
        VN2CN5_sign => VN_sign_out(10151),
        codeword => codeword(1691),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1692 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10157 downto 10152),
        Din0 => VN1692_in0,
        Din1 => VN1692_in1,
        Din2 => VN1692_in2,
        Din3 => VN1692_in3,
        Din4 => VN1692_in4,
        Din5 => VN1692_in5,
        VN2CN0_bit => VN_data_out(10152),
        VN2CN1_bit => VN_data_out(10153),
        VN2CN2_bit => VN_data_out(10154),
        VN2CN3_bit => VN_data_out(10155),
        VN2CN4_bit => VN_data_out(10156),
        VN2CN5_bit => VN_data_out(10157),
        VN2CN0_sign => VN_sign_out(10152),
        VN2CN1_sign => VN_sign_out(10153),
        VN2CN2_sign => VN_sign_out(10154),
        VN2CN3_sign => VN_sign_out(10155),
        VN2CN4_sign => VN_sign_out(10156),
        VN2CN5_sign => VN_sign_out(10157),
        codeword => codeword(1692),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1693 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10163 downto 10158),
        Din0 => VN1693_in0,
        Din1 => VN1693_in1,
        Din2 => VN1693_in2,
        Din3 => VN1693_in3,
        Din4 => VN1693_in4,
        Din5 => VN1693_in5,
        VN2CN0_bit => VN_data_out(10158),
        VN2CN1_bit => VN_data_out(10159),
        VN2CN2_bit => VN_data_out(10160),
        VN2CN3_bit => VN_data_out(10161),
        VN2CN4_bit => VN_data_out(10162),
        VN2CN5_bit => VN_data_out(10163),
        VN2CN0_sign => VN_sign_out(10158),
        VN2CN1_sign => VN_sign_out(10159),
        VN2CN2_sign => VN_sign_out(10160),
        VN2CN3_sign => VN_sign_out(10161),
        VN2CN4_sign => VN_sign_out(10162),
        VN2CN5_sign => VN_sign_out(10163),
        codeword => codeword(1693),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1694 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10169 downto 10164),
        Din0 => VN1694_in0,
        Din1 => VN1694_in1,
        Din2 => VN1694_in2,
        Din3 => VN1694_in3,
        Din4 => VN1694_in4,
        Din5 => VN1694_in5,
        VN2CN0_bit => VN_data_out(10164),
        VN2CN1_bit => VN_data_out(10165),
        VN2CN2_bit => VN_data_out(10166),
        VN2CN3_bit => VN_data_out(10167),
        VN2CN4_bit => VN_data_out(10168),
        VN2CN5_bit => VN_data_out(10169),
        VN2CN0_sign => VN_sign_out(10164),
        VN2CN1_sign => VN_sign_out(10165),
        VN2CN2_sign => VN_sign_out(10166),
        VN2CN3_sign => VN_sign_out(10167),
        VN2CN4_sign => VN_sign_out(10168),
        VN2CN5_sign => VN_sign_out(10169),
        codeword => codeword(1694),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1695 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10175 downto 10170),
        Din0 => VN1695_in0,
        Din1 => VN1695_in1,
        Din2 => VN1695_in2,
        Din3 => VN1695_in3,
        Din4 => VN1695_in4,
        Din5 => VN1695_in5,
        VN2CN0_bit => VN_data_out(10170),
        VN2CN1_bit => VN_data_out(10171),
        VN2CN2_bit => VN_data_out(10172),
        VN2CN3_bit => VN_data_out(10173),
        VN2CN4_bit => VN_data_out(10174),
        VN2CN5_bit => VN_data_out(10175),
        VN2CN0_sign => VN_sign_out(10170),
        VN2CN1_sign => VN_sign_out(10171),
        VN2CN2_sign => VN_sign_out(10172),
        VN2CN3_sign => VN_sign_out(10173),
        VN2CN4_sign => VN_sign_out(10174),
        VN2CN5_sign => VN_sign_out(10175),
        codeword => codeword(1695),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1696 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10181 downto 10176),
        Din0 => VN1696_in0,
        Din1 => VN1696_in1,
        Din2 => VN1696_in2,
        Din3 => VN1696_in3,
        Din4 => VN1696_in4,
        Din5 => VN1696_in5,
        VN2CN0_bit => VN_data_out(10176),
        VN2CN1_bit => VN_data_out(10177),
        VN2CN2_bit => VN_data_out(10178),
        VN2CN3_bit => VN_data_out(10179),
        VN2CN4_bit => VN_data_out(10180),
        VN2CN5_bit => VN_data_out(10181),
        VN2CN0_sign => VN_sign_out(10176),
        VN2CN1_sign => VN_sign_out(10177),
        VN2CN2_sign => VN_sign_out(10178),
        VN2CN3_sign => VN_sign_out(10179),
        VN2CN4_sign => VN_sign_out(10180),
        VN2CN5_sign => VN_sign_out(10181),
        codeword => codeword(1696),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1697 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10187 downto 10182),
        Din0 => VN1697_in0,
        Din1 => VN1697_in1,
        Din2 => VN1697_in2,
        Din3 => VN1697_in3,
        Din4 => VN1697_in4,
        Din5 => VN1697_in5,
        VN2CN0_bit => VN_data_out(10182),
        VN2CN1_bit => VN_data_out(10183),
        VN2CN2_bit => VN_data_out(10184),
        VN2CN3_bit => VN_data_out(10185),
        VN2CN4_bit => VN_data_out(10186),
        VN2CN5_bit => VN_data_out(10187),
        VN2CN0_sign => VN_sign_out(10182),
        VN2CN1_sign => VN_sign_out(10183),
        VN2CN2_sign => VN_sign_out(10184),
        VN2CN3_sign => VN_sign_out(10185),
        VN2CN4_sign => VN_sign_out(10186),
        VN2CN5_sign => VN_sign_out(10187),
        codeword => codeword(1697),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1698 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10193 downto 10188),
        Din0 => VN1698_in0,
        Din1 => VN1698_in1,
        Din2 => VN1698_in2,
        Din3 => VN1698_in3,
        Din4 => VN1698_in4,
        Din5 => VN1698_in5,
        VN2CN0_bit => VN_data_out(10188),
        VN2CN1_bit => VN_data_out(10189),
        VN2CN2_bit => VN_data_out(10190),
        VN2CN3_bit => VN_data_out(10191),
        VN2CN4_bit => VN_data_out(10192),
        VN2CN5_bit => VN_data_out(10193),
        VN2CN0_sign => VN_sign_out(10188),
        VN2CN1_sign => VN_sign_out(10189),
        VN2CN2_sign => VN_sign_out(10190),
        VN2CN3_sign => VN_sign_out(10191),
        VN2CN4_sign => VN_sign_out(10192),
        VN2CN5_sign => VN_sign_out(10193),
        codeword => codeword(1698),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1699 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10199 downto 10194),
        Din0 => VN1699_in0,
        Din1 => VN1699_in1,
        Din2 => VN1699_in2,
        Din3 => VN1699_in3,
        Din4 => VN1699_in4,
        Din5 => VN1699_in5,
        VN2CN0_bit => VN_data_out(10194),
        VN2CN1_bit => VN_data_out(10195),
        VN2CN2_bit => VN_data_out(10196),
        VN2CN3_bit => VN_data_out(10197),
        VN2CN4_bit => VN_data_out(10198),
        VN2CN5_bit => VN_data_out(10199),
        VN2CN0_sign => VN_sign_out(10194),
        VN2CN1_sign => VN_sign_out(10195),
        VN2CN2_sign => VN_sign_out(10196),
        VN2CN3_sign => VN_sign_out(10197),
        VN2CN4_sign => VN_sign_out(10198),
        VN2CN5_sign => VN_sign_out(10199),
        codeword => codeword(1699),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1700 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10205 downto 10200),
        Din0 => VN1700_in0,
        Din1 => VN1700_in1,
        Din2 => VN1700_in2,
        Din3 => VN1700_in3,
        Din4 => VN1700_in4,
        Din5 => VN1700_in5,
        VN2CN0_bit => VN_data_out(10200),
        VN2CN1_bit => VN_data_out(10201),
        VN2CN2_bit => VN_data_out(10202),
        VN2CN3_bit => VN_data_out(10203),
        VN2CN4_bit => VN_data_out(10204),
        VN2CN5_bit => VN_data_out(10205),
        VN2CN0_sign => VN_sign_out(10200),
        VN2CN1_sign => VN_sign_out(10201),
        VN2CN2_sign => VN_sign_out(10202),
        VN2CN3_sign => VN_sign_out(10203),
        VN2CN4_sign => VN_sign_out(10204),
        VN2CN5_sign => VN_sign_out(10205),
        codeword => codeword(1700),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1701 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10211 downto 10206),
        Din0 => VN1701_in0,
        Din1 => VN1701_in1,
        Din2 => VN1701_in2,
        Din3 => VN1701_in3,
        Din4 => VN1701_in4,
        Din5 => VN1701_in5,
        VN2CN0_bit => VN_data_out(10206),
        VN2CN1_bit => VN_data_out(10207),
        VN2CN2_bit => VN_data_out(10208),
        VN2CN3_bit => VN_data_out(10209),
        VN2CN4_bit => VN_data_out(10210),
        VN2CN5_bit => VN_data_out(10211),
        VN2CN0_sign => VN_sign_out(10206),
        VN2CN1_sign => VN_sign_out(10207),
        VN2CN2_sign => VN_sign_out(10208),
        VN2CN3_sign => VN_sign_out(10209),
        VN2CN4_sign => VN_sign_out(10210),
        VN2CN5_sign => VN_sign_out(10211),
        codeword => codeword(1701),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1702 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10217 downto 10212),
        Din0 => VN1702_in0,
        Din1 => VN1702_in1,
        Din2 => VN1702_in2,
        Din3 => VN1702_in3,
        Din4 => VN1702_in4,
        Din5 => VN1702_in5,
        VN2CN0_bit => VN_data_out(10212),
        VN2CN1_bit => VN_data_out(10213),
        VN2CN2_bit => VN_data_out(10214),
        VN2CN3_bit => VN_data_out(10215),
        VN2CN4_bit => VN_data_out(10216),
        VN2CN5_bit => VN_data_out(10217),
        VN2CN0_sign => VN_sign_out(10212),
        VN2CN1_sign => VN_sign_out(10213),
        VN2CN2_sign => VN_sign_out(10214),
        VN2CN3_sign => VN_sign_out(10215),
        VN2CN4_sign => VN_sign_out(10216),
        VN2CN5_sign => VN_sign_out(10217),
        codeword => codeword(1702),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1703 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10223 downto 10218),
        Din0 => VN1703_in0,
        Din1 => VN1703_in1,
        Din2 => VN1703_in2,
        Din3 => VN1703_in3,
        Din4 => VN1703_in4,
        Din5 => VN1703_in5,
        VN2CN0_bit => VN_data_out(10218),
        VN2CN1_bit => VN_data_out(10219),
        VN2CN2_bit => VN_data_out(10220),
        VN2CN3_bit => VN_data_out(10221),
        VN2CN4_bit => VN_data_out(10222),
        VN2CN5_bit => VN_data_out(10223),
        VN2CN0_sign => VN_sign_out(10218),
        VN2CN1_sign => VN_sign_out(10219),
        VN2CN2_sign => VN_sign_out(10220),
        VN2CN3_sign => VN_sign_out(10221),
        VN2CN4_sign => VN_sign_out(10222),
        VN2CN5_sign => VN_sign_out(10223),
        codeword => codeword(1703),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1704 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10229 downto 10224),
        Din0 => VN1704_in0,
        Din1 => VN1704_in1,
        Din2 => VN1704_in2,
        Din3 => VN1704_in3,
        Din4 => VN1704_in4,
        Din5 => VN1704_in5,
        VN2CN0_bit => VN_data_out(10224),
        VN2CN1_bit => VN_data_out(10225),
        VN2CN2_bit => VN_data_out(10226),
        VN2CN3_bit => VN_data_out(10227),
        VN2CN4_bit => VN_data_out(10228),
        VN2CN5_bit => VN_data_out(10229),
        VN2CN0_sign => VN_sign_out(10224),
        VN2CN1_sign => VN_sign_out(10225),
        VN2CN2_sign => VN_sign_out(10226),
        VN2CN3_sign => VN_sign_out(10227),
        VN2CN4_sign => VN_sign_out(10228),
        VN2CN5_sign => VN_sign_out(10229),
        codeword => codeword(1704),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1705 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10235 downto 10230),
        Din0 => VN1705_in0,
        Din1 => VN1705_in1,
        Din2 => VN1705_in2,
        Din3 => VN1705_in3,
        Din4 => VN1705_in4,
        Din5 => VN1705_in5,
        VN2CN0_bit => VN_data_out(10230),
        VN2CN1_bit => VN_data_out(10231),
        VN2CN2_bit => VN_data_out(10232),
        VN2CN3_bit => VN_data_out(10233),
        VN2CN4_bit => VN_data_out(10234),
        VN2CN5_bit => VN_data_out(10235),
        VN2CN0_sign => VN_sign_out(10230),
        VN2CN1_sign => VN_sign_out(10231),
        VN2CN2_sign => VN_sign_out(10232),
        VN2CN3_sign => VN_sign_out(10233),
        VN2CN4_sign => VN_sign_out(10234),
        VN2CN5_sign => VN_sign_out(10235),
        codeword => codeword(1705),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1706 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10241 downto 10236),
        Din0 => VN1706_in0,
        Din1 => VN1706_in1,
        Din2 => VN1706_in2,
        Din3 => VN1706_in3,
        Din4 => VN1706_in4,
        Din5 => VN1706_in5,
        VN2CN0_bit => VN_data_out(10236),
        VN2CN1_bit => VN_data_out(10237),
        VN2CN2_bit => VN_data_out(10238),
        VN2CN3_bit => VN_data_out(10239),
        VN2CN4_bit => VN_data_out(10240),
        VN2CN5_bit => VN_data_out(10241),
        VN2CN0_sign => VN_sign_out(10236),
        VN2CN1_sign => VN_sign_out(10237),
        VN2CN2_sign => VN_sign_out(10238),
        VN2CN3_sign => VN_sign_out(10239),
        VN2CN4_sign => VN_sign_out(10240),
        VN2CN5_sign => VN_sign_out(10241),
        codeword => codeword(1706),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1707 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10247 downto 10242),
        Din0 => VN1707_in0,
        Din1 => VN1707_in1,
        Din2 => VN1707_in2,
        Din3 => VN1707_in3,
        Din4 => VN1707_in4,
        Din5 => VN1707_in5,
        VN2CN0_bit => VN_data_out(10242),
        VN2CN1_bit => VN_data_out(10243),
        VN2CN2_bit => VN_data_out(10244),
        VN2CN3_bit => VN_data_out(10245),
        VN2CN4_bit => VN_data_out(10246),
        VN2CN5_bit => VN_data_out(10247),
        VN2CN0_sign => VN_sign_out(10242),
        VN2CN1_sign => VN_sign_out(10243),
        VN2CN2_sign => VN_sign_out(10244),
        VN2CN3_sign => VN_sign_out(10245),
        VN2CN4_sign => VN_sign_out(10246),
        VN2CN5_sign => VN_sign_out(10247),
        codeword => codeword(1707),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1708 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10253 downto 10248),
        Din0 => VN1708_in0,
        Din1 => VN1708_in1,
        Din2 => VN1708_in2,
        Din3 => VN1708_in3,
        Din4 => VN1708_in4,
        Din5 => VN1708_in5,
        VN2CN0_bit => VN_data_out(10248),
        VN2CN1_bit => VN_data_out(10249),
        VN2CN2_bit => VN_data_out(10250),
        VN2CN3_bit => VN_data_out(10251),
        VN2CN4_bit => VN_data_out(10252),
        VN2CN5_bit => VN_data_out(10253),
        VN2CN0_sign => VN_sign_out(10248),
        VN2CN1_sign => VN_sign_out(10249),
        VN2CN2_sign => VN_sign_out(10250),
        VN2CN3_sign => VN_sign_out(10251),
        VN2CN4_sign => VN_sign_out(10252),
        VN2CN5_sign => VN_sign_out(10253),
        codeword => codeword(1708),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1709 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10259 downto 10254),
        Din0 => VN1709_in0,
        Din1 => VN1709_in1,
        Din2 => VN1709_in2,
        Din3 => VN1709_in3,
        Din4 => VN1709_in4,
        Din5 => VN1709_in5,
        VN2CN0_bit => VN_data_out(10254),
        VN2CN1_bit => VN_data_out(10255),
        VN2CN2_bit => VN_data_out(10256),
        VN2CN3_bit => VN_data_out(10257),
        VN2CN4_bit => VN_data_out(10258),
        VN2CN5_bit => VN_data_out(10259),
        VN2CN0_sign => VN_sign_out(10254),
        VN2CN1_sign => VN_sign_out(10255),
        VN2CN2_sign => VN_sign_out(10256),
        VN2CN3_sign => VN_sign_out(10257),
        VN2CN4_sign => VN_sign_out(10258),
        VN2CN5_sign => VN_sign_out(10259),
        codeword => codeword(1709),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1710 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10265 downto 10260),
        Din0 => VN1710_in0,
        Din1 => VN1710_in1,
        Din2 => VN1710_in2,
        Din3 => VN1710_in3,
        Din4 => VN1710_in4,
        Din5 => VN1710_in5,
        VN2CN0_bit => VN_data_out(10260),
        VN2CN1_bit => VN_data_out(10261),
        VN2CN2_bit => VN_data_out(10262),
        VN2CN3_bit => VN_data_out(10263),
        VN2CN4_bit => VN_data_out(10264),
        VN2CN5_bit => VN_data_out(10265),
        VN2CN0_sign => VN_sign_out(10260),
        VN2CN1_sign => VN_sign_out(10261),
        VN2CN2_sign => VN_sign_out(10262),
        VN2CN3_sign => VN_sign_out(10263),
        VN2CN4_sign => VN_sign_out(10264),
        VN2CN5_sign => VN_sign_out(10265),
        codeword => codeword(1710),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1711 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10271 downto 10266),
        Din0 => VN1711_in0,
        Din1 => VN1711_in1,
        Din2 => VN1711_in2,
        Din3 => VN1711_in3,
        Din4 => VN1711_in4,
        Din5 => VN1711_in5,
        VN2CN0_bit => VN_data_out(10266),
        VN2CN1_bit => VN_data_out(10267),
        VN2CN2_bit => VN_data_out(10268),
        VN2CN3_bit => VN_data_out(10269),
        VN2CN4_bit => VN_data_out(10270),
        VN2CN5_bit => VN_data_out(10271),
        VN2CN0_sign => VN_sign_out(10266),
        VN2CN1_sign => VN_sign_out(10267),
        VN2CN2_sign => VN_sign_out(10268),
        VN2CN3_sign => VN_sign_out(10269),
        VN2CN4_sign => VN_sign_out(10270),
        VN2CN5_sign => VN_sign_out(10271),
        codeword => codeword(1711),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1712 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10277 downto 10272),
        Din0 => VN1712_in0,
        Din1 => VN1712_in1,
        Din2 => VN1712_in2,
        Din3 => VN1712_in3,
        Din4 => VN1712_in4,
        Din5 => VN1712_in5,
        VN2CN0_bit => VN_data_out(10272),
        VN2CN1_bit => VN_data_out(10273),
        VN2CN2_bit => VN_data_out(10274),
        VN2CN3_bit => VN_data_out(10275),
        VN2CN4_bit => VN_data_out(10276),
        VN2CN5_bit => VN_data_out(10277),
        VN2CN0_sign => VN_sign_out(10272),
        VN2CN1_sign => VN_sign_out(10273),
        VN2CN2_sign => VN_sign_out(10274),
        VN2CN3_sign => VN_sign_out(10275),
        VN2CN4_sign => VN_sign_out(10276),
        VN2CN5_sign => VN_sign_out(10277),
        codeword => codeword(1712),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1713 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10283 downto 10278),
        Din0 => VN1713_in0,
        Din1 => VN1713_in1,
        Din2 => VN1713_in2,
        Din3 => VN1713_in3,
        Din4 => VN1713_in4,
        Din5 => VN1713_in5,
        VN2CN0_bit => VN_data_out(10278),
        VN2CN1_bit => VN_data_out(10279),
        VN2CN2_bit => VN_data_out(10280),
        VN2CN3_bit => VN_data_out(10281),
        VN2CN4_bit => VN_data_out(10282),
        VN2CN5_bit => VN_data_out(10283),
        VN2CN0_sign => VN_sign_out(10278),
        VN2CN1_sign => VN_sign_out(10279),
        VN2CN2_sign => VN_sign_out(10280),
        VN2CN3_sign => VN_sign_out(10281),
        VN2CN4_sign => VN_sign_out(10282),
        VN2CN5_sign => VN_sign_out(10283),
        codeword => codeword(1713),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1714 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10289 downto 10284),
        Din0 => VN1714_in0,
        Din1 => VN1714_in1,
        Din2 => VN1714_in2,
        Din3 => VN1714_in3,
        Din4 => VN1714_in4,
        Din5 => VN1714_in5,
        VN2CN0_bit => VN_data_out(10284),
        VN2CN1_bit => VN_data_out(10285),
        VN2CN2_bit => VN_data_out(10286),
        VN2CN3_bit => VN_data_out(10287),
        VN2CN4_bit => VN_data_out(10288),
        VN2CN5_bit => VN_data_out(10289),
        VN2CN0_sign => VN_sign_out(10284),
        VN2CN1_sign => VN_sign_out(10285),
        VN2CN2_sign => VN_sign_out(10286),
        VN2CN3_sign => VN_sign_out(10287),
        VN2CN4_sign => VN_sign_out(10288),
        VN2CN5_sign => VN_sign_out(10289),
        codeword => codeword(1714),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1715 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10295 downto 10290),
        Din0 => VN1715_in0,
        Din1 => VN1715_in1,
        Din2 => VN1715_in2,
        Din3 => VN1715_in3,
        Din4 => VN1715_in4,
        Din5 => VN1715_in5,
        VN2CN0_bit => VN_data_out(10290),
        VN2CN1_bit => VN_data_out(10291),
        VN2CN2_bit => VN_data_out(10292),
        VN2CN3_bit => VN_data_out(10293),
        VN2CN4_bit => VN_data_out(10294),
        VN2CN5_bit => VN_data_out(10295),
        VN2CN0_sign => VN_sign_out(10290),
        VN2CN1_sign => VN_sign_out(10291),
        VN2CN2_sign => VN_sign_out(10292),
        VN2CN3_sign => VN_sign_out(10293),
        VN2CN4_sign => VN_sign_out(10294),
        VN2CN5_sign => VN_sign_out(10295),
        codeword => codeword(1715),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1716 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10301 downto 10296),
        Din0 => VN1716_in0,
        Din1 => VN1716_in1,
        Din2 => VN1716_in2,
        Din3 => VN1716_in3,
        Din4 => VN1716_in4,
        Din5 => VN1716_in5,
        VN2CN0_bit => VN_data_out(10296),
        VN2CN1_bit => VN_data_out(10297),
        VN2CN2_bit => VN_data_out(10298),
        VN2CN3_bit => VN_data_out(10299),
        VN2CN4_bit => VN_data_out(10300),
        VN2CN5_bit => VN_data_out(10301),
        VN2CN0_sign => VN_sign_out(10296),
        VN2CN1_sign => VN_sign_out(10297),
        VN2CN2_sign => VN_sign_out(10298),
        VN2CN3_sign => VN_sign_out(10299),
        VN2CN4_sign => VN_sign_out(10300),
        VN2CN5_sign => VN_sign_out(10301),
        codeword => codeword(1716),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1717 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10307 downto 10302),
        Din0 => VN1717_in0,
        Din1 => VN1717_in1,
        Din2 => VN1717_in2,
        Din3 => VN1717_in3,
        Din4 => VN1717_in4,
        Din5 => VN1717_in5,
        VN2CN0_bit => VN_data_out(10302),
        VN2CN1_bit => VN_data_out(10303),
        VN2CN2_bit => VN_data_out(10304),
        VN2CN3_bit => VN_data_out(10305),
        VN2CN4_bit => VN_data_out(10306),
        VN2CN5_bit => VN_data_out(10307),
        VN2CN0_sign => VN_sign_out(10302),
        VN2CN1_sign => VN_sign_out(10303),
        VN2CN2_sign => VN_sign_out(10304),
        VN2CN3_sign => VN_sign_out(10305),
        VN2CN4_sign => VN_sign_out(10306),
        VN2CN5_sign => VN_sign_out(10307),
        codeword => codeword(1717),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1718 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10313 downto 10308),
        Din0 => VN1718_in0,
        Din1 => VN1718_in1,
        Din2 => VN1718_in2,
        Din3 => VN1718_in3,
        Din4 => VN1718_in4,
        Din5 => VN1718_in5,
        VN2CN0_bit => VN_data_out(10308),
        VN2CN1_bit => VN_data_out(10309),
        VN2CN2_bit => VN_data_out(10310),
        VN2CN3_bit => VN_data_out(10311),
        VN2CN4_bit => VN_data_out(10312),
        VN2CN5_bit => VN_data_out(10313),
        VN2CN0_sign => VN_sign_out(10308),
        VN2CN1_sign => VN_sign_out(10309),
        VN2CN2_sign => VN_sign_out(10310),
        VN2CN3_sign => VN_sign_out(10311),
        VN2CN4_sign => VN_sign_out(10312),
        VN2CN5_sign => VN_sign_out(10313),
        codeword => codeword(1718),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1719 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10319 downto 10314),
        Din0 => VN1719_in0,
        Din1 => VN1719_in1,
        Din2 => VN1719_in2,
        Din3 => VN1719_in3,
        Din4 => VN1719_in4,
        Din5 => VN1719_in5,
        VN2CN0_bit => VN_data_out(10314),
        VN2CN1_bit => VN_data_out(10315),
        VN2CN2_bit => VN_data_out(10316),
        VN2CN3_bit => VN_data_out(10317),
        VN2CN4_bit => VN_data_out(10318),
        VN2CN5_bit => VN_data_out(10319),
        VN2CN0_sign => VN_sign_out(10314),
        VN2CN1_sign => VN_sign_out(10315),
        VN2CN2_sign => VN_sign_out(10316),
        VN2CN3_sign => VN_sign_out(10317),
        VN2CN4_sign => VN_sign_out(10318),
        VN2CN5_sign => VN_sign_out(10319),
        codeword => codeword(1719),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1720 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10325 downto 10320),
        Din0 => VN1720_in0,
        Din1 => VN1720_in1,
        Din2 => VN1720_in2,
        Din3 => VN1720_in3,
        Din4 => VN1720_in4,
        Din5 => VN1720_in5,
        VN2CN0_bit => VN_data_out(10320),
        VN2CN1_bit => VN_data_out(10321),
        VN2CN2_bit => VN_data_out(10322),
        VN2CN3_bit => VN_data_out(10323),
        VN2CN4_bit => VN_data_out(10324),
        VN2CN5_bit => VN_data_out(10325),
        VN2CN0_sign => VN_sign_out(10320),
        VN2CN1_sign => VN_sign_out(10321),
        VN2CN2_sign => VN_sign_out(10322),
        VN2CN3_sign => VN_sign_out(10323),
        VN2CN4_sign => VN_sign_out(10324),
        VN2CN5_sign => VN_sign_out(10325),
        codeword => codeword(1720),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1721 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10331 downto 10326),
        Din0 => VN1721_in0,
        Din1 => VN1721_in1,
        Din2 => VN1721_in2,
        Din3 => VN1721_in3,
        Din4 => VN1721_in4,
        Din5 => VN1721_in5,
        VN2CN0_bit => VN_data_out(10326),
        VN2CN1_bit => VN_data_out(10327),
        VN2CN2_bit => VN_data_out(10328),
        VN2CN3_bit => VN_data_out(10329),
        VN2CN4_bit => VN_data_out(10330),
        VN2CN5_bit => VN_data_out(10331),
        VN2CN0_sign => VN_sign_out(10326),
        VN2CN1_sign => VN_sign_out(10327),
        VN2CN2_sign => VN_sign_out(10328),
        VN2CN3_sign => VN_sign_out(10329),
        VN2CN4_sign => VN_sign_out(10330),
        VN2CN5_sign => VN_sign_out(10331),
        codeword => codeword(1721),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1722 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10337 downto 10332),
        Din0 => VN1722_in0,
        Din1 => VN1722_in1,
        Din2 => VN1722_in2,
        Din3 => VN1722_in3,
        Din4 => VN1722_in4,
        Din5 => VN1722_in5,
        VN2CN0_bit => VN_data_out(10332),
        VN2CN1_bit => VN_data_out(10333),
        VN2CN2_bit => VN_data_out(10334),
        VN2CN3_bit => VN_data_out(10335),
        VN2CN4_bit => VN_data_out(10336),
        VN2CN5_bit => VN_data_out(10337),
        VN2CN0_sign => VN_sign_out(10332),
        VN2CN1_sign => VN_sign_out(10333),
        VN2CN2_sign => VN_sign_out(10334),
        VN2CN3_sign => VN_sign_out(10335),
        VN2CN4_sign => VN_sign_out(10336),
        VN2CN5_sign => VN_sign_out(10337),
        codeword => codeword(1722),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1723 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10343 downto 10338),
        Din0 => VN1723_in0,
        Din1 => VN1723_in1,
        Din2 => VN1723_in2,
        Din3 => VN1723_in3,
        Din4 => VN1723_in4,
        Din5 => VN1723_in5,
        VN2CN0_bit => VN_data_out(10338),
        VN2CN1_bit => VN_data_out(10339),
        VN2CN2_bit => VN_data_out(10340),
        VN2CN3_bit => VN_data_out(10341),
        VN2CN4_bit => VN_data_out(10342),
        VN2CN5_bit => VN_data_out(10343),
        VN2CN0_sign => VN_sign_out(10338),
        VN2CN1_sign => VN_sign_out(10339),
        VN2CN2_sign => VN_sign_out(10340),
        VN2CN3_sign => VN_sign_out(10341),
        VN2CN4_sign => VN_sign_out(10342),
        VN2CN5_sign => VN_sign_out(10343),
        codeword => codeword(1723),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1724 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10349 downto 10344),
        Din0 => VN1724_in0,
        Din1 => VN1724_in1,
        Din2 => VN1724_in2,
        Din3 => VN1724_in3,
        Din4 => VN1724_in4,
        Din5 => VN1724_in5,
        VN2CN0_bit => VN_data_out(10344),
        VN2CN1_bit => VN_data_out(10345),
        VN2CN2_bit => VN_data_out(10346),
        VN2CN3_bit => VN_data_out(10347),
        VN2CN4_bit => VN_data_out(10348),
        VN2CN5_bit => VN_data_out(10349),
        VN2CN0_sign => VN_sign_out(10344),
        VN2CN1_sign => VN_sign_out(10345),
        VN2CN2_sign => VN_sign_out(10346),
        VN2CN3_sign => VN_sign_out(10347),
        VN2CN4_sign => VN_sign_out(10348),
        VN2CN5_sign => VN_sign_out(10349),
        codeword => codeword(1724),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1725 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10355 downto 10350),
        Din0 => VN1725_in0,
        Din1 => VN1725_in1,
        Din2 => VN1725_in2,
        Din3 => VN1725_in3,
        Din4 => VN1725_in4,
        Din5 => VN1725_in5,
        VN2CN0_bit => VN_data_out(10350),
        VN2CN1_bit => VN_data_out(10351),
        VN2CN2_bit => VN_data_out(10352),
        VN2CN3_bit => VN_data_out(10353),
        VN2CN4_bit => VN_data_out(10354),
        VN2CN5_bit => VN_data_out(10355),
        VN2CN0_sign => VN_sign_out(10350),
        VN2CN1_sign => VN_sign_out(10351),
        VN2CN2_sign => VN_sign_out(10352),
        VN2CN3_sign => VN_sign_out(10353),
        VN2CN4_sign => VN_sign_out(10354),
        VN2CN5_sign => VN_sign_out(10355),
        codeword => codeword(1725),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1726 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10361 downto 10356),
        Din0 => VN1726_in0,
        Din1 => VN1726_in1,
        Din2 => VN1726_in2,
        Din3 => VN1726_in3,
        Din4 => VN1726_in4,
        Din5 => VN1726_in5,
        VN2CN0_bit => VN_data_out(10356),
        VN2CN1_bit => VN_data_out(10357),
        VN2CN2_bit => VN_data_out(10358),
        VN2CN3_bit => VN_data_out(10359),
        VN2CN4_bit => VN_data_out(10360),
        VN2CN5_bit => VN_data_out(10361),
        VN2CN0_sign => VN_sign_out(10356),
        VN2CN1_sign => VN_sign_out(10357),
        VN2CN2_sign => VN_sign_out(10358),
        VN2CN3_sign => VN_sign_out(10359),
        VN2CN4_sign => VN_sign_out(10360),
        VN2CN5_sign => VN_sign_out(10361),
        codeword => codeword(1726),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1727 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10367 downto 10362),
        Din0 => VN1727_in0,
        Din1 => VN1727_in1,
        Din2 => VN1727_in2,
        Din3 => VN1727_in3,
        Din4 => VN1727_in4,
        Din5 => VN1727_in5,
        VN2CN0_bit => VN_data_out(10362),
        VN2CN1_bit => VN_data_out(10363),
        VN2CN2_bit => VN_data_out(10364),
        VN2CN3_bit => VN_data_out(10365),
        VN2CN4_bit => VN_data_out(10366),
        VN2CN5_bit => VN_data_out(10367),
        VN2CN0_sign => VN_sign_out(10362),
        VN2CN1_sign => VN_sign_out(10363),
        VN2CN2_sign => VN_sign_out(10364),
        VN2CN3_sign => VN_sign_out(10365),
        VN2CN4_sign => VN_sign_out(10366),
        VN2CN5_sign => VN_sign_out(10367),
        codeword => codeword(1727),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1728 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10373 downto 10368),
        Din0 => VN1728_in0,
        Din1 => VN1728_in1,
        Din2 => VN1728_in2,
        Din3 => VN1728_in3,
        Din4 => VN1728_in4,
        Din5 => VN1728_in5,
        VN2CN0_bit => VN_data_out(10368),
        VN2CN1_bit => VN_data_out(10369),
        VN2CN2_bit => VN_data_out(10370),
        VN2CN3_bit => VN_data_out(10371),
        VN2CN4_bit => VN_data_out(10372),
        VN2CN5_bit => VN_data_out(10373),
        VN2CN0_sign => VN_sign_out(10368),
        VN2CN1_sign => VN_sign_out(10369),
        VN2CN2_sign => VN_sign_out(10370),
        VN2CN3_sign => VN_sign_out(10371),
        VN2CN4_sign => VN_sign_out(10372),
        VN2CN5_sign => VN_sign_out(10373),
        codeword => codeword(1728),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1729 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10379 downto 10374),
        Din0 => VN1729_in0,
        Din1 => VN1729_in1,
        Din2 => VN1729_in2,
        Din3 => VN1729_in3,
        Din4 => VN1729_in4,
        Din5 => VN1729_in5,
        VN2CN0_bit => VN_data_out(10374),
        VN2CN1_bit => VN_data_out(10375),
        VN2CN2_bit => VN_data_out(10376),
        VN2CN3_bit => VN_data_out(10377),
        VN2CN4_bit => VN_data_out(10378),
        VN2CN5_bit => VN_data_out(10379),
        VN2CN0_sign => VN_sign_out(10374),
        VN2CN1_sign => VN_sign_out(10375),
        VN2CN2_sign => VN_sign_out(10376),
        VN2CN3_sign => VN_sign_out(10377),
        VN2CN4_sign => VN_sign_out(10378),
        VN2CN5_sign => VN_sign_out(10379),
        codeword => codeword(1729),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1730 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10385 downto 10380),
        Din0 => VN1730_in0,
        Din1 => VN1730_in1,
        Din2 => VN1730_in2,
        Din3 => VN1730_in3,
        Din4 => VN1730_in4,
        Din5 => VN1730_in5,
        VN2CN0_bit => VN_data_out(10380),
        VN2CN1_bit => VN_data_out(10381),
        VN2CN2_bit => VN_data_out(10382),
        VN2CN3_bit => VN_data_out(10383),
        VN2CN4_bit => VN_data_out(10384),
        VN2CN5_bit => VN_data_out(10385),
        VN2CN0_sign => VN_sign_out(10380),
        VN2CN1_sign => VN_sign_out(10381),
        VN2CN2_sign => VN_sign_out(10382),
        VN2CN3_sign => VN_sign_out(10383),
        VN2CN4_sign => VN_sign_out(10384),
        VN2CN5_sign => VN_sign_out(10385),
        codeword => codeword(1730),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1731 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10391 downto 10386),
        Din0 => VN1731_in0,
        Din1 => VN1731_in1,
        Din2 => VN1731_in2,
        Din3 => VN1731_in3,
        Din4 => VN1731_in4,
        Din5 => VN1731_in5,
        VN2CN0_bit => VN_data_out(10386),
        VN2CN1_bit => VN_data_out(10387),
        VN2CN2_bit => VN_data_out(10388),
        VN2CN3_bit => VN_data_out(10389),
        VN2CN4_bit => VN_data_out(10390),
        VN2CN5_bit => VN_data_out(10391),
        VN2CN0_sign => VN_sign_out(10386),
        VN2CN1_sign => VN_sign_out(10387),
        VN2CN2_sign => VN_sign_out(10388),
        VN2CN3_sign => VN_sign_out(10389),
        VN2CN4_sign => VN_sign_out(10390),
        VN2CN5_sign => VN_sign_out(10391),
        codeword => codeword(1731),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1732 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10397 downto 10392),
        Din0 => VN1732_in0,
        Din1 => VN1732_in1,
        Din2 => VN1732_in2,
        Din3 => VN1732_in3,
        Din4 => VN1732_in4,
        Din5 => VN1732_in5,
        VN2CN0_bit => VN_data_out(10392),
        VN2CN1_bit => VN_data_out(10393),
        VN2CN2_bit => VN_data_out(10394),
        VN2CN3_bit => VN_data_out(10395),
        VN2CN4_bit => VN_data_out(10396),
        VN2CN5_bit => VN_data_out(10397),
        VN2CN0_sign => VN_sign_out(10392),
        VN2CN1_sign => VN_sign_out(10393),
        VN2CN2_sign => VN_sign_out(10394),
        VN2CN3_sign => VN_sign_out(10395),
        VN2CN4_sign => VN_sign_out(10396),
        VN2CN5_sign => VN_sign_out(10397),
        codeword => codeword(1732),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1733 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10403 downto 10398),
        Din0 => VN1733_in0,
        Din1 => VN1733_in1,
        Din2 => VN1733_in2,
        Din3 => VN1733_in3,
        Din4 => VN1733_in4,
        Din5 => VN1733_in5,
        VN2CN0_bit => VN_data_out(10398),
        VN2CN1_bit => VN_data_out(10399),
        VN2CN2_bit => VN_data_out(10400),
        VN2CN3_bit => VN_data_out(10401),
        VN2CN4_bit => VN_data_out(10402),
        VN2CN5_bit => VN_data_out(10403),
        VN2CN0_sign => VN_sign_out(10398),
        VN2CN1_sign => VN_sign_out(10399),
        VN2CN2_sign => VN_sign_out(10400),
        VN2CN3_sign => VN_sign_out(10401),
        VN2CN4_sign => VN_sign_out(10402),
        VN2CN5_sign => VN_sign_out(10403),
        codeword => codeword(1733),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1734 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10409 downto 10404),
        Din0 => VN1734_in0,
        Din1 => VN1734_in1,
        Din2 => VN1734_in2,
        Din3 => VN1734_in3,
        Din4 => VN1734_in4,
        Din5 => VN1734_in5,
        VN2CN0_bit => VN_data_out(10404),
        VN2CN1_bit => VN_data_out(10405),
        VN2CN2_bit => VN_data_out(10406),
        VN2CN3_bit => VN_data_out(10407),
        VN2CN4_bit => VN_data_out(10408),
        VN2CN5_bit => VN_data_out(10409),
        VN2CN0_sign => VN_sign_out(10404),
        VN2CN1_sign => VN_sign_out(10405),
        VN2CN2_sign => VN_sign_out(10406),
        VN2CN3_sign => VN_sign_out(10407),
        VN2CN4_sign => VN_sign_out(10408),
        VN2CN5_sign => VN_sign_out(10409),
        codeword => codeword(1734),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1735 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10415 downto 10410),
        Din0 => VN1735_in0,
        Din1 => VN1735_in1,
        Din2 => VN1735_in2,
        Din3 => VN1735_in3,
        Din4 => VN1735_in4,
        Din5 => VN1735_in5,
        VN2CN0_bit => VN_data_out(10410),
        VN2CN1_bit => VN_data_out(10411),
        VN2CN2_bit => VN_data_out(10412),
        VN2CN3_bit => VN_data_out(10413),
        VN2CN4_bit => VN_data_out(10414),
        VN2CN5_bit => VN_data_out(10415),
        VN2CN0_sign => VN_sign_out(10410),
        VN2CN1_sign => VN_sign_out(10411),
        VN2CN2_sign => VN_sign_out(10412),
        VN2CN3_sign => VN_sign_out(10413),
        VN2CN4_sign => VN_sign_out(10414),
        VN2CN5_sign => VN_sign_out(10415),
        codeword => codeword(1735),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1736 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10421 downto 10416),
        Din0 => VN1736_in0,
        Din1 => VN1736_in1,
        Din2 => VN1736_in2,
        Din3 => VN1736_in3,
        Din4 => VN1736_in4,
        Din5 => VN1736_in5,
        VN2CN0_bit => VN_data_out(10416),
        VN2CN1_bit => VN_data_out(10417),
        VN2CN2_bit => VN_data_out(10418),
        VN2CN3_bit => VN_data_out(10419),
        VN2CN4_bit => VN_data_out(10420),
        VN2CN5_bit => VN_data_out(10421),
        VN2CN0_sign => VN_sign_out(10416),
        VN2CN1_sign => VN_sign_out(10417),
        VN2CN2_sign => VN_sign_out(10418),
        VN2CN3_sign => VN_sign_out(10419),
        VN2CN4_sign => VN_sign_out(10420),
        VN2CN5_sign => VN_sign_out(10421),
        codeword => codeword(1736),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1737 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10427 downto 10422),
        Din0 => VN1737_in0,
        Din1 => VN1737_in1,
        Din2 => VN1737_in2,
        Din3 => VN1737_in3,
        Din4 => VN1737_in4,
        Din5 => VN1737_in5,
        VN2CN0_bit => VN_data_out(10422),
        VN2CN1_bit => VN_data_out(10423),
        VN2CN2_bit => VN_data_out(10424),
        VN2CN3_bit => VN_data_out(10425),
        VN2CN4_bit => VN_data_out(10426),
        VN2CN5_bit => VN_data_out(10427),
        VN2CN0_sign => VN_sign_out(10422),
        VN2CN1_sign => VN_sign_out(10423),
        VN2CN2_sign => VN_sign_out(10424),
        VN2CN3_sign => VN_sign_out(10425),
        VN2CN4_sign => VN_sign_out(10426),
        VN2CN5_sign => VN_sign_out(10427),
        codeword => codeword(1737),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1738 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10433 downto 10428),
        Din0 => VN1738_in0,
        Din1 => VN1738_in1,
        Din2 => VN1738_in2,
        Din3 => VN1738_in3,
        Din4 => VN1738_in4,
        Din5 => VN1738_in5,
        VN2CN0_bit => VN_data_out(10428),
        VN2CN1_bit => VN_data_out(10429),
        VN2CN2_bit => VN_data_out(10430),
        VN2CN3_bit => VN_data_out(10431),
        VN2CN4_bit => VN_data_out(10432),
        VN2CN5_bit => VN_data_out(10433),
        VN2CN0_sign => VN_sign_out(10428),
        VN2CN1_sign => VN_sign_out(10429),
        VN2CN2_sign => VN_sign_out(10430),
        VN2CN3_sign => VN_sign_out(10431),
        VN2CN4_sign => VN_sign_out(10432),
        VN2CN5_sign => VN_sign_out(10433),
        codeword => codeword(1738),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1739 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10439 downto 10434),
        Din0 => VN1739_in0,
        Din1 => VN1739_in1,
        Din2 => VN1739_in2,
        Din3 => VN1739_in3,
        Din4 => VN1739_in4,
        Din5 => VN1739_in5,
        VN2CN0_bit => VN_data_out(10434),
        VN2CN1_bit => VN_data_out(10435),
        VN2CN2_bit => VN_data_out(10436),
        VN2CN3_bit => VN_data_out(10437),
        VN2CN4_bit => VN_data_out(10438),
        VN2CN5_bit => VN_data_out(10439),
        VN2CN0_sign => VN_sign_out(10434),
        VN2CN1_sign => VN_sign_out(10435),
        VN2CN2_sign => VN_sign_out(10436),
        VN2CN3_sign => VN_sign_out(10437),
        VN2CN4_sign => VN_sign_out(10438),
        VN2CN5_sign => VN_sign_out(10439),
        codeword => codeword(1739),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1740 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10445 downto 10440),
        Din0 => VN1740_in0,
        Din1 => VN1740_in1,
        Din2 => VN1740_in2,
        Din3 => VN1740_in3,
        Din4 => VN1740_in4,
        Din5 => VN1740_in5,
        VN2CN0_bit => VN_data_out(10440),
        VN2CN1_bit => VN_data_out(10441),
        VN2CN2_bit => VN_data_out(10442),
        VN2CN3_bit => VN_data_out(10443),
        VN2CN4_bit => VN_data_out(10444),
        VN2CN5_bit => VN_data_out(10445),
        VN2CN0_sign => VN_sign_out(10440),
        VN2CN1_sign => VN_sign_out(10441),
        VN2CN2_sign => VN_sign_out(10442),
        VN2CN3_sign => VN_sign_out(10443),
        VN2CN4_sign => VN_sign_out(10444),
        VN2CN5_sign => VN_sign_out(10445),
        codeword => codeword(1740),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1741 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10451 downto 10446),
        Din0 => VN1741_in0,
        Din1 => VN1741_in1,
        Din2 => VN1741_in2,
        Din3 => VN1741_in3,
        Din4 => VN1741_in4,
        Din5 => VN1741_in5,
        VN2CN0_bit => VN_data_out(10446),
        VN2CN1_bit => VN_data_out(10447),
        VN2CN2_bit => VN_data_out(10448),
        VN2CN3_bit => VN_data_out(10449),
        VN2CN4_bit => VN_data_out(10450),
        VN2CN5_bit => VN_data_out(10451),
        VN2CN0_sign => VN_sign_out(10446),
        VN2CN1_sign => VN_sign_out(10447),
        VN2CN2_sign => VN_sign_out(10448),
        VN2CN3_sign => VN_sign_out(10449),
        VN2CN4_sign => VN_sign_out(10450),
        VN2CN5_sign => VN_sign_out(10451),
        codeword => codeword(1741),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1742 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10457 downto 10452),
        Din0 => VN1742_in0,
        Din1 => VN1742_in1,
        Din2 => VN1742_in2,
        Din3 => VN1742_in3,
        Din4 => VN1742_in4,
        Din5 => VN1742_in5,
        VN2CN0_bit => VN_data_out(10452),
        VN2CN1_bit => VN_data_out(10453),
        VN2CN2_bit => VN_data_out(10454),
        VN2CN3_bit => VN_data_out(10455),
        VN2CN4_bit => VN_data_out(10456),
        VN2CN5_bit => VN_data_out(10457),
        VN2CN0_sign => VN_sign_out(10452),
        VN2CN1_sign => VN_sign_out(10453),
        VN2CN2_sign => VN_sign_out(10454),
        VN2CN3_sign => VN_sign_out(10455),
        VN2CN4_sign => VN_sign_out(10456),
        VN2CN5_sign => VN_sign_out(10457),
        codeword => codeword(1742),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1743 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10463 downto 10458),
        Din0 => VN1743_in0,
        Din1 => VN1743_in1,
        Din2 => VN1743_in2,
        Din3 => VN1743_in3,
        Din4 => VN1743_in4,
        Din5 => VN1743_in5,
        VN2CN0_bit => VN_data_out(10458),
        VN2CN1_bit => VN_data_out(10459),
        VN2CN2_bit => VN_data_out(10460),
        VN2CN3_bit => VN_data_out(10461),
        VN2CN4_bit => VN_data_out(10462),
        VN2CN5_bit => VN_data_out(10463),
        VN2CN0_sign => VN_sign_out(10458),
        VN2CN1_sign => VN_sign_out(10459),
        VN2CN2_sign => VN_sign_out(10460),
        VN2CN3_sign => VN_sign_out(10461),
        VN2CN4_sign => VN_sign_out(10462),
        VN2CN5_sign => VN_sign_out(10463),
        codeword => codeword(1743),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1744 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10469 downto 10464),
        Din0 => VN1744_in0,
        Din1 => VN1744_in1,
        Din2 => VN1744_in2,
        Din3 => VN1744_in3,
        Din4 => VN1744_in4,
        Din5 => VN1744_in5,
        VN2CN0_bit => VN_data_out(10464),
        VN2CN1_bit => VN_data_out(10465),
        VN2CN2_bit => VN_data_out(10466),
        VN2CN3_bit => VN_data_out(10467),
        VN2CN4_bit => VN_data_out(10468),
        VN2CN5_bit => VN_data_out(10469),
        VN2CN0_sign => VN_sign_out(10464),
        VN2CN1_sign => VN_sign_out(10465),
        VN2CN2_sign => VN_sign_out(10466),
        VN2CN3_sign => VN_sign_out(10467),
        VN2CN4_sign => VN_sign_out(10468),
        VN2CN5_sign => VN_sign_out(10469),
        codeword => codeword(1744),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1745 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10475 downto 10470),
        Din0 => VN1745_in0,
        Din1 => VN1745_in1,
        Din2 => VN1745_in2,
        Din3 => VN1745_in3,
        Din4 => VN1745_in4,
        Din5 => VN1745_in5,
        VN2CN0_bit => VN_data_out(10470),
        VN2CN1_bit => VN_data_out(10471),
        VN2CN2_bit => VN_data_out(10472),
        VN2CN3_bit => VN_data_out(10473),
        VN2CN4_bit => VN_data_out(10474),
        VN2CN5_bit => VN_data_out(10475),
        VN2CN0_sign => VN_sign_out(10470),
        VN2CN1_sign => VN_sign_out(10471),
        VN2CN2_sign => VN_sign_out(10472),
        VN2CN3_sign => VN_sign_out(10473),
        VN2CN4_sign => VN_sign_out(10474),
        VN2CN5_sign => VN_sign_out(10475),
        codeword => codeword(1745),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1746 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10481 downto 10476),
        Din0 => VN1746_in0,
        Din1 => VN1746_in1,
        Din2 => VN1746_in2,
        Din3 => VN1746_in3,
        Din4 => VN1746_in4,
        Din5 => VN1746_in5,
        VN2CN0_bit => VN_data_out(10476),
        VN2CN1_bit => VN_data_out(10477),
        VN2CN2_bit => VN_data_out(10478),
        VN2CN3_bit => VN_data_out(10479),
        VN2CN4_bit => VN_data_out(10480),
        VN2CN5_bit => VN_data_out(10481),
        VN2CN0_sign => VN_sign_out(10476),
        VN2CN1_sign => VN_sign_out(10477),
        VN2CN2_sign => VN_sign_out(10478),
        VN2CN3_sign => VN_sign_out(10479),
        VN2CN4_sign => VN_sign_out(10480),
        VN2CN5_sign => VN_sign_out(10481),
        codeword => codeword(1746),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1747 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10487 downto 10482),
        Din0 => VN1747_in0,
        Din1 => VN1747_in1,
        Din2 => VN1747_in2,
        Din3 => VN1747_in3,
        Din4 => VN1747_in4,
        Din5 => VN1747_in5,
        VN2CN0_bit => VN_data_out(10482),
        VN2CN1_bit => VN_data_out(10483),
        VN2CN2_bit => VN_data_out(10484),
        VN2CN3_bit => VN_data_out(10485),
        VN2CN4_bit => VN_data_out(10486),
        VN2CN5_bit => VN_data_out(10487),
        VN2CN0_sign => VN_sign_out(10482),
        VN2CN1_sign => VN_sign_out(10483),
        VN2CN2_sign => VN_sign_out(10484),
        VN2CN3_sign => VN_sign_out(10485),
        VN2CN4_sign => VN_sign_out(10486),
        VN2CN5_sign => VN_sign_out(10487),
        codeword => codeword(1747),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1748 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10493 downto 10488),
        Din0 => VN1748_in0,
        Din1 => VN1748_in1,
        Din2 => VN1748_in2,
        Din3 => VN1748_in3,
        Din4 => VN1748_in4,
        Din5 => VN1748_in5,
        VN2CN0_bit => VN_data_out(10488),
        VN2CN1_bit => VN_data_out(10489),
        VN2CN2_bit => VN_data_out(10490),
        VN2CN3_bit => VN_data_out(10491),
        VN2CN4_bit => VN_data_out(10492),
        VN2CN5_bit => VN_data_out(10493),
        VN2CN0_sign => VN_sign_out(10488),
        VN2CN1_sign => VN_sign_out(10489),
        VN2CN2_sign => VN_sign_out(10490),
        VN2CN3_sign => VN_sign_out(10491),
        VN2CN4_sign => VN_sign_out(10492),
        VN2CN5_sign => VN_sign_out(10493),
        codeword => codeword(1748),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1749 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10499 downto 10494),
        Din0 => VN1749_in0,
        Din1 => VN1749_in1,
        Din2 => VN1749_in2,
        Din3 => VN1749_in3,
        Din4 => VN1749_in4,
        Din5 => VN1749_in5,
        VN2CN0_bit => VN_data_out(10494),
        VN2CN1_bit => VN_data_out(10495),
        VN2CN2_bit => VN_data_out(10496),
        VN2CN3_bit => VN_data_out(10497),
        VN2CN4_bit => VN_data_out(10498),
        VN2CN5_bit => VN_data_out(10499),
        VN2CN0_sign => VN_sign_out(10494),
        VN2CN1_sign => VN_sign_out(10495),
        VN2CN2_sign => VN_sign_out(10496),
        VN2CN3_sign => VN_sign_out(10497),
        VN2CN4_sign => VN_sign_out(10498),
        VN2CN5_sign => VN_sign_out(10499),
        codeword => codeword(1749),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1750 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10505 downto 10500),
        Din0 => VN1750_in0,
        Din1 => VN1750_in1,
        Din2 => VN1750_in2,
        Din3 => VN1750_in3,
        Din4 => VN1750_in4,
        Din5 => VN1750_in5,
        VN2CN0_bit => VN_data_out(10500),
        VN2CN1_bit => VN_data_out(10501),
        VN2CN2_bit => VN_data_out(10502),
        VN2CN3_bit => VN_data_out(10503),
        VN2CN4_bit => VN_data_out(10504),
        VN2CN5_bit => VN_data_out(10505),
        VN2CN0_sign => VN_sign_out(10500),
        VN2CN1_sign => VN_sign_out(10501),
        VN2CN2_sign => VN_sign_out(10502),
        VN2CN3_sign => VN_sign_out(10503),
        VN2CN4_sign => VN_sign_out(10504),
        VN2CN5_sign => VN_sign_out(10505),
        codeword => codeword(1750),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1751 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10511 downto 10506),
        Din0 => VN1751_in0,
        Din1 => VN1751_in1,
        Din2 => VN1751_in2,
        Din3 => VN1751_in3,
        Din4 => VN1751_in4,
        Din5 => VN1751_in5,
        VN2CN0_bit => VN_data_out(10506),
        VN2CN1_bit => VN_data_out(10507),
        VN2CN2_bit => VN_data_out(10508),
        VN2CN3_bit => VN_data_out(10509),
        VN2CN4_bit => VN_data_out(10510),
        VN2CN5_bit => VN_data_out(10511),
        VN2CN0_sign => VN_sign_out(10506),
        VN2CN1_sign => VN_sign_out(10507),
        VN2CN2_sign => VN_sign_out(10508),
        VN2CN3_sign => VN_sign_out(10509),
        VN2CN4_sign => VN_sign_out(10510),
        VN2CN5_sign => VN_sign_out(10511),
        codeword => codeword(1751),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1752 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10517 downto 10512),
        Din0 => VN1752_in0,
        Din1 => VN1752_in1,
        Din2 => VN1752_in2,
        Din3 => VN1752_in3,
        Din4 => VN1752_in4,
        Din5 => VN1752_in5,
        VN2CN0_bit => VN_data_out(10512),
        VN2CN1_bit => VN_data_out(10513),
        VN2CN2_bit => VN_data_out(10514),
        VN2CN3_bit => VN_data_out(10515),
        VN2CN4_bit => VN_data_out(10516),
        VN2CN5_bit => VN_data_out(10517),
        VN2CN0_sign => VN_sign_out(10512),
        VN2CN1_sign => VN_sign_out(10513),
        VN2CN2_sign => VN_sign_out(10514),
        VN2CN3_sign => VN_sign_out(10515),
        VN2CN4_sign => VN_sign_out(10516),
        VN2CN5_sign => VN_sign_out(10517),
        codeword => codeword(1752),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1753 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10523 downto 10518),
        Din0 => VN1753_in0,
        Din1 => VN1753_in1,
        Din2 => VN1753_in2,
        Din3 => VN1753_in3,
        Din4 => VN1753_in4,
        Din5 => VN1753_in5,
        VN2CN0_bit => VN_data_out(10518),
        VN2CN1_bit => VN_data_out(10519),
        VN2CN2_bit => VN_data_out(10520),
        VN2CN3_bit => VN_data_out(10521),
        VN2CN4_bit => VN_data_out(10522),
        VN2CN5_bit => VN_data_out(10523),
        VN2CN0_sign => VN_sign_out(10518),
        VN2CN1_sign => VN_sign_out(10519),
        VN2CN2_sign => VN_sign_out(10520),
        VN2CN3_sign => VN_sign_out(10521),
        VN2CN4_sign => VN_sign_out(10522),
        VN2CN5_sign => VN_sign_out(10523),
        codeword => codeword(1753),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1754 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10529 downto 10524),
        Din0 => VN1754_in0,
        Din1 => VN1754_in1,
        Din2 => VN1754_in2,
        Din3 => VN1754_in3,
        Din4 => VN1754_in4,
        Din5 => VN1754_in5,
        VN2CN0_bit => VN_data_out(10524),
        VN2CN1_bit => VN_data_out(10525),
        VN2CN2_bit => VN_data_out(10526),
        VN2CN3_bit => VN_data_out(10527),
        VN2CN4_bit => VN_data_out(10528),
        VN2CN5_bit => VN_data_out(10529),
        VN2CN0_sign => VN_sign_out(10524),
        VN2CN1_sign => VN_sign_out(10525),
        VN2CN2_sign => VN_sign_out(10526),
        VN2CN3_sign => VN_sign_out(10527),
        VN2CN4_sign => VN_sign_out(10528),
        VN2CN5_sign => VN_sign_out(10529),
        codeword => codeword(1754),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1755 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10535 downto 10530),
        Din0 => VN1755_in0,
        Din1 => VN1755_in1,
        Din2 => VN1755_in2,
        Din3 => VN1755_in3,
        Din4 => VN1755_in4,
        Din5 => VN1755_in5,
        VN2CN0_bit => VN_data_out(10530),
        VN2CN1_bit => VN_data_out(10531),
        VN2CN2_bit => VN_data_out(10532),
        VN2CN3_bit => VN_data_out(10533),
        VN2CN4_bit => VN_data_out(10534),
        VN2CN5_bit => VN_data_out(10535),
        VN2CN0_sign => VN_sign_out(10530),
        VN2CN1_sign => VN_sign_out(10531),
        VN2CN2_sign => VN_sign_out(10532),
        VN2CN3_sign => VN_sign_out(10533),
        VN2CN4_sign => VN_sign_out(10534),
        VN2CN5_sign => VN_sign_out(10535),
        codeword => codeword(1755),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1756 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10541 downto 10536),
        Din0 => VN1756_in0,
        Din1 => VN1756_in1,
        Din2 => VN1756_in2,
        Din3 => VN1756_in3,
        Din4 => VN1756_in4,
        Din5 => VN1756_in5,
        VN2CN0_bit => VN_data_out(10536),
        VN2CN1_bit => VN_data_out(10537),
        VN2CN2_bit => VN_data_out(10538),
        VN2CN3_bit => VN_data_out(10539),
        VN2CN4_bit => VN_data_out(10540),
        VN2CN5_bit => VN_data_out(10541),
        VN2CN0_sign => VN_sign_out(10536),
        VN2CN1_sign => VN_sign_out(10537),
        VN2CN2_sign => VN_sign_out(10538),
        VN2CN3_sign => VN_sign_out(10539),
        VN2CN4_sign => VN_sign_out(10540),
        VN2CN5_sign => VN_sign_out(10541),
        codeword => codeword(1756),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1757 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10547 downto 10542),
        Din0 => VN1757_in0,
        Din1 => VN1757_in1,
        Din2 => VN1757_in2,
        Din3 => VN1757_in3,
        Din4 => VN1757_in4,
        Din5 => VN1757_in5,
        VN2CN0_bit => VN_data_out(10542),
        VN2CN1_bit => VN_data_out(10543),
        VN2CN2_bit => VN_data_out(10544),
        VN2CN3_bit => VN_data_out(10545),
        VN2CN4_bit => VN_data_out(10546),
        VN2CN5_bit => VN_data_out(10547),
        VN2CN0_sign => VN_sign_out(10542),
        VN2CN1_sign => VN_sign_out(10543),
        VN2CN2_sign => VN_sign_out(10544),
        VN2CN3_sign => VN_sign_out(10545),
        VN2CN4_sign => VN_sign_out(10546),
        VN2CN5_sign => VN_sign_out(10547),
        codeword => codeword(1757),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1758 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10553 downto 10548),
        Din0 => VN1758_in0,
        Din1 => VN1758_in1,
        Din2 => VN1758_in2,
        Din3 => VN1758_in3,
        Din4 => VN1758_in4,
        Din5 => VN1758_in5,
        VN2CN0_bit => VN_data_out(10548),
        VN2CN1_bit => VN_data_out(10549),
        VN2CN2_bit => VN_data_out(10550),
        VN2CN3_bit => VN_data_out(10551),
        VN2CN4_bit => VN_data_out(10552),
        VN2CN5_bit => VN_data_out(10553),
        VN2CN0_sign => VN_sign_out(10548),
        VN2CN1_sign => VN_sign_out(10549),
        VN2CN2_sign => VN_sign_out(10550),
        VN2CN3_sign => VN_sign_out(10551),
        VN2CN4_sign => VN_sign_out(10552),
        VN2CN5_sign => VN_sign_out(10553),
        codeword => codeword(1758),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1759 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10559 downto 10554),
        Din0 => VN1759_in0,
        Din1 => VN1759_in1,
        Din2 => VN1759_in2,
        Din3 => VN1759_in3,
        Din4 => VN1759_in4,
        Din5 => VN1759_in5,
        VN2CN0_bit => VN_data_out(10554),
        VN2CN1_bit => VN_data_out(10555),
        VN2CN2_bit => VN_data_out(10556),
        VN2CN3_bit => VN_data_out(10557),
        VN2CN4_bit => VN_data_out(10558),
        VN2CN5_bit => VN_data_out(10559),
        VN2CN0_sign => VN_sign_out(10554),
        VN2CN1_sign => VN_sign_out(10555),
        VN2CN2_sign => VN_sign_out(10556),
        VN2CN3_sign => VN_sign_out(10557),
        VN2CN4_sign => VN_sign_out(10558),
        VN2CN5_sign => VN_sign_out(10559),
        codeword => codeword(1759),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1760 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10565 downto 10560),
        Din0 => VN1760_in0,
        Din1 => VN1760_in1,
        Din2 => VN1760_in2,
        Din3 => VN1760_in3,
        Din4 => VN1760_in4,
        Din5 => VN1760_in5,
        VN2CN0_bit => VN_data_out(10560),
        VN2CN1_bit => VN_data_out(10561),
        VN2CN2_bit => VN_data_out(10562),
        VN2CN3_bit => VN_data_out(10563),
        VN2CN4_bit => VN_data_out(10564),
        VN2CN5_bit => VN_data_out(10565),
        VN2CN0_sign => VN_sign_out(10560),
        VN2CN1_sign => VN_sign_out(10561),
        VN2CN2_sign => VN_sign_out(10562),
        VN2CN3_sign => VN_sign_out(10563),
        VN2CN4_sign => VN_sign_out(10564),
        VN2CN5_sign => VN_sign_out(10565),
        codeword => codeword(1760),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1761 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10571 downto 10566),
        Din0 => VN1761_in0,
        Din1 => VN1761_in1,
        Din2 => VN1761_in2,
        Din3 => VN1761_in3,
        Din4 => VN1761_in4,
        Din5 => VN1761_in5,
        VN2CN0_bit => VN_data_out(10566),
        VN2CN1_bit => VN_data_out(10567),
        VN2CN2_bit => VN_data_out(10568),
        VN2CN3_bit => VN_data_out(10569),
        VN2CN4_bit => VN_data_out(10570),
        VN2CN5_bit => VN_data_out(10571),
        VN2CN0_sign => VN_sign_out(10566),
        VN2CN1_sign => VN_sign_out(10567),
        VN2CN2_sign => VN_sign_out(10568),
        VN2CN3_sign => VN_sign_out(10569),
        VN2CN4_sign => VN_sign_out(10570),
        VN2CN5_sign => VN_sign_out(10571),
        codeword => codeword(1761),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1762 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10577 downto 10572),
        Din0 => VN1762_in0,
        Din1 => VN1762_in1,
        Din2 => VN1762_in2,
        Din3 => VN1762_in3,
        Din4 => VN1762_in4,
        Din5 => VN1762_in5,
        VN2CN0_bit => VN_data_out(10572),
        VN2CN1_bit => VN_data_out(10573),
        VN2CN2_bit => VN_data_out(10574),
        VN2CN3_bit => VN_data_out(10575),
        VN2CN4_bit => VN_data_out(10576),
        VN2CN5_bit => VN_data_out(10577),
        VN2CN0_sign => VN_sign_out(10572),
        VN2CN1_sign => VN_sign_out(10573),
        VN2CN2_sign => VN_sign_out(10574),
        VN2CN3_sign => VN_sign_out(10575),
        VN2CN4_sign => VN_sign_out(10576),
        VN2CN5_sign => VN_sign_out(10577),
        codeword => codeword(1762),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1763 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10583 downto 10578),
        Din0 => VN1763_in0,
        Din1 => VN1763_in1,
        Din2 => VN1763_in2,
        Din3 => VN1763_in3,
        Din4 => VN1763_in4,
        Din5 => VN1763_in5,
        VN2CN0_bit => VN_data_out(10578),
        VN2CN1_bit => VN_data_out(10579),
        VN2CN2_bit => VN_data_out(10580),
        VN2CN3_bit => VN_data_out(10581),
        VN2CN4_bit => VN_data_out(10582),
        VN2CN5_bit => VN_data_out(10583),
        VN2CN0_sign => VN_sign_out(10578),
        VN2CN1_sign => VN_sign_out(10579),
        VN2CN2_sign => VN_sign_out(10580),
        VN2CN3_sign => VN_sign_out(10581),
        VN2CN4_sign => VN_sign_out(10582),
        VN2CN5_sign => VN_sign_out(10583),
        codeword => codeword(1763),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1764 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10589 downto 10584),
        Din0 => VN1764_in0,
        Din1 => VN1764_in1,
        Din2 => VN1764_in2,
        Din3 => VN1764_in3,
        Din4 => VN1764_in4,
        Din5 => VN1764_in5,
        VN2CN0_bit => VN_data_out(10584),
        VN2CN1_bit => VN_data_out(10585),
        VN2CN2_bit => VN_data_out(10586),
        VN2CN3_bit => VN_data_out(10587),
        VN2CN4_bit => VN_data_out(10588),
        VN2CN5_bit => VN_data_out(10589),
        VN2CN0_sign => VN_sign_out(10584),
        VN2CN1_sign => VN_sign_out(10585),
        VN2CN2_sign => VN_sign_out(10586),
        VN2CN3_sign => VN_sign_out(10587),
        VN2CN4_sign => VN_sign_out(10588),
        VN2CN5_sign => VN_sign_out(10589),
        codeword => codeword(1764),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1765 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10595 downto 10590),
        Din0 => VN1765_in0,
        Din1 => VN1765_in1,
        Din2 => VN1765_in2,
        Din3 => VN1765_in3,
        Din4 => VN1765_in4,
        Din5 => VN1765_in5,
        VN2CN0_bit => VN_data_out(10590),
        VN2CN1_bit => VN_data_out(10591),
        VN2CN2_bit => VN_data_out(10592),
        VN2CN3_bit => VN_data_out(10593),
        VN2CN4_bit => VN_data_out(10594),
        VN2CN5_bit => VN_data_out(10595),
        VN2CN0_sign => VN_sign_out(10590),
        VN2CN1_sign => VN_sign_out(10591),
        VN2CN2_sign => VN_sign_out(10592),
        VN2CN3_sign => VN_sign_out(10593),
        VN2CN4_sign => VN_sign_out(10594),
        VN2CN5_sign => VN_sign_out(10595),
        codeword => codeword(1765),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1766 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10601 downto 10596),
        Din0 => VN1766_in0,
        Din1 => VN1766_in1,
        Din2 => VN1766_in2,
        Din3 => VN1766_in3,
        Din4 => VN1766_in4,
        Din5 => VN1766_in5,
        VN2CN0_bit => VN_data_out(10596),
        VN2CN1_bit => VN_data_out(10597),
        VN2CN2_bit => VN_data_out(10598),
        VN2CN3_bit => VN_data_out(10599),
        VN2CN4_bit => VN_data_out(10600),
        VN2CN5_bit => VN_data_out(10601),
        VN2CN0_sign => VN_sign_out(10596),
        VN2CN1_sign => VN_sign_out(10597),
        VN2CN2_sign => VN_sign_out(10598),
        VN2CN3_sign => VN_sign_out(10599),
        VN2CN4_sign => VN_sign_out(10600),
        VN2CN5_sign => VN_sign_out(10601),
        codeword => codeword(1766),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1767 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10607 downto 10602),
        Din0 => VN1767_in0,
        Din1 => VN1767_in1,
        Din2 => VN1767_in2,
        Din3 => VN1767_in3,
        Din4 => VN1767_in4,
        Din5 => VN1767_in5,
        VN2CN0_bit => VN_data_out(10602),
        VN2CN1_bit => VN_data_out(10603),
        VN2CN2_bit => VN_data_out(10604),
        VN2CN3_bit => VN_data_out(10605),
        VN2CN4_bit => VN_data_out(10606),
        VN2CN5_bit => VN_data_out(10607),
        VN2CN0_sign => VN_sign_out(10602),
        VN2CN1_sign => VN_sign_out(10603),
        VN2CN2_sign => VN_sign_out(10604),
        VN2CN3_sign => VN_sign_out(10605),
        VN2CN4_sign => VN_sign_out(10606),
        VN2CN5_sign => VN_sign_out(10607),
        codeword => codeword(1767),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1768 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10613 downto 10608),
        Din0 => VN1768_in0,
        Din1 => VN1768_in1,
        Din2 => VN1768_in2,
        Din3 => VN1768_in3,
        Din4 => VN1768_in4,
        Din5 => VN1768_in5,
        VN2CN0_bit => VN_data_out(10608),
        VN2CN1_bit => VN_data_out(10609),
        VN2CN2_bit => VN_data_out(10610),
        VN2CN3_bit => VN_data_out(10611),
        VN2CN4_bit => VN_data_out(10612),
        VN2CN5_bit => VN_data_out(10613),
        VN2CN0_sign => VN_sign_out(10608),
        VN2CN1_sign => VN_sign_out(10609),
        VN2CN2_sign => VN_sign_out(10610),
        VN2CN3_sign => VN_sign_out(10611),
        VN2CN4_sign => VN_sign_out(10612),
        VN2CN5_sign => VN_sign_out(10613),
        codeword => codeword(1768),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1769 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10619 downto 10614),
        Din0 => VN1769_in0,
        Din1 => VN1769_in1,
        Din2 => VN1769_in2,
        Din3 => VN1769_in3,
        Din4 => VN1769_in4,
        Din5 => VN1769_in5,
        VN2CN0_bit => VN_data_out(10614),
        VN2CN1_bit => VN_data_out(10615),
        VN2CN2_bit => VN_data_out(10616),
        VN2CN3_bit => VN_data_out(10617),
        VN2CN4_bit => VN_data_out(10618),
        VN2CN5_bit => VN_data_out(10619),
        VN2CN0_sign => VN_sign_out(10614),
        VN2CN1_sign => VN_sign_out(10615),
        VN2CN2_sign => VN_sign_out(10616),
        VN2CN3_sign => VN_sign_out(10617),
        VN2CN4_sign => VN_sign_out(10618),
        VN2CN5_sign => VN_sign_out(10619),
        codeword => codeword(1769),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1770 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10625 downto 10620),
        Din0 => VN1770_in0,
        Din1 => VN1770_in1,
        Din2 => VN1770_in2,
        Din3 => VN1770_in3,
        Din4 => VN1770_in4,
        Din5 => VN1770_in5,
        VN2CN0_bit => VN_data_out(10620),
        VN2CN1_bit => VN_data_out(10621),
        VN2CN2_bit => VN_data_out(10622),
        VN2CN3_bit => VN_data_out(10623),
        VN2CN4_bit => VN_data_out(10624),
        VN2CN5_bit => VN_data_out(10625),
        VN2CN0_sign => VN_sign_out(10620),
        VN2CN1_sign => VN_sign_out(10621),
        VN2CN2_sign => VN_sign_out(10622),
        VN2CN3_sign => VN_sign_out(10623),
        VN2CN4_sign => VN_sign_out(10624),
        VN2CN5_sign => VN_sign_out(10625),
        codeword => codeword(1770),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1771 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10631 downto 10626),
        Din0 => VN1771_in0,
        Din1 => VN1771_in1,
        Din2 => VN1771_in2,
        Din3 => VN1771_in3,
        Din4 => VN1771_in4,
        Din5 => VN1771_in5,
        VN2CN0_bit => VN_data_out(10626),
        VN2CN1_bit => VN_data_out(10627),
        VN2CN2_bit => VN_data_out(10628),
        VN2CN3_bit => VN_data_out(10629),
        VN2CN4_bit => VN_data_out(10630),
        VN2CN5_bit => VN_data_out(10631),
        VN2CN0_sign => VN_sign_out(10626),
        VN2CN1_sign => VN_sign_out(10627),
        VN2CN2_sign => VN_sign_out(10628),
        VN2CN3_sign => VN_sign_out(10629),
        VN2CN4_sign => VN_sign_out(10630),
        VN2CN5_sign => VN_sign_out(10631),
        codeword => codeword(1771),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1772 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10637 downto 10632),
        Din0 => VN1772_in0,
        Din1 => VN1772_in1,
        Din2 => VN1772_in2,
        Din3 => VN1772_in3,
        Din4 => VN1772_in4,
        Din5 => VN1772_in5,
        VN2CN0_bit => VN_data_out(10632),
        VN2CN1_bit => VN_data_out(10633),
        VN2CN2_bit => VN_data_out(10634),
        VN2CN3_bit => VN_data_out(10635),
        VN2CN4_bit => VN_data_out(10636),
        VN2CN5_bit => VN_data_out(10637),
        VN2CN0_sign => VN_sign_out(10632),
        VN2CN1_sign => VN_sign_out(10633),
        VN2CN2_sign => VN_sign_out(10634),
        VN2CN3_sign => VN_sign_out(10635),
        VN2CN4_sign => VN_sign_out(10636),
        VN2CN5_sign => VN_sign_out(10637),
        codeword => codeword(1772),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1773 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10643 downto 10638),
        Din0 => VN1773_in0,
        Din1 => VN1773_in1,
        Din2 => VN1773_in2,
        Din3 => VN1773_in3,
        Din4 => VN1773_in4,
        Din5 => VN1773_in5,
        VN2CN0_bit => VN_data_out(10638),
        VN2CN1_bit => VN_data_out(10639),
        VN2CN2_bit => VN_data_out(10640),
        VN2CN3_bit => VN_data_out(10641),
        VN2CN4_bit => VN_data_out(10642),
        VN2CN5_bit => VN_data_out(10643),
        VN2CN0_sign => VN_sign_out(10638),
        VN2CN1_sign => VN_sign_out(10639),
        VN2CN2_sign => VN_sign_out(10640),
        VN2CN3_sign => VN_sign_out(10641),
        VN2CN4_sign => VN_sign_out(10642),
        VN2CN5_sign => VN_sign_out(10643),
        codeword => codeword(1773),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1774 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10649 downto 10644),
        Din0 => VN1774_in0,
        Din1 => VN1774_in1,
        Din2 => VN1774_in2,
        Din3 => VN1774_in3,
        Din4 => VN1774_in4,
        Din5 => VN1774_in5,
        VN2CN0_bit => VN_data_out(10644),
        VN2CN1_bit => VN_data_out(10645),
        VN2CN2_bit => VN_data_out(10646),
        VN2CN3_bit => VN_data_out(10647),
        VN2CN4_bit => VN_data_out(10648),
        VN2CN5_bit => VN_data_out(10649),
        VN2CN0_sign => VN_sign_out(10644),
        VN2CN1_sign => VN_sign_out(10645),
        VN2CN2_sign => VN_sign_out(10646),
        VN2CN3_sign => VN_sign_out(10647),
        VN2CN4_sign => VN_sign_out(10648),
        VN2CN5_sign => VN_sign_out(10649),
        codeword => codeword(1774),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1775 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10655 downto 10650),
        Din0 => VN1775_in0,
        Din1 => VN1775_in1,
        Din2 => VN1775_in2,
        Din3 => VN1775_in3,
        Din4 => VN1775_in4,
        Din5 => VN1775_in5,
        VN2CN0_bit => VN_data_out(10650),
        VN2CN1_bit => VN_data_out(10651),
        VN2CN2_bit => VN_data_out(10652),
        VN2CN3_bit => VN_data_out(10653),
        VN2CN4_bit => VN_data_out(10654),
        VN2CN5_bit => VN_data_out(10655),
        VN2CN0_sign => VN_sign_out(10650),
        VN2CN1_sign => VN_sign_out(10651),
        VN2CN2_sign => VN_sign_out(10652),
        VN2CN3_sign => VN_sign_out(10653),
        VN2CN4_sign => VN_sign_out(10654),
        VN2CN5_sign => VN_sign_out(10655),
        codeword => codeword(1775),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1776 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10661 downto 10656),
        Din0 => VN1776_in0,
        Din1 => VN1776_in1,
        Din2 => VN1776_in2,
        Din3 => VN1776_in3,
        Din4 => VN1776_in4,
        Din5 => VN1776_in5,
        VN2CN0_bit => VN_data_out(10656),
        VN2CN1_bit => VN_data_out(10657),
        VN2CN2_bit => VN_data_out(10658),
        VN2CN3_bit => VN_data_out(10659),
        VN2CN4_bit => VN_data_out(10660),
        VN2CN5_bit => VN_data_out(10661),
        VN2CN0_sign => VN_sign_out(10656),
        VN2CN1_sign => VN_sign_out(10657),
        VN2CN2_sign => VN_sign_out(10658),
        VN2CN3_sign => VN_sign_out(10659),
        VN2CN4_sign => VN_sign_out(10660),
        VN2CN5_sign => VN_sign_out(10661),
        codeword => codeword(1776),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1777 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10667 downto 10662),
        Din0 => VN1777_in0,
        Din1 => VN1777_in1,
        Din2 => VN1777_in2,
        Din3 => VN1777_in3,
        Din4 => VN1777_in4,
        Din5 => VN1777_in5,
        VN2CN0_bit => VN_data_out(10662),
        VN2CN1_bit => VN_data_out(10663),
        VN2CN2_bit => VN_data_out(10664),
        VN2CN3_bit => VN_data_out(10665),
        VN2CN4_bit => VN_data_out(10666),
        VN2CN5_bit => VN_data_out(10667),
        VN2CN0_sign => VN_sign_out(10662),
        VN2CN1_sign => VN_sign_out(10663),
        VN2CN2_sign => VN_sign_out(10664),
        VN2CN3_sign => VN_sign_out(10665),
        VN2CN4_sign => VN_sign_out(10666),
        VN2CN5_sign => VN_sign_out(10667),
        codeword => codeword(1777),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1778 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10673 downto 10668),
        Din0 => VN1778_in0,
        Din1 => VN1778_in1,
        Din2 => VN1778_in2,
        Din3 => VN1778_in3,
        Din4 => VN1778_in4,
        Din5 => VN1778_in5,
        VN2CN0_bit => VN_data_out(10668),
        VN2CN1_bit => VN_data_out(10669),
        VN2CN2_bit => VN_data_out(10670),
        VN2CN3_bit => VN_data_out(10671),
        VN2CN4_bit => VN_data_out(10672),
        VN2CN5_bit => VN_data_out(10673),
        VN2CN0_sign => VN_sign_out(10668),
        VN2CN1_sign => VN_sign_out(10669),
        VN2CN2_sign => VN_sign_out(10670),
        VN2CN3_sign => VN_sign_out(10671),
        VN2CN4_sign => VN_sign_out(10672),
        VN2CN5_sign => VN_sign_out(10673),
        codeword => codeword(1778),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1779 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10679 downto 10674),
        Din0 => VN1779_in0,
        Din1 => VN1779_in1,
        Din2 => VN1779_in2,
        Din3 => VN1779_in3,
        Din4 => VN1779_in4,
        Din5 => VN1779_in5,
        VN2CN0_bit => VN_data_out(10674),
        VN2CN1_bit => VN_data_out(10675),
        VN2CN2_bit => VN_data_out(10676),
        VN2CN3_bit => VN_data_out(10677),
        VN2CN4_bit => VN_data_out(10678),
        VN2CN5_bit => VN_data_out(10679),
        VN2CN0_sign => VN_sign_out(10674),
        VN2CN1_sign => VN_sign_out(10675),
        VN2CN2_sign => VN_sign_out(10676),
        VN2CN3_sign => VN_sign_out(10677),
        VN2CN4_sign => VN_sign_out(10678),
        VN2CN5_sign => VN_sign_out(10679),
        codeword => codeword(1779),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1780 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10685 downto 10680),
        Din0 => VN1780_in0,
        Din1 => VN1780_in1,
        Din2 => VN1780_in2,
        Din3 => VN1780_in3,
        Din4 => VN1780_in4,
        Din5 => VN1780_in5,
        VN2CN0_bit => VN_data_out(10680),
        VN2CN1_bit => VN_data_out(10681),
        VN2CN2_bit => VN_data_out(10682),
        VN2CN3_bit => VN_data_out(10683),
        VN2CN4_bit => VN_data_out(10684),
        VN2CN5_bit => VN_data_out(10685),
        VN2CN0_sign => VN_sign_out(10680),
        VN2CN1_sign => VN_sign_out(10681),
        VN2CN2_sign => VN_sign_out(10682),
        VN2CN3_sign => VN_sign_out(10683),
        VN2CN4_sign => VN_sign_out(10684),
        VN2CN5_sign => VN_sign_out(10685),
        codeword => codeword(1780),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1781 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10691 downto 10686),
        Din0 => VN1781_in0,
        Din1 => VN1781_in1,
        Din2 => VN1781_in2,
        Din3 => VN1781_in3,
        Din4 => VN1781_in4,
        Din5 => VN1781_in5,
        VN2CN0_bit => VN_data_out(10686),
        VN2CN1_bit => VN_data_out(10687),
        VN2CN2_bit => VN_data_out(10688),
        VN2CN3_bit => VN_data_out(10689),
        VN2CN4_bit => VN_data_out(10690),
        VN2CN5_bit => VN_data_out(10691),
        VN2CN0_sign => VN_sign_out(10686),
        VN2CN1_sign => VN_sign_out(10687),
        VN2CN2_sign => VN_sign_out(10688),
        VN2CN3_sign => VN_sign_out(10689),
        VN2CN4_sign => VN_sign_out(10690),
        VN2CN5_sign => VN_sign_out(10691),
        codeword => codeword(1781),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1782 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10697 downto 10692),
        Din0 => VN1782_in0,
        Din1 => VN1782_in1,
        Din2 => VN1782_in2,
        Din3 => VN1782_in3,
        Din4 => VN1782_in4,
        Din5 => VN1782_in5,
        VN2CN0_bit => VN_data_out(10692),
        VN2CN1_bit => VN_data_out(10693),
        VN2CN2_bit => VN_data_out(10694),
        VN2CN3_bit => VN_data_out(10695),
        VN2CN4_bit => VN_data_out(10696),
        VN2CN5_bit => VN_data_out(10697),
        VN2CN0_sign => VN_sign_out(10692),
        VN2CN1_sign => VN_sign_out(10693),
        VN2CN2_sign => VN_sign_out(10694),
        VN2CN3_sign => VN_sign_out(10695),
        VN2CN4_sign => VN_sign_out(10696),
        VN2CN5_sign => VN_sign_out(10697),
        codeword => codeword(1782),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1783 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10703 downto 10698),
        Din0 => VN1783_in0,
        Din1 => VN1783_in1,
        Din2 => VN1783_in2,
        Din3 => VN1783_in3,
        Din4 => VN1783_in4,
        Din5 => VN1783_in5,
        VN2CN0_bit => VN_data_out(10698),
        VN2CN1_bit => VN_data_out(10699),
        VN2CN2_bit => VN_data_out(10700),
        VN2CN3_bit => VN_data_out(10701),
        VN2CN4_bit => VN_data_out(10702),
        VN2CN5_bit => VN_data_out(10703),
        VN2CN0_sign => VN_sign_out(10698),
        VN2CN1_sign => VN_sign_out(10699),
        VN2CN2_sign => VN_sign_out(10700),
        VN2CN3_sign => VN_sign_out(10701),
        VN2CN4_sign => VN_sign_out(10702),
        VN2CN5_sign => VN_sign_out(10703),
        codeword => codeword(1783),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1784 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10709 downto 10704),
        Din0 => VN1784_in0,
        Din1 => VN1784_in1,
        Din2 => VN1784_in2,
        Din3 => VN1784_in3,
        Din4 => VN1784_in4,
        Din5 => VN1784_in5,
        VN2CN0_bit => VN_data_out(10704),
        VN2CN1_bit => VN_data_out(10705),
        VN2CN2_bit => VN_data_out(10706),
        VN2CN3_bit => VN_data_out(10707),
        VN2CN4_bit => VN_data_out(10708),
        VN2CN5_bit => VN_data_out(10709),
        VN2CN0_sign => VN_sign_out(10704),
        VN2CN1_sign => VN_sign_out(10705),
        VN2CN2_sign => VN_sign_out(10706),
        VN2CN3_sign => VN_sign_out(10707),
        VN2CN4_sign => VN_sign_out(10708),
        VN2CN5_sign => VN_sign_out(10709),
        codeword => codeword(1784),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1785 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10715 downto 10710),
        Din0 => VN1785_in0,
        Din1 => VN1785_in1,
        Din2 => VN1785_in2,
        Din3 => VN1785_in3,
        Din4 => VN1785_in4,
        Din5 => VN1785_in5,
        VN2CN0_bit => VN_data_out(10710),
        VN2CN1_bit => VN_data_out(10711),
        VN2CN2_bit => VN_data_out(10712),
        VN2CN3_bit => VN_data_out(10713),
        VN2CN4_bit => VN_data_out(10714),
        VN2CN5_bit => VN_data_out(10715),
        VN2CN0_sign => VN_sign_out(10710),
        VN2CN1_sign => VN_sign_out(10711),
        VN2CN2_sign => VN_sign_out(10712),
        VN2CN3_sign => VN_sign_out(10713),
        VN2CN4_sign => VN_sign_out(10714),
        VN2CN5_sign => VN_sign_out(10715),
        codeword => codeword(1785),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1786 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10721 downto 10716),
        Din0 => VN1786_in0,
        Din1 => VN1786_in1,
        Din2 => VN1786_in2,
        Din3 => VN1786_in3,
        Din4 => VN1786_in4,
        Din5 => VN1786_in5,
        VN2CN0_bit => VN_data_out(10716),
        VN2CN1_bit => VN_data_out(10717),
        VN2CN2_bit => VN_data_out(10718),
        VN2CN3_bit => VN_data_out(10719),
        VN2CN4_bit => VN_data_out(10720),
        VN2CN5_bit => VN_data_out(10721),
        VN2CN0_sign => VN_sign_out(10716),
        VN2CN1_sign => VN_sign_out(10717),
        VN2CN2_sign => VN_sign_out(10718),
        VN2CN3_sign => VN_sign_out(10719),
        VN2CN4_sign => VN_sign_out(10720),
        VN2CN5_sign => VN_sign_out(10721),
        codeword => codeword(1786),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1787 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10727 downto 10722),
        Din0 => VN1787_in0,
        Din1 => VN1787_in1,
        Din2 => VN1787_in2,
        Din3 => VN1787_in3,
        Din4 => VN1787_in4,
        Din5 => VN1787_in5,
        VN2CN0_bit => VN_data_out(10722),
        VN2CN1_bit => VN_data_out(10723),
        VN2CN2_bit => VN_data_out(10724),
        VN2CN3_bit => VN_data_out(10725),
        VN2CN4_bit => VN_data_out(10726),
        VN2CN5_bit => VN_data_out(10727),
        VN2CN0_sign => VN_sign_out(10722),
        VN2CN1_sign => VN_sign_out(10723),
        VN2CN2_sign => VN_sign_out(10724),
        VN2CN3_sign => VN_sign_out(10725),
        VN2CN4_sign => VN_sign_out(10726),
        VN2CN5_sign => VN_sign_out(10727),
        codeword => codeword(1787),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1788 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10733 downto 10728),
        Din0 => VN1788_in0,
        Din1 => VN1788_in1,
        Din2 => VN1788_in2,
        Din3 => VN1788_in3,
        Din4 => VN1788_in4,
        Din5 => VN1788_in5,
        VN2CN0_bit => VN_data_out(10728),
        VN2CN1_bit => VN_data_out(10729),
        VN2CN2_bit => VN_data_out(10730),
        VN2CN3_bit => VN_data_out(10731),
        VN2CN4_bit => VN_data_out(10732),
        VN2CN5_bit => VN_data_out(10733),
        VN2CN0_sign => VN_sign_out(10728),
        VN2CN1_sign => VN_sign_out(10729),
        VN2CN2_sign => VN_sign_out(10730),
        VN2CN3_sign => VN_sign_out(10731),
        VN2CN4_sign => VN_sign_out(10732),
        VN2CN5_sign => VN_sign_out(10733),
        codeword => codeword(1788),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1789 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10739 downto 10734),
        Din0 => VN1789_in0,
        Din1 => VN1789_in1,
        Din2 => VN1789_in2,
        Din3 => VN1789_in3,
        Din4 => VN1789_in4,
        Din5 => VN1789_in5,
        VN2CN0_bit => VN_data_out(10734),
        VN2CN1_bit => VN_data_out(10735),
        VN2CN2_bit => VN_data_out(10736),
        VN2CN3_bit => VN_data_out(10737),
        VN2CN4_bit => VN_data_out(10738),
        VN2CN5_bit => VN_data_out(10739),
        VN2CN0_sign => VN_sign_out(10734),
        VN2CN1_sign => VN_sign_out(10735),
        VN2CN2_sign => VN_sign_out(10736),
        VN2CN3_sign => VN_sign_out(10737),
        VN2CN4_sign => VN_sign_out(10738),
        VN2CN5_sign => VN_sign_out(10739),
        codeword => codeword(1789),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1790 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10745 downto 10740),
        Din0 => VN1790_in0,
        Din1 => VN1790_in1,
        Din2 => VN1790_in2,
        Din3 => VN1790_in3,
        Din4 => VN1790_in4,
        Din5 => VN1790_in5,
        VN2CN0_bit => VN_data_out(10740),
        VN2CN1_bit => VN_data_out(10741),
        VN2CN2_bit => VN_data_out(10742),
        VN2CN3_bit => VN_data_out(10743),
        VN2CN4_bit => VN_data_out(10744),
        VN2CN5_bit => VN_data_out(10745),
        VN2CN0_sign => VN_sign_out(10740),
        VN2CN1_sign => VN_sign_out(10741),
        VN2CN2_sign => VN_sign_out(10742),
        VN2CN3_sign => VN_sign_out(10743),
        VN2CN4_sign => VN_sign_out(10744),
        VN2CN5_sign => VN_sign_out(10745),
        codeword => codeword(1790),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1791 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10751 downto 10746),
        Din0 => VN1791_in0,
        Din1 => VN1791_in1,
        Din2 => VN1791_in2,
        Din3 => VN1791_in3,
        Din4 => VN1791_in4,
        Din5 => VN1791_in5,
        VN2CN0_bit => VN_data_out(10746),
        VN2CN1_bit => VN_data_out(10747),
        VN2CN2_bit => VN_data_out(10748),
        VN2CN3_bit => VN_data_out(10749),
        VN2CN4_bit => VN_data_out(10750),
        VN2CN5_bit => VN_data_out(10751),
        VN2CN0_sign => VN_sign_out(10746),
        VN2CN1_sign => VN_sign_out(10747),
        VN2CN2_sign => VN_sign_out(10748),
        VN2CN3_sign => VN_sign_out(10749),
        VN2CN4_sign => VN_sign_out(10750),
        VN2CN5_sign => VN_sign_out(10751),
        codeword => codeword(1791),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1792 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10757 downto 10752),
        Din0 => VN1792_in0,
        Din1 => VN1792_in1,
        Din2 => VN1792_in2,
        Din3 => VN1792_in3,
        Din4 => VN1792_in4,
        Din5 => VN1792_in5,
        VN2CN0_bit => VN_data_out(10752),
        VN2CN1_bit => VN_data_out(10753),
        VN2CN2_bit => VN_data_out(10754),
        VN2CN3_bit => VN_data_out(10755),
        VN2CN4_bit => VN_data_out(10756),
        VN2CN5_bit => VN_data_out(10757),
        VN2CN0_sign => VN_sign_out(10752),
        VN2CN1_sign => VN_sign_out(10753),
        VN2CN2_sign => VN_sign_out(10754),
        VN2CN3_sign => VN_sign_out(10755),
        VN2CN4_sign => VN_sign_out(10756),
        VN2CN5_sign => VN_sign_out(10757),
        codeword => codeword(1792),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1793 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10763 downto 10758),
        Din0 => VN1793_in0,
        Din1 => VN1793_in1,
        Din2 => VN1793_in2,
        Din3 => VN1793_in3,
        Din4 => VN1793_in4,
        Din5 => VN1793_in5,
        VN2CN0_bit => VN_data_out(10758),
        VN2CN1_bit => VN_data_out(10759),
        VN2CN2_bit => VN_data_out(10760),
        VN2CN3_bit => VN_data_out(10761),
        VN2CN4_bit => VN_data_out(10762),
        VN2CN5_bit => VN_data_out(10763),
        VN2CN0_sign => VN_sign_out(10758),
        VN2CN1_sign => VN_sign_out(10759),
        VN2CN2_sign => VN_sign_out(10760),
        VN2CN3_sign => VN_sign_out(10761),
        VN2CN4_sign => VN_sign_out(10762),
        VN2CN5_sign => VN_sign_out(10763),
        codeword => codeword(1793),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1794 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10769 downto 10764),
        Din0 => VN1794_in0,
        Din1 => VN1794_in1,
        Din2 => VN1794_in2,
        Din3 => VN1794_in3,
        Din4 => VN1794_in4,
        Din5 => VN1794_in5,
        VN2CN0_bit => VN_data_out(10764),
        VN2CN1_bit => VN_data_out(10765),
        VN2CN2_bit => VN_data_out(10766),
        VN2CN3_bit => VN_data_out(10767),
        VN2CN4_bit => VN_data_out(10768),
        VN2CN5_bit => VN_data_out(10769),
        VN2CN0_sign => VN_sign_out(10764),
        VN2CN1_sign => VN_sign_out(10765),
        VN2CN2_sign => VN_sign_out(10766),
        VN2CN3_sign => VN_sign_out(10767),
        VN2CN4_sign => VN_sign_out(10768),
        VN2CN5_sign => VN_sign_out(10769),
        codeword => codeword(1794),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1795 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10775 downto 10770),
        Din0 => VN1795_in0,
        Din1 => VN1795_in1,
        Din2 => VN1795_in2,
        Din3 => VN1795_in3,
        Din4 => VN1795_in4,
        Din5 => VN1795_in5,
        VN2CN0_bit => VN_data_out(10770),
        VN2CN1_bit => VN_data_out(10771),
        VN2CN2_bit => VN_data_out(10772),
        VN2CN3_bit => VN_data_out(10773),
        VN2CN4_bit => VN_data_out(10774),
        VN2CN5_bit => VN_data_out(10775),
        VN2CN0_sign => VN_sign_out(10770),
        VN2CN1_sign => VN_sign_out(10771),
        VN2CN2_sign => VN_sign_out(10772),
        VN2CN3_sign => VN_sign_out(10773),
        VN2CN4_sign => VN_sign_out(10774),
        VN2CN5_sign => VN_sign_out(10775),
        codeword => codeword(1795),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1796 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10781 downto 10776),
        Din0 => VN1796_in0,
        Din1 => VN1796_in1,
        Din2 => VN1796_in2,
        Din3 => VN1796_in3,
        Din4 => VN1796_in4,
        Din5 => VN1796_in5,
        VN2CN0_bit => VN_data_out(10776),
        VN2CN1_bit => VN_data_out(10777),
        VN2CN2_bit => VN_data_out(10778),
        VN2CN3_bit => VN_data_out(10779),
        VN2CN4_bit => VN_data_out(10780),
        VN2CN5_bit => VN_data_out(10781),
        VN2CN0_sign => VN_sign_out(10776),
        VN2CN1_sign => VN_sign_out(10777),
        VN2CN2_sign => VN_sign_out(10778),
        VN2CN3_sign => VN_sign_out(10779),
        VN2CN4_sign => VN_sign_out(10780),
        VN2CN5_sign => VN_sign_out(10781),
        codeword => codeword(1796),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1797 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10787 downto 10782),
        Din0 => VN1797_in0,
        Din1 => VN1797_in1,
        Din2 => VN1797_in2,
        Din3 => VN1797_in3,
        Din4 => VN1797_in4,
        Din5 => VN1797_in5,
        VN2CN0_bit => VN_data_out(10782),
        VN2CN1_bit => VN_data_out(10783),
        VN2CN2_bit => VN_data_out(10784),
        VN2CN3_bit => VN_data_out(10785),
        VN2CN4_bit => VN_data_out(10786),
        VN2CN5_bit => VN_data_out(10787),
        VN2CN0_sign => VN_sign_out(10782),
        VN2CN1_sign => VN_sign_out(10783),
        VN2CN2_sign => VN_sign_out(10784),
        VN2CN3_sign => VN_sign_out(10785),
        VN2CN4_sign => VN_sign_out(10786),
        VN2CN5_sign => VN_sign_out(10787),
        codeword => codeword(1797),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1798 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10793 downto 10788),
        Din0 => VN1798_in0,
        Din1 => VN1798_in1,
        Din2 => VN1798_in2,
        Din3 => VN1798_in3,
        Din4 => VN1798_in4,
        Din5 => VN1798_in5,
        VN2CN0_bit => VN_data_out(10788),
        VN2CN1_bit => VN_data_out(10789),
        VN2CN2_bit => VN_data_out(10790),
        VN2CN3_bit => VN_data_out(10791),
        VN2CN4_bit => VN_data_out(10792),
        VN2CN5_bit => VN_data_out(10793),
        VN2CN0_sign => VN_sign_out(10788),
        VN2CN1_sign => VN_sign_out(10789),
        VN2CN2_sign => VN_sign_out(10790),
        VN2CN3_sign => VN_sign_out(10791),
        VN2CN4_sign => VN_sign_out(10792),
        VN2CN5_sign => VN_sign_out(10793),
        codeword => codeword(1798),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1799 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10799 downto 10794),
        Din0 => VN1799_in0,
        Din1 => VN1799_in1,
        Din2 => VN1799_in2,
        Din3 => VN1799_in3,
        Din4 => VN1799_in4,
        Din5 => VN1799_in5,
        VN2CN0_bit => VN_data_out(10794),
        VN2CN1_bit => VN_data_out(10795),
        VN2CN2_bit => VN_data_out(10796),
        VN2CN3_bit => VN_data_out(10797),
        VN2CN4_bit => VN_data_out(10798),
        VN2CN5_bit => VN_data_out(10799),
        VN2CN0_sign => VN_sign_out(10794),
        VN2CN1_sign => VN_sign_out(10795),
        VN2CN2_sign => VN_sign_out(10796),
        VN2CN3_sign => VN_sign_out(10797),
        VN2CN4_sign => VN_sign_out(10798),
        VN2CN5_sign => VN_sign_out(10799),
        codeword => codeword(1799),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1800 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10805 downto 10800),
        Din0 => VN1800_in0,
        Din1 => VN1800_in1,
        Din2 => VN1800_in2,
        Din3 => VN1800_in3,
        Din4 => VN1800_in4,
        Din5 => VN1800_in5,
        VN2CN0_bit => VN_data_out(10800),
        VN2CN1_bit => VN_data_out(10801),
        VN2CN2_bit => VN_data_out(10802),
        VN2CN3_bit => VN_data_out(10803),
        VN2CN4_bit => VN_data_out(10804),
        VN2CN5_bit => VN_data_out(10805),
        VN2CN0_sign => VN_sign_out(10800),
        VN2CN1_sign => VN_sign_out(10801),
        VN2CN2_sign => VN_sign_out(10802),
        VN2CN3_sign => VN_sign_out(10803),
        VN2CN4_sign => VN_sign_out(10804),
        VN2CN5_sign => VN_sign_out(10805),
        codeword => codeword(1800),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1801 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10811 downto 10806),
        Din0 => VN1801_in0,
        Din1 => VN1801_in1,
        Din2 => VN1801_in2,
        Din3 => VN1801_in3,
        Din4 => VN1801_in4,
        Din5 => VN1801_in5,
        VN2CN0_bit => VN_data_out(10806),
        VN2CN1_bit => VN_data_out(10807),
        VN2CN2_bit => VN_data_out(10808),
        VN2CN3_bit => VN_data_out(10809),
        VN2CN4_bit => VN_data_out(10810),
        VN2CN5_bit => VN_data_out(10811),
        VN2CN0_sign => VN_sign_out(10806),
        VN2CN1_sign => VN_sign_out(10807),
        VN2CN2_sign => VN_sign_out(10808),
        VN2CN3_sign => VN_sign_out(10809),
        VN2CN4_sign => VN_sign_out(10810),
        VN2CN5_sign => VN_sign_out(10811),
        codeword => codeword(1801),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1802 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10817 downto 10812),
        Din0 => VN1802_in0,
        Din1 => VN1802_in1,
        Din2 => VN1802_in2,
        Din3 => VN1802_in3,
        Din4 => VN1802_in4,
        Din5 => VN1802_in5,
        VN2CN0_bit => VN_data_out(10812),
        VN2CN1_bit => VN_data_out(10813),
        VN2CN2_bit => VN_data_out(10814),
        VN2CN3_bit => VN_data_out(10815),
        VN2CN4_bit => VN_data_out(10816),
        VN2CN5_bit => VN_data_out(10817),
        VN2CN0_sign => VN_sign_out(10812),
        VN2CN1_sign => VN_sign_out(10813),
        VN2CN2_sign => VN_sign_out(10814),
        VN2CN3_sign => VN_sign_out(10815),
        VN2CN4_sign => VN_sign_out(10816),
        VN2CN5_sign => VN_sign_out(10817),
        codeword => codeword(1802),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1803 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10823 downto 10818),
        Din0 => VN1803_in0,
        Din1 => VN1803_in1,
        Din2 => VN1803_in2,
        Din3 => VN1803_in3,
        Din4 => VN1803_in4,
        Din5 => VN1803_in5,
        VN2CN0_bit => VN_data_out(10818),
        VN2CN1_bit => VN_data_out(10819),
        VN2CN2_bit => VN_data_out(10820),
        VN2CN3_bit => VN_data_out(10821),
        VN2CN4_bit => VN_data_out(10822),
        VN2CN5_bit => VN_data_out(10823),
        VN2CN0_sign => VN_sign_out(10818),
        VN2CN1_sign => VN_sign_out(10819),
        VN2CN2_sign => VN_sign_out(10820),
        VN2CN3_sign => VN_sign_out(10821),
        VN2CN4_sign => VN_sign_out(10822),
        VN2CN5_sign => VN_sign_out(10823),
        codeword => codeword(1803),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1804 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10829 downto 10824),
        Din0 => VN1804_in0,
        Din1 => VN1804_in1,
        Din2 => VN1804_in2,
        Din3 => VN1804_in3,
        Din4 => VN1804_in4,
        Din5 => VN1804_in5,
        VN2CN0_bit => VN_data_out(10824),
        VN2CN1_bit => VN_data_out(10825),
        VN2CN2_bit => VN_data_out(10826),
        VN2CN3_bit => VN_data_out(10827),
        VN2CN4_bit => VN_data_out(10828),
        VN2CN5_bit => VN_data_out(10829),
        VN2CN0_sign => VN_sign_out(10824),
        VN2CN1_sign => VN_sign_out(10825),
        VN2CN2_sign => VN_sign_out(10826),
        VN2CN3_sign => VN_sign_out(10827),
        VN2CN4_sign => VN_sign_out(10828),
        VN2CN5_sign => VN_sign_out(10829),
        codeword => codeword(1804),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1805 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10835 downto 10830),
        Din0 => VN1805_in0,
        Din1 => VN1805_in1,
        Din2 => VN1805_in2,
        Din3 => VN1805_in3,
        Din4 => VN1805_in4,
        Din5 => VN1805_in5,
        VN2CN0_bit => VN_data_out(10830),
        VN2CN1_bit => VN_data_out(10831),
        VN2CN2_bit => VN_data_out(10832),
        VN2CN3_bit => VN_data_out(10833),
        VN2CN4_bit => VN_data_out(10834),
        VN2CN5_bit => VN_data_out(10835),
        VN2CN0_sign => VN_sign_out(10830),
        VN2CN1_sign => VN_sign_out(10831),
        VN2CN2_sign => VN_sign_out(10832),
        VN2CN3_sign => VN_sign_out(10833),
        VN2CN4_sign => VN_sign_out(10834),
        VN2CN5_sign => VN_sign_out(10835),
        codeword => codeword(1805),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1806 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10841 downto 10836),
        Din0 => VN1806_in0,
        Din1 => VN1806_in1,
        Din2 => VN1806_in2,
        Din3 => VN1806_in3,
        Din4 => VN1806_in4,
        Din5 => VN1806_in5,
        VN2CN0_bit => VN_data_out(10836),
        VN2CN1_bit => VN_data_out(10837),
        VN2CN2_bit => VN_data_out(10838),
        VN2CN3_bit => VN_data_out(10839),
        VN2CN4_bit => VN_data_out(10840),
        VN2CN5_bit => VN_data_out(10841),
        VN2CN0_sign => VN_sign_out(10836),
        VN2CN1_sign => VN_sign_out(10837),
        VN2CN2_sign => VN_sign_out(10838),
        VN2CN3_sign => VN_sign_out(10839),
        VN2CN4_sign => VN_sign_out(10840),
        VN2CN5_sign => VN_sign_out(10841),
        codeword => codeword(1806),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1807 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10847 downto 10842),
        Din0 => VN1807_in0,
        Din1 => VN1807_in1,
        Din2 => VN1807_in2,
        Din3 => VN1807_in3,
        Din4 => VN1807_in4,
        Din5 => VN1807_in5,
        VN2CN0_bit => VN_data_out(10842),
        VN2CN1_bit => VN_data_out(10843),
        VN2CN2_bit => VN_data_out(10844),
        VN2CN3_bit => VN_data_out(10845),
        VN2CN4_bit => VN_data_out(10846),
        VN2CN5_bit => VN_data_out(10847),
        VN2CN0_sign => VN_sign_out(10842),
        VN2CN1_sign => VN_sign_out(10843),
        VN2CN2_sign => VN_sign_out(10844),
        VN2CN3_sign => VN_sign_out(10845),
        VN2CN4_sign => VN_sign_out(10846),
        VN2CN5_sign => VN_sign_out(10847),
        codeword => codeword(1807),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1808 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10853 downto 10848),
        Din0 => VN1808_in0,
        Din1 => VN1808_in1,
        Din2 => VN1808_in2,
        Din3 => VN1808_in3,
        Din4 => VN1808_in4,
        Din5 => VN1808_in5,
        VN2CN0_bit => VN_data_out(10848),
        VN2CN1_bit => VN_data_out(10849),
        VN2CN2_bit => VN_data_out(10850),
        VN2CN3_bit => VN_data_out(10851),
        VN2CN4_bit => VN_data_out(10852),
        VN2CN5_bit => VN_data_out(10853),
        VN2CN0_sign => VN_sign_out(10848),
        VN2CN1_sign => VN_sign_out(10849),
        VN2CN2_sign => VN_sign_out(10850),
        VN2CN3_sign => VN_sign_out(10851),
        VN2CN4_sign => VN_sign_out(10852),
        VN2CN5_sign => VN_sign_out(10853),
        codeword => codeword(1808),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1809 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10859 downto 10854),
        Din0 => VN1809_in0,
        Din1 => VN1809_in1,
        Din2 => VN1809_in2,
        Din3 => VN1809_in3,
        Din4 => VN1809_in4,
        Din5 => VN1809_in5,
        VN2CN0_bit => VN_data_out(10854),
        VN2CN1_bit => VN_data_out(10855),
        VN2CN2_bit => VN_data_out(10856),
        VN2CN3_bit => VN_data_out(10857),
        VN2CN4_bit => VN_data_out(10858),
        VN2CN5_bit => VN_data_out(10859),
        VN2CN0_sign => VN_sign_out(10854),
        VN2CN1_sign => VN_sign_out(10855),
        VN2CN2_sign => VN_sign_out(10856),
        VN2CN3_sign => VN_sign_out(10857),
        VN2CN4_sign => VN_sign_out(10858),
        VN2CN5_sign => VN_sign_out(10859),
        codeword => codeword(1809),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1810 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10865 downto 10860),
        Din0 => VN1810_in0,
        Din1 => VN1810_in1,
        Din2 => VN1810_in2,
        Din3 => VN1810_in3,
        Din4 => VN1810_in4,
        Din5 => VN1810_in5,
        VN2CN0_bit => VN_data_out(10860),
        VN2CN1_bit => VN_data_out(10861),
        VN2CN2_bit => VN_data_out(10862),
        VN2CN3_bit => VN_data_out(10863),
        VN2CN4_bit => VN_data_out(10864),
        VN2CN5_bit => VN_data_out(10865),
        VN2CN0_sign => VN_sign_out(10860),
        VN2CN1_sign => VN_sign_out(10861),
        VN2CN2_sign => VN_sign_out(10862),
        VN2CN3_sign => VN_sign_out(10863),
        VN2CN4_sign => VN_sign_out(10864),
        VN2CN5_sign => VN_sign_out(10865),
        codeword => codeword(1810),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1811 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10871 downto 10866),
        Din0 => VN1811_in0,
        Din1 => VN1811_in1,
        Din2 => VN1811_in2,
        Din3 => VN1811_in3,
        Din4 => VN1811_in4,
        Din5 => VN1811_in5,
        VN2CN0_bit => VN_data_out(10866),
        VN2CN1_bit => VN_data_out(10867),
        VN2CN2_bit => VN_data_out(10868),
        VN2CN3_bit => VN_data_out(10869),
        VN2CN4_bit => VN_data_out(10870),
        VN2CN5_bit => VN_data_out(10871),
        VN2CN0_sign => VN_sign_out(10866),
        VN2CN1_sign => VN_sign_out(10867),
        VN2CN2_sign => VN_sign_out(10868),
        VN2CN3_sign => VN_sign_out(10869),
        VN2CN4_sign => VN_sign_out(10870),
        VN2CN5_sign => VN_sign_out(10871),
        codeword => codeword(1811),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1812 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10877 downto 10872),
        Din0 => VN1812_in0,
        Din1 => VN1812_in1,
        Din2 => VN1812_in2,
        Din3 => VN1812_in3,
        Din4 => VN1812_in4,
        Din5 => VN1812_in5,
        VN2CN0_bit => VN_data_out(10872),
        VN2CN1_bit => VN_data_out(10873),
        VN2CN2_bit => VN_data_out(10874),
        VN2CN3_bit => VN_data_out(10875),
        VN2CN4_bit => VN_data_out(10876),
        VN2CN5_bit => VN_data_out(10877),
        VN2CN0_sign => VN_sign_out(10872),
        VN2CN1_sign => VN_sign_out(10873),
        VN2CN2_sign => VN_sign_out(10874),
        VN2CN3_sign => VN_sign_out(10875),
        VN2CN4_sign => VN_sign_out(10876),
        VN2CN5_sign => VN_sign_out(10877),
        codeword => codeword(1812),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1813 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10883 downto 10878),
        Din0 => VN1813_in0,
        Din1 => VN1813_in1,
        Din2 => VN1813_in2,
        Din3 => VN1813_in3,
        Din4 => VN1813_in4,
        Din5 => VN1813_in5,
        VN2CN0_bit => VN_data_out(10878),
        VN2CN1_bit => VN_data_out(10879),
        VN2CN2_bit => VN_data_out(10880),
        VN2CN3_bit => VN_data_out(10881),
        VN2CN4_bit => VN_data_out(10882),
        VN2CN5_bit => VN_data_out(10883),
        VN2CN0_sign => VN_sign_out(10878),
        VN2CN1_sign => VN_sign_out(10879),
        VN2CN2_sign => VN_sign_out(10880),
        VN2CN3_sign => VN_sign_out(10881),
        VN2CN4_sign => VN_sign_out(10882),
        VN2CN5_sign => VN_sign_out(10883),
        codeword => codeword(1813),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1814 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10889 downto 10884),
        Din0 => VN1814_in0,
        Din1 => VN1814_in1,
        Din2 => VN1814_in2,
        Din3 => VN1814_in3,
        Din4 => VN1814_in4,
        Din5 => VN1814_in5,
        VN2CN0_bit => VN_data_out(10884),
        VN2CN1_bit => VN_data_out(10885),
        VN2CN2_bit => VN_data_out(10886),
        VN2CN3_bit => VN_data_out(10887),
        VN2CN4_bit => VN_data_out(10888),
        VN2CN5_bit => VN_data_out(10889),
        VN2CN0_sign => VN_sign_out(10884),
        VN2CN1_sign => VN_sign_out(10885),
        VN2CN2_sign => VN_sign_out(10886),
        VN2CN3_sign => VN_sign_out(10887),
        VN2CN4_sign => VN_sign_out(10888),
        VN2CN5_sign => VN_sign_out(10889),
        codeword => codeword(1814),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1815 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10895 downto 10890),
        Din0 => VN1815_in0,
        Din1 => VN1815_in1,
        Din2 => VN1815_in2,
        Din3 => VN1815_in3,
        Din4 => VN1815_in4,
        Din5 => VN1815_in5,
        VN2CN0_bit => VN_data_out(10890),
        VN2CN1_bit => VN_data_out(10891),
        VN2CN2_bit => VN_data_out(10892),
        VN2CN3_bit => VN_data_out(10893),
        VN2CN4_bit => VN_data_out(10894),
        VN2CN5_bit => VN_data_out(10895),
        VN2CN0_sign => VN_sign_out(10890),
        VN2CN1_sign => VN_sign_out(10891),
        VN2CN2_sign => VN_sign_out(10892),
        VN2CN3_sign => VN_sign_out(10893),
        VN2CN4_sign => VN_sign_out(10894),
        VN2CN5_sign => VN_sign_out(10895),
        codeword => codeword(1815),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1816 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10901 downto 10896),
        Din0 => VN1816_in0,
        Din1 => VN1816_in1,
        Din2 => VN1816_in2,
        Din3 => VN1816_in3,
        Din4 => VN1816_in4,
        Din5 => VN1816_in5,
        VN2CN0_bit => VN_data_out(10896),
        VN2CN1_bit => VN_data_out(10897),
        VN2CN2_bit => VN_data_out(10898),
        VN2CN3_bit => VN_data_out(10899),
        VN2CN4_bit => VN_data_out(10900),
        VN2CN5_bit => VN_data_out(10901),
        VN2CN0_sign => VN_sign_out(10896),
        VN2CN1_sign => VN_sign_out(10897),
        VN2CN2_sign => VN_sign_out(10898),
        VN2CN3_sign => VN_sign_out(10899),
        VN2CN4_sign => VN_sign_out(10900),
        VN2CN5_sign => VN_sign_out(10901),
        codeword => codeword(1816),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1817 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10907 downto 10902),
        Din0 => VN1817_in0,
        Din1 => VN1817_in1,
        Din2 => VN1817_in2,
        Din3 => VN1817_in3,
        Din4 => VN1817_in4,
        Din5 => VN1817_in5,
        VN2CN0_bit => VN_data_out(10902),
        VN2CN1_bit => VN_data_out(10903),
        VN2CN2_bit => VN_data_out(10904),
        VN2CN3_bit => VN_data_out(10905),
        VN2CN4_bit => VN_data_out(10906),
        VN2CN5_bit => VN_data_out(10907),
        VN2CN0_sign => VN_sign_out(10902),
        VN2CN1_sign => VN_sign_out(10903),
        VN2CN2_sign => VN_sign_out(10904),
        VN2CN3_sign => VN_sign_out(10905),
        VN2CN4_sign => VN_sign_out(10906),
        VN2CN5_sign => VN_sign_out(10907),
        codeword => codeword(1817),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1818 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10913 downto 10908),
        Din0 => VN1818_in0,
        Din1 => VN1818_in1,
        Din2 => VN1818_in2,
        Din3 => VN1818_in3,
        Din4 => VN1818_in4,
        Din5 => VN1818_in5,
        VN2CN0_bit => VN_data_out(10908),
        VN2CN1_bit => VN_data_out(10909),
        VN2CN2_bit => VN_data_out(10910),
        VN2CN3_bit => VN_data_out(10911),
        VN2CN4_bit => VN_data_out(10912),
        VN2CN5_bit => VN_data_out(10913),
        VN2CN0_sign => VN_sign_out(10908),
        VN2CN1_sign => VN_sign_out(10909),
        VN2CN2_sign => VN_sign_out(10910),
        VN2CN3_sign => VN_sign_out(10911),
        VN2CN4_sign => VN_sign_out(10912),
        VN2CN5_sign => VN_sign_out(10913),
        codeword => codeword(1818),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1819 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10919 downto 10914),
        Din0 => VN1819_in0,
        Din1 => VN1819_in1,
        Din2 => VN1819_in2,
        Din3 => VN1819_in3,
        Din4 => VN1819_in4,
        Din5 => VN1819_in5,
        VN2CN0_bit => VN_data_out(10914),
        VN2CN1_bit => VN_data_out(10915),
        VN2CN2_bit => VN_data_out(10916),
        VN2CN3_bit => VN_data_out(10917),
        VN2CN4_bit => VN_data_out(10918),
        VN2CN5_bit => VN_data_out(10919),
        VN2CN0_sign => VN_sign_out(10914),
        VN2CN1_sign => VN_sign_out(10915),
        VN2CN2_sign => VN_sign_out(10916),
        VN2CN3_sign => VN_sign_out(10917),
        VN2CN4_sign => VN_sign_out(10918),
        VN2CN5_sign => VN_sign_out(10919),
        codeword => codeword(1819),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1820 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10925 downto 10920),
        Din0 => VN1820_in0,
        Din1 => VN1820_in1,
        Din2 => VN1820_in2,
        Din3 => VN1820_in3,
        Din4 => VN1820_in4,
        Din5 => VN1820_in5,
        VN2CN0_bit => VN_data_out(10920),
        VN2CN1_bit => VN_data_out(10921),
        VN2CN2_bit => VN_data_out(10922),
        VN2CN3_bit => VN_data_out(10923),
        VN2CN4_bit => VN_data_out(10924),
        VN2CN5_bit => VN_data_out(10925),
        VN2CN0_sign => VN_sign_out(10920),
        VN2CN1_sign => VN_sign_out(10921),
        VN2CN2_sign => VN_sign_out(10922),
        VN2CN3_sign => VN_sign_out(10923),
        VN2CN4_sign => VN_sign_out(10924),
        VN2CN5_sign => VN_sign_out(10925),
        codeword => codeword(1820),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1821 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10931 downto 10926),
        Din0 => VN1821_in0,
        Din1 => VN1821_in1,
        Din2 => VN1821_in2,
        Din3 => VN1821_in3,
        Din4 => VN1821_in4,
        Din5 => VN1821_in5,
        VN2CN0_bit => VN_data_out(10926),
        VN2CN1_bit => VN_data_out(10927),
        VN2CN2_bit => VN_data_out(10928),
        VN2CN3_bit => VN_data_out(10929),
        VN2CN4_bit => VN_data_out(10930),
        VN2CN5_bit => VN_data_out(10931),
        VN2CN0_sign => VN_sign_out(10926),
        VN2CN1_sign => VN_sign_out(10927),
        VN2CN2_sign => VN_sign_out(10928),
        VN2CN3_sign => VN_sign_out(10929),
        VN2CN4_sign => VN_sign_out(10930),
        VN2CN5_sign => VN_sign_out(10931),
        codeword => codeword(1821),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1822 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10937 downto 10932),
        Din0 => VN1822_in0,
        Din1 => VN1822_in1,
        Din2 => VN1822_in2,
        Din3 => VN1822_in3,
        Din4 => VN1822_in4,
        Din5 => VN1822_in5,
        VN2CN0_bit => VN_data_out(10932),
        VN2CN1_bit => VN_data_out(10933),
        VN2CN2_bit => VN_data_out(10934),
        VN2CN3_bit => VN_data_out(10935),
        VN2CN4_bit => VN_data_out(10936),
        VN2CN5_bit => VN_data_out(10937),
        VN2CN0_sign => VN_sign_out(10932),
        VN2CN1_sign => VN_sign_out(10933),
        VN2CN2_sign => VN_sign_out(10934),
        VN2CN3_sign => VN_sign_out(10935),
        VN2CN4_sign => VN_sign_out(10936),
        VN2CN5_sign => VN_sign_out(10937),
        codeword => codeword(1822),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1823 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10943 downto 10938),
        Din0 => VN1823_in0,
        Din1 => VN1823_in1,
        Din2 => VN1823_in2,
        Din3 => VN1823_in3,
        Din4 => VN1823_in4,
        Din5 => VN1823_in5,
        VN2CN0_bit => VN_data_out(10938),
        VN2CN1_bit => VN_data_out(10939),
        VN2CN2_bit => VN_data_out(10940),
        VN2CN3_bit => VN_data_out(10941),
        VN2CN4_bit => VN_data_out(10942),
        VN2CN5_bit => VN_data_out(10943),
        VN2CN0_sign => VN_sign_out(10938),
        VN2CN1_sign => VN_sign_out(10939),
        VN2CN2_sign => VN_sign_out(10940),
        VN2CN3_sign => VN_sign_out(10941),
        VN2CN4_sign => VN_sign_out(10942),
        VN2CN5_sign => VN_sign_out(10943),
        codeword => codeword(1823),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1824 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10949 downto 10944),
        Din0 => VN1824_in0,
        Din1 => VN1824_in1,
        Din2 => VN1824_in2,
        Din3 => VN1824_in3,
        Din4 => VN1824_in4,
        Din5 => VN1824_in5,
        VN2CN0_bit => VN_data_out(10944),
        VN2CN1_bit => VN_data_out(10945),
        VN2CN2_bit => VN_data_out(10946),
        VN2CN3_bit => VN_data_out(10947),
        VN2CN4_bit => VN_data_out(10948),
        VN2CN5_bit => VN_data_out(10949),
        VN2CN0_sign => VN_sign_out(10944),
        VN2CN1_sign => VN_sign_out(10945),
        VN2CN2_sign => VN_sign_out(10946),
        VN2CN3_sign => VN_sign_out(10947),
        VN2CN4_sign => VN_sign_out(10948),
        VN2CN5_sign => VN_sign_out(10949),
        codeword => codeword(1824),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1825 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10955 downto 10950),
        Din0 => VN1825_in0,
        Din1 => VN1825_in1,
        Din2 => VN1825_in2,
        Din3 => VN1825_in3,
        Din4 => VN1825_in4,
        Din5 => VN1825_in5,
        VN2CN0_bit => VN_data_out(10950),
        VN2CN1_bit => VN_data_out(10951),
        VN2CN2_bit => VN_data_out(10952),
        VN2CN3_bit => VN_data_out(10953),
        VN2CN4_bit => VN_data_out(10954),
        VN2CN5_bit => VN_data_out(10955),
        VN2CN0_sign => VN_sign_out(10950),
        VN2CN1_sign => VN_sign_out(10951),
        VN2CN2_sign => VN_sign_out(10952),
        VN2CN3_sign => VN_sign_out(10953),
        VN2CN4_sign => VN_sign_out(10954),
        VN2CN5_sign => VN_sign_out(10955),
        codeword => codeword(1825),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1826 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10961 downto 10956),
        Din0 => VN1826_in0,
        Din1 => VN1826_in1,
        Din2 => VN1826_in2,
        Din3 => VN1826_in3,
        Din4 => VN1826_in4,
        Din5 => VN1826_in5,
        VN2CN0_bit => VN_data_out(10956),
        VN2CN1_bit => VN_data_out(10957),
        VN2CN2_bit => VN_data_out(10958),
        VN2CN3_bit => VN_data_out(10959),
        VN2CN4_bit => VN_data_out(10960),
        VN2CN5_bit => VN_data_out(10961),
        VN2CN0_sign => VN_sign_out(10956),
        VN2CN1_sign => VN_sign_out(10957),
        VN2CN2_sign => VN_sign_out(10958),
        VN2CN3_sign => VN_sign_out(10959),
        VN2CN4_sign => VN_sign_out(10960),
        VN2CN5_sign => VN_sign_out(10961),
        codeword => codeword(1826),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1827 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10967 downto 10962),
        Din0 => VN1827_in0,
        Din1 => VN1827_in1,
        Din2 => VN1827_in2,
        Din3 => VN1827_in3,
        Din4 => VN1827_in4,
        Din5 => VN1827_in5,
        VN2CN0_bit => VN_data_out(10962),
        VN2CN1_bit => VN_data_out(10963),
        VN2CN2_bit => VN_data_out(10964),
        VN2CN3_bit => VN_data_out(10965),
        VN2CN4_bit => VN_data_out(10966),
        VN2CN5_bit => VN_data_out(10967),
        VN2CN0_sign => VN_sign_out(10962),
        VN2CN1_sign => VN_sign_out(10963),
        VN2CN2_sign => VN_sign_out(10964),
        VN2CN3_sign => VN_sign_out(10965),
        VN2CN4_sign => VN_sign_out(10966),
        VN2CN5_sign => VN_sign_out(10967),
        codeword => codeword(1827),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1828 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10973 downto 10968),
        Din0 => VN1828_in0,
        Din1 => VN1828_in1,
        Din2 => VN1828_in2,
        Din3 => VN1828_in3,
        Din4 => VN1828_in4,
        Din5 => VN1828_in5,
        VN2CN0_bit => VN_data_out(10968),
        VN2CN1_bit => VN_data_out(10969),
        VN2CN2_bit => VN_data_out(10970),
        VN2CN3_bit => VN_data_out(10971),
        VN2CN4_bit => VN_data_out(10972),
        VN2CN5_bit => VN_data_out(10973),
        VN2CN0_sign => VN_sign_out(10968),
        VN2CN1_sign => VN_sign_out(10969),
        VN2CN2_sign => VN_sign_out(10970),
        VN2CN3_sign => VN_sign_out(10971),
        VN2CN4_sign => VN_sign_out(10972),
        VN2CN5_sign => VN_sign_out(10973),
        codeword => codeword(1828),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1829 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10979 downto 10974),
        Din0 => VN1829_in0,
        Din1 => VN1829_in1,
        Din2 => VN1829_in2,
        Din3 => VN1829_in3,
        Din4 => VN1829_in4,
        Din5 => VN1829_in5,
        VN2CN0_bit => VN_data_out(10974),
        VN2CN1_bit => VN_data_out(10975),
        VN2CN2_bit => VN_data_out(10976),
        VN2CN3_bit => VN_data_out(10977),
        VN2CN4_bit => VN_data_out(10978),
        VN2CN5_bit => VN_data_out(10979),
        VN2CN0_sign => VN_sign_out(10974),
        VN2CN1_sign => VN_sign_out(10975),
        VN2CN2_sign => VN_sign_out(10976),
        VN2CN3_sign => VN_sign_out(10977),
        VN2CN4_sign => VN_sign_out(10978),
        VN2CN5_sign => VN_sign_out(10979),
        codeword => codeword(1829),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1830 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10985 downto 10980),
        Din0 => VN1830_in0,
        Din1 => VN1830_in1,
        Din2 => VN1830_in2,
        Din3 => VN1830_in3,
        Din4 => VN1830_in4,
        Din5 => VN1830_in5,
        VN2CN0_bit => VN_data_out(10980),
        VN2CN1_bit => VN_data_out(10981),
        VN2CN2_bit => VN_data_out(10982),
        VN2CN3_bit => VN_data_out(10983),
        VN2CN4_bit => VN_data_out(10984),
        VN2CN5_bit => VN_data_out(10985),
        VN2CN0_sign => VN_sign_out(10980),
        VN2CN1_sign => VN_sign_out(10981),
        VN2CN2_sign => VN_sign_out(10982),
        VN2CN3_sign => VN_sign_out(10983),
        VN2CN4_sign => VN_sign_out(10984),
        VN2CN5_sign => VN_sign_out(10985),
        codeword => codeword(1830),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1831 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10991 downto 10986),
        Din0 => VN1831_in0,
        Din1 => VN1831_in1,
        Din2 => VN1831_in2,
        Din3 => VN1831_in3,
        Din4 => VN1831_in4,
        Din5 => VN1831_in5,
        VN2CN0_bit => VN_data_out(10986),
        VN2CN1_bit => VN_data_out(10987),
        VN2CN2_bit => VN_data_out(10988),
        VN2CN3_bit => VN_data_out(10989),
        VN2CN4_bit => VN_data_out(10990),
        VN2CN5_bit => VN_data_out(10991),
        VN2CN0_sign => VN_sign_out(10986),
        VN2CN1_sign => VN_sign_out(10987),
        VN2CN2_sign => VN_sign_out(10988),
        VN2CN3_sign => VN_sign_out(10989),
        VN2CN4_sign => VN_sign_out(10990),
        VN2CN5_sign => VN_sign_out(10991),
        codeword => codeword(1831),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1832 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(10997 downto 10992),
        Din0 => VN1832_in0,
        Din1 => VN1832_in1,
        Din2 => VN1832_in2,
        Din3 => VN1832_in3,
        Din4 => VN1832_in4,
        Din5 => VN1832_in5,
        VN2CN0_bit => VN_data_out(10992),
        VN2CN1_bit => VN_data_out(10993),
        VN2CN2_bit => VN_data_out(10994),
        VN2CN3_bit => VN_data_out(10995),
        VN2CN4_bit => VN_data_out(10996),
        VN2CN5_bit => VN_data_out(10997),
        VN2CN0_sign => VN_sign_out(10992),
        VN2CN1_sign => VN_sign_out(10993),
        VN2CN2_sign => VN_sign_out(10994),
        VN2CN3_sign => VN_sign_out(10995),
        VN2CN4_sign => VN_sign_out(10996),
        VN2CN5_sign => VN_sign_out(10997),
        codeword => codeword(1832),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1833 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11003 downto 10998),
        Din0 => VN1833_in0,
        Din1 => VN1833_in1,
        Din2 => VN1833_in2,
        Din3 => VN1833_in3,
        Din4 => VN1833_in4,
        Din5 => VN1833_in5,
        VN2CN0_bit => VN_data_out(10998),
        VN2CN1_bit => VN_data_out(10999),
        VN2CN2_bit => VN_data_out(11000),
        VN2CN3_bit => VN_data_out(11001),
        VN2CN4_bit => VN_data_out(11002),
        VN2CN5_bit => VN_data_out(11003),
        VN2CN0_sign => VN_sign_out(10998),
        VN2CN1_sign => VN_sign_out(10999),
        VN2CN2_sign => VN_sign_out(11000),
        VN2CN3_sign => VN_sign_out(11001),
        VN2CN4_sign => VN_sign_out(11002),
        VN2CN5_sign => VN_sign_out(11003),
        codeword => codeword(1833),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1834 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11009 downto 11004),
        Din0 => VN1834_in0,
        Din1 => VN1834_in1,
        Din2 => VN1834_in2,
        Din3 => VN1834_in3,
        Din4 => VN1834_in4,
        Din5 => VN1834_in5,
        VN2CN0_bit => VN_data_out(11004),
        VN2CN1_bit => VN_data_out(11005),
        VN2CN2_bit => VN_data_out(11006),
        VN2CN3_bit => VN_data_out(11007),
        VN2CN4_bit => VN_data_out(11008),
        VN2CN5_bit => VN_data_out(11009),
        VN2CN0_sign => VN_sign_out(11004),
        VN2CN1_sign => VN_sign_out(11005),
        VN2CN2_sign => VN_sign_out(11006),
        VN2CN3_sign => VN_sign_out(11007),
        VN2CN4_sign => VN_sign_out(11008),
        VN2CN5_sign => VN_sign_out(11009),
        codeword => codeword(1834),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1835 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11015 downto 11010),
        Din0 => VN1835_in0,
        Din1 => VN1835_in1,
        Din2 => VN1835_in2,
        Din3 => VN1835_in3,
        Din4 => VN1835_in4,
        Din5 => VN1835_in5,
        VN2CN0_bit => VN_data_out(11010),
        VN2CN1_bit => VN_data_out(11011),
        VN2CN2_bit => VN_data_out(11012),
        VN2CN3_bit => VN_data_out(11013),
        VN2CN4_bit => VN_data_out(11014),
        VN2CN5_bit => VN_data_out(11015),
        VN2CN0_sign => VN_sign_out(11010),
        VN2CN1_sign => VN_sign_out(11011),
        VN2CN2_sign => VN_sign_out(11012),
        VN2CN3_sign => VN_sign_out(11013),
        VN2CN4_sign => VN_sign_out(11014),
        VN2CN5_sign => VN_sign_out(11015),
        codeword => codeword(1835),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1836 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11021 downto 11016),
        Din0 => VN1836_in0,
        Din1 => VN1836_in1,
        Din2 => VN1836_in2,
        Din3 => VN1836_in3,
        Din4 => VN1836_in4,
        Din5 => VN1836_in5,
        VN2CN0_bit => VN_data_out(11016),
        VN2CN1_bit => VN_data_out(11017),
        VN2CN2_bit => VN_data_out(11018),
        VN2CN3_bit => VN_data_out(11019),
        VN2CN4_bit => VN_data_out(11020),
        VN2CN5_bit => VN_data_out(11021),
        VN2CN0_sign => VN_sign_out(11016),
        VN2CN1_sign => VN_sign_out(11017),
        VN2CN2_sign => VN_sign_out(11018),
        VN2CN3_sign => VN_sign_out(11019),
        VN2CN4_sign => VN_sign_out(11020),
        VN2CN5_sign => VN_sign_out(11021),
        codeword => codeword(1836),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1837 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11027 downto 11022),
        Din0 => VN1837_in0,
        Din1 => VN1837_in1,
        Din2 => VN1837_in2,
        Din3 => VN1837_in3,
        Din4 => VN1837_in4,
        Din5 => VN1837_in5,
        VN2CN0_bit => VN_data_out(11022),
        VN2CN1_bit => VN_data_out(11023),
        VN2CN2_bit => VN_data_out(11024),
        VN2CN3_bit => VN_data_out(11025),
        VN2CN4_bit => VN_data_out(11026),
        VN2CN5_bit => VN_data_out(11027),
        VN2CN0_sign => VN_sign_out(11022),
        VN2CN1_sign => VN_sign_out(11023),
        VN2CN2_sign => VN_sign_out(11024),
        VN2CN3_sign => VN_sign_out(11025),
        VN2CN4_sign => VN_sign_out(11026),
        VN2CN5_sign => VN_sign_out(11027),
        codeword => codeword(1837),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1838 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11033 downto 11028),
        Din0 => VN1838_in0,
        Din1 => VN1838_in1,
        Din2 => VN1838_in2,
        Din3 => VN1838_in3,
        Din4 => VN1838_in4,
        Din5 => VN1838_in5,
        VN2CN0_bit => VN_data_out(11028),
        VN2CN1_bit => VN_data_out(11029),
        VN2CN2_bit => VN_data_out(11030),
        VN2CN3_bit => VN_data_out(11031),
        VN2CN4_bit => VN_data_out(11032),
        VN2CN5_bit => VN_data_out(11033),
        VN2CN0_sign => VN_sign_out(11028),
        VN2CN1_sign => VN_sign_out(11029),
        VN2CN2_sign => VN_sign_out(11030),
        VN2CN3_sign => VN_sign_out(11031),
        VN2CN4_sign => VN_sign_out(11032),
        VN2CN5_sign => VN_sign_out(11033),
        codeword => codeword(1838),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1839 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11039 downto 11034),
        Din0 => VN1839_in0,
        Din1 => VN1839_in1,
        Din2 => VN1839_in2,
        Din3 => VN1839_in3,
        Din4 => VN1839_in4,
        Din5 => VN1839_in5,
        VN2CN0_bit => VN_data_out(11034),
        VN2CN1_bit => VN_data_out(11035),
        VN2CN2_bit => VN_data_out(11036),
        VN2CN3_bit => VN_data_out(11037),
        VN2CN4_bit => VN_data_out(11038),
        VN2CN5_bit => VN_data_out(11039),
        VN2CN0_sign => VN_sign_out(11034),
        VN2CN1_sign => VN_sign_out(11035),
        VN2CN2_sign => VN_sign_out(11036),
        VN2CN3_sign => VN_sign_out(11037),
        VN2CN4_sign => VN_sign_out(11038),
        VN2CN5_sign => VN_sign_out(11039),
        codeword => codeword(1839),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1840 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11045 downto 11040),
        Din0 => VN1840_in0,
        Din1 => VN1840_in1,
        Din2 => VN1840_in2,
        Din3 => VN1840_in3,
        Din4 => VN1840_in4,
        Din5 => VN1840_in5,
        VN2CN0_bit => VN_data_out(11040),
        VN2CN1_bit => VN_data_out(11041),
        VN2CN2_bit => VN_data_out(11042),
        VN2CN3_bit => VN_data_out(11043),
        VN2CN4_bit => VN_data_out(11044),
        VN2CN5_bit => VN_data_out(11045),
        VN2CN0_sign => VN_sign_out(11040),
        VN2CN1_sign => VN_sign_out(11041),
        VN2CN2_sign => VN_sign_out(11042),
        VN2CN3_sign => VN_sign_out(11043),
        VN2CN4_sign => VN_sign_out(11044),
        VN2CN5_sign => VN_sign_out(11045),
        codeword => codeword(1840),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1841 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11051 downto 11046),
        Din0 => VN1841_in0,
        Din1 => VN1841_in1,
        Din2 => VN1841_in2,
        Din3 => VN1841_in3,
        Din4 => VN1841_in4,
        Din5 => VN1841_in5,
        VN2CN0_bit => VN_data_out(11046),
        VN2CN1_bit => VN_data_out(11047),
        VN2CN2_bit => VN_data_out(11048),
        VN2CN3_bit => VN_data_out(11049),
        VN2CN4_bit => VN_data_out(11050),
        VN2CN5_bit => VN_data_out(11051),
        VN2CN0_sign => VN_sign_out(11046),
        VN2CN1_sign => VN_sign_out(11047),
        VN2CN2_sign => VN_sign_out(11048),
        VN2CN3_sign => VN_sign_out(11049),
        VN2CN4_sign => VN_sign_out(11050),
        VN2CN5_sign => VN_sign_out(11051),
        codeword => codeword(1841),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1842 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11057 downto 11052),
        Din0 => VN1842_in0,
        Din1 => VN1842_in1,
        Din2 => VN1842_in2,
        Din3 => VN1842_in3,
        Din4 => VN1842_in4,
        Din5 => VN1842_in5,
        VN2CN0_bit => VN_data_out(11052),
        VN2CN1_bit => VN_data_out(11053),
        VN2CN2_bit => VN_data_out(11054),
        VN2CN3_bit => VN_data_out(11055),
        VN2CN4_bit => VN_data_out(11056),
        VN2CN5_bit => VN_data_out(11057),
        VN2CN0_sign => VN_sign_out(11052),
        VN2CN1_sign => VN_sign_out(11053),
        VN2CN2_sign => VN_sign_out(11054),
        VN2CN3_sign => VN_sign_out(11055),
        VN2CN4_sign => VN_sign_out(11056),
        VN2CN5_sign => VN_sign_out(11057),
        codeword => codeword(1842),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1843 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11063 downto 11058),
        Din0 => VN1843_in0,
        Din1 => VN1843_in1,
        Din2 => VN1843_in2,
        Din3 => VN1843_in3,
        Din4 => VN1843_in4,
        Din5 => VN1843_in5,
        VN2CN0_bit => VN_data_out(11058),
        VN2CN1_bit => VN_data_out(11059),
        VN2CN2_bit => VN_data_out(11060),
        VN2CN3_bit => VN_data_out(11061),
        VN2CN4_bit => VN_data_out(11062),
        VN2CN5_bit => VN_data_out(11063),
        VN2CN0_sign => VN_sign_out(11058),
        VN2CN1_sign => VN_sign_out(11059),
        VN2CN2_sign => VN_sign_out(11060),
        VN2CN3_sign => VN_sign_out(11061),
        VN2CN4_sign => VN_sign_out(11062),
        VN2CN5_sign => VN_sign_out(11063),
        codeword => codeword(1843),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1844 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11069 downto 11064),
        Din0 => VN1844_in0,
        Din1 => VN1844_in1,
        Din2 => VN1844_in2,
        Din3 => VN1844_in3,
        Din4 => VN1844_in4,
        Din5 => VN1844_in5,
        VN2CN0_bit => VN_data_out(11064),
        VN2CN1_bit => VN_data_out(11065),
        VN2CN2_bit => VN_data_out(11066),
        VN2CN3_bit => VN_data_out(11067),
        VN2CN4_bit => VN_data_out(11068),
        VN2CN5_bit => VN_data_out(11069),
        VN2CN0_sign => VN_sign_out(11064),
        VN2CN1_sign => VN_sign_out(11065),
        VN2CN2_sign => VN_sign_out(11066),
        VN2CN3_sign => VN_sign_out(11067),
        VN2CN4_sign => VN_sign_out(11068),
        VN2CN5_sign => VN_sign_out(11069),
        codeword => codeword(1844),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1845 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11075 downto 11070),
        Din0 => VN1845_in0,
        Din1 => VN1845_in1,
        Din2 => VN1845_in2,
        Din3 => VN1845_in3,
        Din4 => VN1845_in4,
        Din5 => VN1845_in5,
        VN2CN0_bit => VN_data_out(11070),
        VN2CN1_bit => VN_data_out(11071),
        VN2CN2_bit => VN_data_out(11072),
        VN2CN3_bit => VN_data_out(11073),
        VN2CN4_bit => VN_data_out(11074),
        VN2CN5_bit => VN_data_out(11075),
        VN2CN0_sign => VN_sign_out(11070),
        VN2CN1_sign => VN_sign_out(11071),
        VN2CN2_sign => VN_sign_out(11072),
        VN2CN3_sign => VN_sign_out(11073),
        VN2CN4_sign => VN_sign_out(11074),
        VN2CN5_sign => VN_sign_out(11075),
        codeword => codeword(1845),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1846 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11081 downto 11076),
        Din0 => VN1846_in0,
        Din1 => VN1846_in1,
        Din2 => VN1846_in2,
        Din3 => VN1846_in3,
        Din4 => VN1846_in4,
        Din5 => VN1846_in5,
        VN2CN0_bit => VN_data_out(11076),
        VN2CN1_bit => VN_data_out(11077),
        VN2CN2_bit => VN_data_out(11078),
        VN2CN3_bit => VN_data_out(11079),
        VN2CN4_bit => VN_data_out(11080),
        VN2CN5_bit => VN_data_out(11081),
        VN2CN0_sign => VN_sign_out(11076),
        VN2CN1_sign => VN_sign_out(11077),
        VN2CN2_sign => VN_sign_out(11078),
        VN2CN3_sign => VN_sign_out(11079),
        VN2CN4_sign => VN_sign_out(11080),
        VN2CN5_sign => VN_sign_out(11081),
        codeword => codeword(1846),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1847 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11087 downto 11082),
        Din0 => VN1847_in0,
        Din1 => VN1847_in1,
        Din2 => VN1847_in2,
        Din3 => VN1847_in3,
        Din4 => VN1847_in4,
        Din5 => VN1847_in5,
        VN2CN0_bit => VN_data_out(11082),
        VN2CN1_bit => VN_data_out(11083),
        VN2CN2_bit => VN_data_out(11084),
        VN2CN3_bit => VN_data_out(11085),
        VN2CN4_bit => VN_data_out(11086),
        VN2CN5_bit => VN_data_out(11087),
        VN2CN0_sign => VN_sign_out(11082),
        VN2CN1_sign => VN_sign_out(11083),
        VN2CN2_sign => VN_sign_out(11084),
        VN2CN3_sign => VN_sign_out(11085),
        VN2CN4_sign => VN_sign_out(11086),
        VN2CN5_sign => VN_sign_out(11087),
        codeword => codeword(1847),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1848 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11093 downto 11088),
        Din0 => VN1848_in0,
        Din1 => VN1848_in1,
        Din2 => VN1848_in2,
        Din3 => VN1848_in3,
        Din4 => VN1848_in4,
        Din5 => VN1848_in5,
        VN2CN0_bit => VN_data_out(11088),
        VN2CN1_bit => VN_data_out(11089),
        VN2CN2_bit => VN_data_out(11090),
        VN2CN3_bit => VN_data_out(11091),
        VN2CN4_bit => VN_data_out(11092),
        VN2CN5_bit => VN_data_out(11093),
        VN2CN0_sign => VN_sign_out(11088),
        VN2CN1_sign => VN_sign_out(11089),
        VN2CN2_sign => VN_sign_out(11090),
        VN2CN3_sign => VN_sign_out(11091),
        VN2CN4_sign => VN_sign_out(11092),
        VN2CN5_sign => VN_sign_out(11093),
        codeword => codeword(1848),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1849 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11099 downto 11094),
        Din0 => VN1849_in0,
        Din1 => VN1849_in1,
        Din2 => VN1849_in2,
        Din3 => VN1849_in3,
        Din4 => VN1849_in4,
        Din5 => VN1849_in5,
        VN2CN0_bit => VN_data_out(11094),
        VN2CN1_bit => VN_data_out(11095),
        VN2CN2_bit => VN_data_out(11096),
        VN2CN3_bit => VN_data_out(11097),
        VN2CN4_bit => VN_data_out(11098),
        VN2CN5_bit => VN_data_out(11099),
        VN2CN0_sign => VN_sign_out(11094),
        VN2CN1_sign => VN_sign_out(11095),
        VN2CN2_sign => VN_sign_out(11096),
        VN2CN3_sign => VN_sign_out(11097),
        VN2CN4_sign => VN_sign_out(11098),
        VN2CN5_sign => VN_sign_out(11099),
        codeword => codeword(1849),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1850 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11105 downto 11100),
        Din0 => VN1850_in0,
        Din1 => VN1850_in1,
        Din2 => VN1850_in2,
        Din3 => VN1850_in3,
        Din4 => VN1850_in4,
        Din5 => VN1850_in5,
        VN2CN0_bit => VN_data_out(11100),
        VN2CN1_bit => VN_data_out(11101),
        VN2CN2_bit => VN_data_out(11102),
        VN2CN3_bit => VN_data_out(11103),
        VN2CN4_bit => VN_data_out(11104),
        VN2CN5_bit => VN_data_out(11105),
        VN2CN0_sign => VN_sign_out(11100),
        VN2CN1_sign => VN_sign_out(11101),
        VN2CN2_sign => VN_sign_out(11102),
        VN2CN3_sign => VN_sign_out(11103),
        VN2CN4_sign => VN_sign_out(11104),
        VN2CN5_sign => VN_sign_out(11105),
        codeword => codeword(1850),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1851 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11111 downto 11106),
        Din0 => VN1851_in0,
        Din1 => VN1851_in1,
        Din2 => VN1851_in2,
        Din3 => VN1851_in3,
        Din4 => VN1851_in4,
        Din5 => VN1851_in5,
        VN2CN0_bit => VN_data_out(11106),
        VN2CN1_bit => VN_data_out(11107),
        VN2CN2_bit => VN_data_out(11108),
        VN2CN3_bit => VN_data_out(11109),
        VN2CN4_bit => VN_data_out(11110),
        VN2CN5_bit => VN_data_out(11111),
        VN2CN0_sign => VN_sign_out(11106),
        VN2CN1_sign => VN_sign_out(11107),
        VN2CN2_sign => VN_sign_out(11108),
        VN2CN3_sign => VN_sign_out(11109),
        VN2CN4_sign => VN_sign_out(11110),
        VN2CN5_sign => VN_sign_out(11111),
        codeword => codeword(1851),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1852 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11117 downto 11112),
        Din0 => VN1852_in0,
        Din1 => VN1852_in1,
        Din2 => VN1852_in2,
        Din3 => VN1852_in3,
        Din4 => VN1852_in4,
        Din5 => VN1852_in5,
        VN2CN0_bit => VN_data_out(11112),
        VN2CN1_bit => VN_data_out(11113),
        VN2CN2_bit => VN_data_out(11114),
        VN2CN3_bit => VN_data_out(11115),
        VN2CN4_bit => VN_data_out(11116),
        VN2CN5_bit => VN_data_out(11117),
        VN2CN0_sign => VN_sign_out(11112),
        VN2CN1_sign => VN_sign_out(11113),
        VN2CN2_sign => VN_sign_out(11114),
        VN2CN3_sign => VN_sign_out(11115),
        VN2CN4_sign => VN_sign_out(11116),
        VN2CN5_sign => VN_sign_out(11117),
        codeword => codeword(1852),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1853 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11123 downto 11118),
        Din0 => VN1853_in0,
        Din1 => VN1853_in1,
        Din2 => VN1853_in2,
        Din3 => VN1853_in3,
        Din4 => VN1853_in4,
        Din5 => VN1853_in5,
        VN2CN0_bit => VN_data_out(11118),
        VN2CN1_bit => VN_data_out(11119),
        VN2CN2_bit => VN_data_out(11120),
        VN2CN3_bit => VN_data_out(11121),
        VN2CN4_bit => VN_data_out(11122),
        VN2CN5_bit => VN_data_out(11123),
        VN2CN0_sign => VN_sign_out(11118),
        VN2CN1_sign => VN_sign_out(11119),
        VN2CN2_sign => VN_sign_out(11120),
        VN2CN3_sign => VN_sign_out(11121),
        VN2CN4_sign => VN_sign_out(11122),
        VN2CN5_sign => VN_sign_out(11123),
        codeword => codeword(1853),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1854 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11129 downto 11124),
        Din0 => VN1854_in0,
        Din1 => VN1854_in1,
        Din2 => VN1854_in2,
        Din3 => VN1854_in3,
        Din4 => VN1854_in4,
        Din5 => VN1854_in5,
        VN2CN0_bit => VN_data_out(11124),
        VN2CN1_bit => VN_data_out(11125),
        VN2CN2_bit => VN_data_out(11126),
        VN2CN3_bit => VN_data_out(11127),
        VN2CN4_bit => VN_data_out(11128),
        VN2CN5_bit => VN_data_out(11129),
        VN2CN0_sign => VN_sign_out(11124),
        VN2CN1_sign => VN_sign_out(11125),
        VN2CN2_sign => VN_sign_out(11126),
        VN2CN3_sign => VN_sign_out(11127),
        VN2CN4_sign => VN_sign_out(11128),
        VN2CN5_sign => VN_sign_out(11129),
        codeword => codeword(1854),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1855 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11135 downto 11130),
        Din0 => VN1855_in0,
        Din1 => VN1855_in1,
        Din2 => VN1855_in2,
        Din3 => VN1855_in3,
        Din4 => VN1855_in4,
        Din5 => VN1855_in5,
        VN2CN0_bit => VN_data_out(11130),
        VN2CN1_bit => VN_data_out(11131),
        VN2CN2_bit => VN_data_out(11132),
        VN2CN3_bit => VN_data_out(11133),
        VN2CN4_bit => VN_data_out(11134),
        VN2CN5_bit => VN_data_out(11135),
        VN2CN0_sign => VN_sign_out(11130),
        VN2CN1_sign => VN_sign_out(11131),
        VN2CN2_sign => VN_sign_out(11132),
        VN2CN3_sign => VN_sign_out(11133),
        VN2CN4_sign => VN_sign_out(11134),
        VN2CN5_sign => VN_sign_out(11135),
        codeword => codeword(1855),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1856 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11141 downto 11136),
        Din0 => VN1856_in0,
        Din1 => VN1856_in1,
        Din2 => VN1856_in2,
        Din3 => VN1856_in3,
        Din4 => VN1856_in4,
        Din5 => VN1856_in5,
        VN2CN0_bit => VN_data_out(11136),
        VN2CN1_bit => VN_data_out(11137),
        VN2CN2_bit => VN_data_out(11138),
        VN2CN3_bit => VN_data_out(11139),
        VN2CN4_bit => VN_data_out(11140),
        VN2CN5_bit => VN_data_out(11141),
        VN2CN0_sign => VN_sign_out(11136),
        VN2CN1_sign => VN_sign_out(11137),
        VN2CN2_sign => VN_sign_out(11138),
        VN2CN3_sign => VN_sign_out(11139),
        VN2CN4_sign => VN_sign_out(11140),
        VN2CN5_sign => VN_sign_out(11141),
        codeword => codeword(1856),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1857 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11147 downto 11142),
        Din0 => VN1857_in0,
        Din1 => VN1857_in1,
        Din2 => VN1857_in2,
        Din3 => VN1857_in3,
        Din4 => VN1857_in4,
        Din5 => VN1857_in5,
        VN2CN0_bit => VN_data_out(11142),
        VN2CN1_bit => VN_data_out(11143),
        VN2CN2_bit => VN_data_out(11144),
        VN2CN3_bit => VN_data_out(11145),
        VN2CN4_bit => VN_data_out(11146),
        VN2CN5_bit => VN_data_out(11147),
        VN2CN0_sign => VN_sign_out(11142),
        VN2CN1_sign => VN_sign_out(11143),
        VN2CN2_sign => VN_sign_out(11144),
        VN2CN3_sign => VN_sign_out(11145),
        VN2CN4_sign => VN_sign_out(11146),
        VN2CN5_sign => VN_sign_out(11147),
        codeword => codeword(1857),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1858 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11153 downto 11148),
        Din0 => VN1858_in0,
        Din1 => VN1858_in1,
        Din2 => VN1858_in2,
        Din3 => VN1858_in3,
        Din4 => VN1858_in4,
        Din5 => VN1858_in5,
        VN2CN0_bit => VN_data_out(11148),
        VN2CN1_bit => VN_data_out(11149),
        VN2CN2_bit => VN_data_out(11150),
        VN2CN3_bit => VN_data_out(11151),
        VN2CN4_bit => VN_data_out(11152),
        VN2CN5_bit => VN_data_out(11153),
        VN2CN0_sign => VN_sign_out(11148),
        VN2CN1_sign => VN_sign_out(11149),
        VN2CN2_sign => VN_sign_out(11150),
        VN2CN3_sign => VN_sign_out(11151),
        VN2CN4_sign => VN_sign_out(11152),
        VN2CN5_sign => VN_sign_out(11153),
        codeword => codeword(1858),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1859 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11159 downto 11154),
        Din0 => VN1859_in0,
        Din1 => VN1859_in1,
        Din2 => VN1859_in2,
        Din3 => VN1859_in3,
        Din4 => VN1859_in4,
        Din5 => VN1859_in5,
        VN2CN0_bit => VN_data_out(11154),
        VN2CN1_bit => VN_data_out(11155),
        VN2CN2_bit => VN_data_out(11156),
        VN2CN3_bit => VN_data_out(11157),
        VN2CN4_bit => VN_data_out(11158),
        VN2CN5_bit => VN_data_out(11159),
        VN2CN0_sign => VN_sign_out(11154),
        VN2CN1_sign => VN_sign_out(11155),
        VN2CN2_sign => VN_sign_out(11156),
        VN2CN3_sign => VN_sign_out(11157),
        VN2CN4_sign => VN_sign_out(11158),
        VN2CN5_sign => VN_sign_out(11159),
        codeword => codeword(1859),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1860 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11165 downto 11160),
        Din0 => VN1860_in0,
        Din1 => VN1860_in1,
        Din2 => VN1860_in2,
        Din3 => VN1860_in3,
        Din4 => VN1860_in4,
        Din5 => VN1860_in5,
        VN2CN0_bit => VN_data_out(11160),
        VN2CN1_bit => VN_data_out(11161),
        VN2CN2_bit => VN_data_out(11162),
        VN2CN3_bit => VN_data_out(11163),
        VN2CN4_bit => VN_data_out(11164),
        VN2CN5_bit => VN_data_out(11165),
        VN2CN0_sign => VN_sign_out(11160),
        VN2CN1_sign => VN_sign_out(11161),
        VN2CN2_sign => VN_sign_out(11162),
        VN2CN3_sign => VN_sign_out(11163),
        VN2CN4_sign => VN_sign_out(11164),
        VN2CN5_sign => VN_sign_out(11165),
        codeword => codeword(1860),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1861 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11171 downto 11166),
        Din0 => VN1861_in0,
        Din1 => VN1861_in1,
        Din2 => VN1861_in2,
        Din3 => VN1861_in3,
        Din4 => VN1861_in4,
        Din5 => VN1861_in5,
        VN2CN0_bit => VN_data_out(11166),
        VN2CN1_bit => VN_data_out(11167),
        VN2CN2_bit => VN_data_out(11168),
        VN2CN3_bit => VN_data_out(11169),
        VN2CN4_bit => VN_data_out(11170),
        VN2CN5_bit => VN_data_out(11171),
        VN2CN0_sign => VN_sign_out(11166),
        VN2CN1_sign => VN_sign_out(11167),
        VN2CN2_sign => VN_sign_out(11168),
        VN2CN3_sign => VN_sign_out(11169),
        VN2CN4_sign => VN_sign_out(11170),
        VN2CN5_sign => VN_sign_out(11171),
        codeword => codeword(1861),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1862 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11177 downto 11172),
        Din0 => VN1862_in0,
        Din1 => VN1862_in1,
        Din2 => VN1862_in2,
        Din3 => VN1862_in3,
        Din4 => VN1862_in4,
        Din5 => VN1862_in5,
        VN2CN0_bit => VN_data_out(11172),
        VN2CN1_bit => VN_data_out(11173),
        VN2CN2_bit => VN_data_out(11174),
        VN2CN3_bit => VN_data_out(11175),
        VN2CN4_bit => VN_data_out(11176),
        VN2CN5_bit => VN_data_out(11177),
        VN2CN0_sign => VN_sign_out(11172),
        VN2CN1_sign => VN_sign_out(11173),
        VN2CN2_sign => VN_sign_out(11174),
        VN2CN3_sign => VN_sign_out(11175),
        VN2CN4_sign => VN_sign_out(11176),
        VN2CN5_sign => VN_sign_out(11177),
        codeword => codeword(1862),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1863 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11183 downto 11178),
        Din0 => VN1863_in0,
        Din1 => VN1863_in1,
        Din2 => VN1863_in2,
        Din3 => VN1863_in3,
        Din4 => VN1863_in4,
        Din5 => VN1863_in5,
        VN2CN0_bit => VN_data_out(11178),
        VN2CN1_bit => VN_data_out(11179),
        VN2CN2_bit => VN_data_out(11180),
        VN2CN3_bit => VN_data_out(11181),
        VN2CN4_bit => VN_data_out(11182),
        VN2CN5_bit => VN_data_out(11183),
        VN2CN0_sign => VN_sign_out(11178),
        VN2CN1_sign => VN_sign_out(11179),
        VN2CN2_sign => VN_sign_out(11180),
        VN2CN3_sign => VN_sign_out(11181),
        VN2CN4_sign => VN_sign_out(11182),
        VN2CN5_sign => VN_sign_out(11183),
        codeword => codeword(1863),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1864 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11189 downto 11184),
        Din0 => VN1864_in0,
        Din1 => VN1864_in1,
        Din2 => VN1864_in2,
        Din3 => VN1864_in3,
        Din4 => VN1864_in4,
        Din5 => VN1864_in5,
        VN2CN0_bit => VN_data_out(11184),
        VN2CN1_bit => VN_data_out(11185),
        VN2CN2_bit => VN_data_out(11186),
        VN2CN3_bit => VN_data_out(11187),
        VN2CN4_bit => VN_data_out(11188),
        VN2CN5_bit => VN_data_out(11189),
        VN2CN0_sign => VN_sign_out(11184),
        VN2CN1_sign => VN_sign_out(11185),
        VN2CN2_sign => VN_sign_out(11186),
        VN2CN3_sign => VN_sign_out(11187),
        VN2CN4_sign => VN_sign_out(11188),
        VN2CN5_sign => VN_sign_out(11189),
        codeword => codeword(1864),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1865 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11195 downto 11190),
        Din0 => VN1865_in0,
        Din1 => VN1865_in1,
        Din2 => VN1865_in2,
        Din3 => VN1865_in3,
        Din4 => VN1865_in4,
        Din5 => VN1865_in5,
        VN2CN0_bit => VN_data_out(11190),
        VN2CN1_bit => VN_data_out(11191),
        VN2CN2_bit => VN_data_out(11192),
        VN2CN3_bit => VN_data_out(11193),
        VN2CN4_bit => VN_data_out(11194),
        VN2CN5_bit => VN_data_out(11195),
        VN2CN0_sign => VN_sign_out(11190),
        VN2CN1_sign => VN_sign_out(11191),
        VN2CN2_sign => VN_sign_out(11192),
        VN2CN3_sign => VN_sign_out(11193),
        VN2CN4_sign => VN_sign_out(11194),
        VN2CN5_sign => VN_sign_out(11195),
        codeword => codeword(1865),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1866 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11201 downto 11196),
        Din0 => VN1866_in0,
        Din1 => VN1866_in1,
        Din2 => VN1866_in2,
        Din3 => VN1866_in3,
        Din4 => VN1866_in4,
        Din5 => VN1866_in5,
        VN2CN0_bit => VN_data_out(11196),
        VN2CN1_bit => VN_data_out(11197),
        VN2CN2_bit => VN_data_out(11198),
        VN2CN3_bit => VN_data_out(11199),
        VN2CN4_bit => VN_data_out(11200),
        VN2CN5_bit => VN_data_out(11201),
        VN2CN0_sign => VN_sign_out(11196),
        VN2CN1_sign => VN_sign_out(11197),
        VN2CN2_sign => VN_sign_out(11198),
        VN2CN3_sign => VN_sign_out(11199),
        VN2CN4_sign => VN_sign_out(11200),
        VN2CN5_sign => VN_sign_out(11201),
        codeword => codeword(1866),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1867 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11207 downto 11202),
        Din0 => VN1867_in0,
        Din1 => VN1867_in1,
        Din2 => VN1867_in2,
        Din3 => VN1867_in3,
        Din4 => VN1867_in4,
        Din5 => VN1867_in5,
        VN2CN0_bit => VN_data_out(11202),
        VN2CN1_bit => VN_data_out(11203),
        VN2CN2_bit => VN_data_out(11204),
        VN2CN3_bit => VN_data_out(11205),
        VN2CN4_bit => VN_data_out(11206),
        VN2CN5_bit => VN_data_out(11207),
        VN2CN0_sign => VN_sign_out(11202),
        VN2CN1_sign => VN_sign_out(11203),
        VN2CN2_sign => VN_sign_out(11204),
        VN2CN3_sign => VN_sign_out(11205),
        VN2CN4_sign => VN_sign_out(11206),
        VN2CN5_sign => VN_sign_out(11207),
        codeword => codeword(1867),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1868 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11213 downto 11208),
        Din0 => VN1868_in0,
        Din1 => VN1868_in1,
        Din2 => VN1868_in2,
        Din3 => VN1868_in3,
        Din4 => VN1868_in4,
        Din5 => VN1868_in5,
        VN2CN0_bit => VN_data_out(11208),
        VN2CN1_bit => VN_data_out(11209),
        VN2CN2_bit => VN_data_out(11210),
        VN2CN3_bit => VN_data_out(11211),
        VN2CN4_bit => VN_data_out(11212),
        VN2CN5_bit => VN_data_out(11213),
        VN2CN0_sign => VN_sign_out(11208),
        VN2CN1_sign => VN_sign_out(11209),
        VN2CN2_sign => VN_sign_out(11210),
        VN2CN3_sign => VN_sign_out(11211),
        VN2CN4_sign => VN_sign_out(11212),
        VN2CN5_sign => VN_sign_out(11213),
        codeword => codeword(1868),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1869 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11219 downto 11214),
        Din0 => VN1869_in0,
        Din1 => VN1869_in1,
        Din2 => VN1869_in2,
        Din3 => VN1869_in3,
        Din4 => VN1869_in4,
        Din5 => VN1869_in5,
        VN2CN0_bit => VN_data_out(11214),
        VN2CN1_bit => VN_data_out(11215),
        VN2CN2_bit => VN_data_out(11216),
        VN2CN3_bit => VN_data_out(11217),
        VN2CN4_bit => VN_data_out(11218),
        VN2CN5_bit => VN_data_out(11219),
        VN2CN0_sign => VN_sign_out(11214),
        VN2CN1_sign => VN_sign_out(11215),
        VN2CN2_sign => VN_sign_out(11216),
        VN2CN3_sign => VN_sign_out(11217),
        VN2CN4_sign => VN_sign_out(11218),
        VN2CN5_sign => VN_sign_out(11219),
        codeword => codeword(1869),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1870 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11225 downto 11220),
        Din0 => VN1870_in0,
        Din1 => VN1870_in1,
        Din2 => VN1870_in2,
        Din3 => VN1870_in3,
        Din4 => VN1870_in4,
        Din5 => VN1870_in5,
        VN2CN0_bit => VN_data_out(11220),
        VN2CN1_bit => VN_data_out(11221),
        VN2CN2_bit => VN_data_out(11222),
        VN2CN3_bit => VN_data_out(11223),
        VN2CN4_bit => VN_data_out(11224),
        VN2CN5_bit => VN_data_out(11225),
        VN2CN0_sign => VN_sign_out(11220),
        VN2CN1_sign => VN_sign_out(11221),
        VN2CN2_sign => VN_sign_out(11222),
        VN2CN3_sign => VN_sign_out(11223),
        VN2CN4_sign => VN_sign_out(11224),
        VN2CN5_sign => VN_sign_out(11225),
        codeword => codeword(1870),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1871 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11231 downto 11226),
        Din0 => VN1871_in0,
        Din1 => VN1871_in1,
        Din2 => VN1871_in2,
        Din3 => VN1871_in3,
        Din4 => VN1871_in4,
        Din5 => VN1871_in5,
        VN2CN0_bit => VN_data_out(11226),
        VN2CN1_bit => VN_data_out(11227),
        VN2CN2_bit => VN_data_out(11228),
        VN2CN3_bit => VN_data_out(11229),
        VN2CN4_bit => VN_data_out(11230),
        VN2CN5_bit => VN_data_out(11231),
        VN2CN0_sign => VN_sign_out(11226),
        VN2CN1_sign => VN_sign_out(11227),
        VN2CN2_sign => VN_sign_out(11228),
        VN2CN3_sign => VN_sign_out(11229),
        VN2CN4_sign => VN_sign_out(11230),
        VN2CN5_sign => VN_sign_out(11231),
        codeword => codeword(1871),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1872 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11237 downto 11232),
        Din0 => VN1872_in0,
        Din1 => VN1872_in1,
        Din2 => VN1872_in2,
        Din3 => VN1872_in3,
        Din4 => VN1872_in4,
        Din5 => VN1872_in5,
        VN2CN0_bit => VN_data_out(11232),
        VN2CN1_bit => VN_data_out(11233),
        VN2CN2_bit => VN_data_out(11234),
        VN2CN3_bit => VN_data_out(11235),
        VN2CN4_bit => VN_data_out(11236),
        VN2CN5_bit => VN_data_out(11237),
        VN2CN0_sign => VN_sign_out(11232),
        VN2CN1_sign => VN_sign_out(11233),
        VN2CN2_sign => VN_sign_out(11234),
        VN2CN3_sign => VN_sign_out(11235),
        VN2CN4_sign => VN_sign_out(11236),
        VN2CN5_sign => VN_sign_out(11237),
        codeword => codeword(1872),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1873 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11243 downto 11238),
        Din0 => VN1873_in0,
        Din1 => VN1873_in1,
        Din2 => VN1873_in2,
        Din3 => VN1873_in3,
        Din4 => VN1873_in4,
        Din5 => VN1873_in5,
        VN2CN0_bit => VN_data_out(11238),
        VN2CN1_bit => VN_data_out(11239),
        VN2CN2_bit => VN_data_out(11240),
        VN2CN3_bit => VN_data_out(11241),
        VN2CN4_bit => VN_data_out(11242),
        VN2CN5_bit => VN_data_out(11243),
        VN2CN0_sign => VN_sign_out(11238),
        VN2CN1_sign => VN_sign_out(11239),
        VN2CN2_sign => VN_sign_out(11240),
        VN2CN3_sign => VN_sign_out(11241),
        VN2CN4_sign => VN_sign_out(11242),
        VN2CN5_sign => VN_sign_out(11243),
        codeword => codeword(1873),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1874 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11249 downto 11244),
        Din0 => VN1874_in0,
        Din1 => VN1874_in1,
        Din2 => VN1874_in2,
        Din3 => VN1874_in3,
        Din4 => VN1874_in4,
        Din5 => VN1874_in5,
        VN2CN0_bit => VN_data_out(11244),
        VN2CN1_bit => VN_data_out(11245),
        VN2CN2_bit => VN_data_out(11246),
        VN2CN3_bit => VN_data_out(11247),
        VN2CN4_bit => VN_data_out(11248),
        VN2CN5_bit => VN_data_out(11249),
        VN2CN0_sign => VN_sign_out(11244),
        VN2CN1_sign => VN_sign_out(11245),
        VN2CN2_sign => VN_sign_out(11246),
        VN2CN3_sign => VN_sign_out(11247),
        VN2CN4_sign => VN_sign_out(11248),
        VN2CN5_sign => VN_sign_out(11249),
        codeword => codeword(1874),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1875 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11255 downto 11250),
        Din0 => VN1875_in0,
        Din1 => VN1875_in1,
        Din2 => VN1875_in2,
        Din3 => VN1875_in3,
        Din4 => VN1875_in4,
        Din5 => VN1875_in5,
        VN2CN0_bit => VN_data_out(11250),
        VN2CN1_bit => VN_data_out(11251),
        VN2CN2_bit => VN_data_out(11252),
        VN2CN3_bit => VN_data_out(11253),
        VN2CN4_bit => VN_data_out(11254),
        VN2CN5_bit => VN_data_out(11255),
        VN2CN0_sign => VN_sign_out(11250),
        VN2CN1_sign => VN_sign_out(11251),
        VN2CN2_sign => VN_sign_out(11252),
        VN2CN3_sign => VN_sign_out(11253),
        VN2CN4_sign => VN_sign_out(11254),
        VN2CN5_sign => VN_sign_out(11255),
        codeword => codeword(1875),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1876 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11261 downto 11256),
        Din0 => VN1876_in0,
        Din1 => VN1876_in1,
        Din2 => VN1876_in2,
        Din3 => VN1876_in3,
        Din4 => VN1876_in4,
        Din5 => VN1876_in5,
        VN2CN0_bit => VN_data_out(11256),
        VN2CN1_bit => VN_data_out(11257),
        VN2CN2_bit => VN_data_out(11258),
        VN2CN3_bit => VN_data_out(11259),
        VN2CN4_bit => VN_data_out(11260),
        VN2CN5_bit => VN_data_out(11261),
        VN2CN0_sign => VN_sign_out(11256),
        VN2CN1_sign => VN_sign_out(11257),
        VN2CN2_sign => VN_sign_out(11258),
        VN2CN3_sign => VN_sign_out(11259),
        VN2CN4_sign => VN_sign_out(11260),
        VN2CN5_sign => VN_sign_out(11261),
        codeword => codeword(1876),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1877 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11267 downto 11262),
        Din0 => VN1877_in0,
        Din1 => VN1877_in1,
        Din2 => VN1877_in2,
        Din3 => VN1877_in3,
        Din4 => VN1877_in4,
        Din5 => VN1877_in5,
        VN2CN0_bit => VN_data_out(11262),
        VN2CN1_bit => VN_data_out(11263),
        VN2CN2_bit => VN_data_out(11264),
        VN2CN3_bit => VN_data_out(11265),
        VN2CN4_bit => VN_data_out(11266),
        VN2CN5_bit => VN_data_out(11267),
        VN2CN0_sign => VN_sign_out(11262),
        VN2CN1_sign => VN_sign_out(11263),
        VN2CN2_sign => VN_sign_out(11264),
        VN2CN3_sign => VN_sign_out(11265),
        VN2CN4_sign => VN_sign_out(11266),
        VN2CN5_sign => VN_sign_out(11267),
        codeword => codeword(1877),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1878 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11273 downto 11268),
        Din0 => VN1878_in0,
        Din1 => VN1878_in1,
        Din2 => VN1878_in2,
        Din3 => VN1878_in3,
        Din4 => VN1878_in4,
        Din5 => VN1878_in5,
        VN2CN0_bit => VN_data_out(11268),
        VN2CN1_bit => VN_data_out(11269),
        VN2CN2_bit => VN_data_out(11270),
        VN2CN3_bit => VN_data_out(11271),
        VN2CN4_bit => VN_data_out(11272),
        VN2CN5_bit => VN_data_out(11273),
        VN2CN0_sign => VN_sign_out(11268),
        VN2CN1_sign => VN_sign_out(11269),
        VN2CN2_sign => VN_sign_out(11270),
        VN2CN3_sign => VN_sign_out(11271),
        VN2CN4_sign => VN_sign_out(11272),
        VN2CN5_sign => VN_sign_out(11273),
        codeword => codeword(1878),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1879 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11279 downto 11274),
        Din0 => VN1879_in0,
        Din1 => VN1879_in1,
        Din2 => VN1879_in2,
        Din3 => VN1879_in3,
        Din4 => VN1879_in4,
        Din5 => VN1879_in5,
        VN2CN0_bit => VN_data_out(11274),
        VN2CN1_bit => VN_data_out(11275),
        VN2CN2_bit => VN_data_out(11276),
        VN2CN3_bit => VN_data_out(11277),
        VN2CN4_bit => VN_data_out(11278),
        VN2CN5_bit => VN_data_out(11279),
        VN2CN0_sign => VN_sign_out(11274),
        VN2CN1_sign => VN_sign_out(11275),
        VN2CN2_sign => VN_sign_out(11276),
        VN2CN3_sign => VN_sign_out(11277),
        VN2CN4_sign => VN_sign_out(11278),
        VN2CN5_sign => VN_sign_out(11279),
        codeword => codeword(1879),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1880 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11285 downto 11280),
        Din0 => VN1880_in0,
        Din1 => VN1880_in1,
        Din2 => VN1880_in2,
        Din3 => VN1880_in3,
        Din4 => VN1880_in4,
        Din5 => VN1880_in5,
        VN2CN0_bit => VN_data_out(11280),
        VN2CN1_bit => VN_data_out(11281),
        VN2CN2_bit => VN_data_out(11282),
        VN2CN3_bit => VN_data_out(11283),
        VN2CN4_bit => VN_data_out(11284),
        VN2CN5_bit => VN_data_out(11285),
        VN2CN0_sign => VN_sign_out(11280),
        VN2CN1_sign => VN_sign_out(11281),
        VN2CN2_sign => VN_sign_out(11282),
        VN2CN3_sign => VN_sign_out(11283),
        VN2CN4_sign => VN_sign_out(11284),
        VN2CN5_sign => VN_sign_out(11285),
        codeword => codeword(1880),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1881 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11291 downto 11286),
        Din0 => VN1881_in0,
        Din1 => VN1881_in1,
        Din2 => VN1881_in2,
        Din3 => VN1881_in3,
        Din4 => VN1881_in4,
        Din5 => VN1881_in5,
        VN2CN0_bit => VN_data_out(11286),
        VN2CN1_bit => VN_data_out(11287),
        VN2CN2_bit => VN_data_out(11288),
        VN2CN3_bit => VN_data_out(11289),
        VN2CN4_bit => VN_data_out(11290),
        VN2CN5_bit => VN_data_out(11291),
        VN2CN0_sign => VN_sign_out(11286),
        VN2CN1_sign => VN_sign_out(11287),
        VN2CN2_sign => VN_sign_out(11288),
        VN2CN3_sign => VN_sign_out(11289),
        VN2CN4_sign => VN_sign_out(11290),
        VN2CN5_sign => VN_sign_out(11291),
        codeword => codeword(1881),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1882 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11297 downto 11292),
        Din0 => VN1882_in0,
        Din1 => VN1882_in1,
        Din2 => VN1882_in2,
        Din3 => VN1882_in3,
        Din4 => VN1882_in4,
        Din5 => VN1882_in5,
        VN2CN0_bit => VN_data_out(11292),
        VN2CN1_bit => VN_data_out(11293),
        VN2CN2_bit => VN_data_out(11294),
        VN2CN3_bit => VN_data_out(11295),
        VN2CN4_bit => VN_data_out(11296),
        VN2CN5_bit => VN_data_out(11297),
        VN2CN0_sign => VN_sign_out(11292),
        VN2CN1_sign => VN_sign_out(11293),
        VN2CN2_sign => VN_sign_out(11294),
        VN2CN3_sign => VN_sign_out(11295),
        VN2CN4_sign => VN_sign_out(11296),
        VN2CN5_sign => VN_sign_out(11297),
        codeword => codeword(1882),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1883 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11303 downto 11298),
        Din0 => VN1883_in0,
        Din1 => VN1883_in1,
        Din2 => VN1883_in2,
        Din3 => VN1883_in3,
        Din4 => VN1883_in4,
        Din5 => VN1883_in5,
        VN2CN0_bit => VN_data_out(11298),
        VN2CN1_bit => VN_data_out(11299),
        VN2CN2_bit => VN_data_out(11300),
        VN2CN3_bit => VN_data_out(11301),
        VN2CN4_bit => VN_data_out(11302),
        VN2CN5_bit => VN_data_out(11303),
        VN2CN0_sign => VN_sign_out(11298),
        VN2CN1_sign => VN_sign_out(11299),
        VN2CN2_sign => VN_sign_out(11300),
        VN2CN3_sign => VN_sign_out(11301),
        VN2CN4_sign => VN_sign_out(11302),
        VN2CN5_sign => VN_sign_out(11303),
        codeword => codeword(1883),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1884 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11309 downto 11304),
        Din0 => VN1884_in0,
        Din1 => VN1884_in1,
        Din2 => VN1884_in2,
        Din3 => VN1884_in3,
        Din4 => VN1884_in4,
        Din5 => VN1884_in5,
        VN2CN0_bit => VN_data_out(11304),
        VN2CN1_bit => VN_data_out(11305),
        VN2CN2_bit => VN_data_out(11306),
        VN2CN3_bit => VN_data_out(11307),
        VN2CN4_bit => VN_data_out(11308),
        VN2CN5_bit => VN_data_out(11309),
        VN2CN0_sign => VN_sign_out(11304),
        VN2CN1_sign => VN_sign_out(11305),
        VN2CN2_sign => VN_sign_out(11306),
        VN2CN3_sign => VN_sign_out(11307),
        VN2CN4_sign => VN_sign_out(11308),
        VN2CN5_sign => VN_sign_out(11309),
        codeword => codeword(1884),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1885 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11315 downto 11310),
        Din0 => VN1885_in0,
        Din1 => VN1885_in1,
        Din2 => VN1885_in2,
        Din3 => VN1885_in3,
        Din4 => VN1885_in4,
        Din5 => VN1885_in5,
        VN2CN0_bit => VN_data_out(11310),
        VN2CN1_bit => VN_data_out(11311),
        VN2CN2_bit => VN_data_out(11312),
        VN2CN3_bit => VN_data_out(11313),
        VN2CN4_bit => VN_data_out(11314),
        VN2CN5_bit => VN_data_out(11315),
        VN2CN0_sign => VN_sign_out(11310),
        VN2CN1_sign => VN_sign_out(11311),
        VN2CN2_sign => VN_sign_out(11312),
        VN2CN3_sign => VN_sign_out(11313),
        VN2CN4_sign => VN_sign_out(11314),
        VN2CN5_sign => VN_sign_out(11315),
        codeword => codeword(1885),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1886 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11321 downto 11316),
        Din0 => VN1886_in0,
        Din1 => VN1886_in1,
        Din2 => VN1886_in2,
        Din3 => VN1886_in3,
        Din4 => VN1886_in4,
        Din5 => VN1886_in5,
        VN2CN0_bit => VN_data_out(11316),
        VN2CN1_bit => VN_data_out(11317),
        VN2CN2_bit => VN_data_out(11318),
        VN2CN3_bit => VN_data_out(11319),
        VN2CN4_bit => VN_data_out(11320),
        VN2CN5_bit => VN_data_out(11321),
        VN2CN0_sign => VN_sign_out(11316),
        VN2CN1_sign => VN_sign_out(11317),
        VN2CN2_sign => VN_sign_out(11318),
        VN2CN3_sign => VN_sign_out(11319),
        VN2CN4_sign => VN_sign_out(11320),
        VN2CN5_sign => VN_sign_out(11321),
        codeword => codeword(1886),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1887 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11327 downto 11322),
        Din0 => VN1887_in0,
        Din1 => VN1887_in1,
        Din2 => VN1887_in2,
        Din3 => VN1887_in3,
        Din4 => VN1887_in4,
        Din5 => VN1887_in5,
        VN2CN0_bit => VN_data_out(11322),
        VN2CN1_bit => VN_data_out(11323),
        VN2CN2_bit => VN_data_out(11324),
        VN2CN3_bit => VN_data_out(11325),
        VN2CN4_bit => VN_data_out(11326),
        VN2CN5_bit => VN_data_out(11327),
        VN2CN0_sign => VN_sign_out(11322),
        VN2CN1_sign => VN_sign_out(11323),
        VN2CN2_sign => VN_sign_out(11324),
        VN2CN3_sign => VN_sign_out(11325),
        VN2CN4_sign => VN_sign_out(11326),
        VN2CN5_sign => VN_sign_out(11327),
        codeword => codeword(1887),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1888 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11333 downto 11328),
        Din0 => VN1888_in0,
        Din1 => VN1888_in1,
        Din2 => VN1888_in2,
        Din3 => VN1888_in3,
        Din4 => VN1888_in4,
        Din5 => VN1888_in5,
        VN2CN0_bit => VN_data_out(11328),
        VN2CN1_bit => VN_data_out(11329),
        VN2CN2_bit => VN_data_out(11330),
        VN2CN3_bit => VN_data_out(11331),
        VN2CN4_bit => VN_data_out(11332),
        VN2CN5_bit => VN_data_out(11333),
        VN2CN0_sign => VN_sign_out(11328),
        VN2CN1_sign => VN_sign_out(11329),
        VN2CN2_sign => VN_sign_out(11330),
        VN2CN3_sign => VN_sign_out(11331),
        VN2CN4_sign => VN_sign_out(11332),
        VN2CN5_sign => VN_sign_out(11333),
        codeword => codeword(1888),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1889 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11339 downto 11334),
        Din0 => VN1889_in0,
        Din1 => VN1889_in1,
        Din2 => VN1889_in2,
        Din3 => VN1889_in3,
        Din4 => VN1889_in4,
        Din5 => VN1889_in5,
        VN2CN0_bit => VN_data_out(11334),
        VN2CN1_bit => VN_data_out(11335),
        VN2CN2_bit => VN_data_out(11336),
        VN2CN3_bit => VN_data_out(11337),
        VN2CN4_bit => VN_data_out(11338),
        VN2CN5_bit => VN_data_out(11339),
        VN2CN0_sign => VN_sign_out(11334),
        VN2CN1_sign => VN_sign_out(11335),
        VN2CN2_sign => VN_sign_out(11336),
        VN2CN3_sign => VN_sign_out(11337),
        VN2CN4_sign => VN_sign_out(11338),
        VN2CN5_sign => VN_sign_out(11339),
        codeword => codeword(1889),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1890 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11345 downto 11340),
        Din0 => VN1890_in0,
        Din1 => VN1890_in1,
        Din2 => VN1890_in2,
        Din3 => VN1890_in3,
        Din4 => VN1890_in4,
        Din5 => VN1890_in5,
        VN2CN0_bit => VN_data_out(11340),
        VN2CN1_bit => VN_data_out(11341),
        VN2CN2_bit => VN_data_out(11342),
        VN2CN3_bit => VN_data_out(11343),
        VN2CN4_bit => VN_data_out(11344),
        VN2CN5_bit => VN_data_out(11345),
        VN2CN0_sign => VN_sign_out(11340),
        VN2CN1_sign => VN_sign_out(11341),
        VN2CN2_sign => VN_sign_out(11342),
        VN2CN3_sign => VN_sign_out(11343),
        VN2CN4_sign => VN_sign_out(11344),
        VN2CN5_sign => VN_sign_out(11345),
        codeword => codeword(1890),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1891 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11351 downto 11346),
        Din0 => VN1891_in0,
        Din1 => VN1891_in1,
        Din2 => VN1891_in2,
        Din3 => VN1891_in3,
        Din4 => VN1891_in4,
        Din5 => VN1891_in5,
        VN2CN0_bit => VN_data_out(11346),
        VN2CN1_bit => VN_data_out(11347),
        VN2CN2_bit => VN_data_out(11348),
        VN2CN3_bit => VN_data_out(11349),
        VN2CN4_bit => VN_data_out(11350),
        VN2CN5_bit => VN_data_out(11351),
        VN2CN0_sign => VN_sign_out(11346),
        VN2CN1_sign => VN_sign_out(11347),
        VN2CN2_sign => VN_sign_out(11348),
        VN2CN3_sign => VN_sign_out(11349),
        VN2CN4_sign => VN_sign_out(11350),
        VN2CN5_sign => VN_sign_out(11351),
        codeword => codeword(1891),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1892 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11357 downto 11352),
        Din0 => VN1892_in0,
        Din1 => VN1892_in1,
        Din2 => VN1892_in2,
        Din3 => VN1892_in3,
        Din4 => VN1892_in4,
        Din5 => VN1892_in5,
        VN2CN0_bit => VN_data_out(11352),
        VN2CN1_bit => VN_data_out(11353),
        VN2CN2_bit => VN_data_out(11354),
        VN2CN3_bit => VN_data_out(11355),
        VN2CN4_bit => VN_data_out(11356),
        VN2CN5_bit => VN_data_out(11357),
        VN2CN0_sign => VN_sign_out(11352),
        VN2CN1_sign => VN_sign_out(11353),
        VN2CN2_sign => VN_sign_out(11354),
        VN2CN3_sign => VN_sign_out(11355),
        VN2CN4_sign => VN_sign_out(11356),
        VN2CN5_sign => VN_sign_out(11357),
        codeword => codeword(1892),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1893 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11363 downto 11358),
        Din0 => VN1893_in0,
        Din1 => VN1893_in1,
        Din2 => VN1893_in2,
        Din3 => VN1893_in3,
        Din4 => VN1893_in4,
        Din5 => VN1893_in5,
        VN2CN0_bit => VN_data_out(11358),
        VN2CN1_bit => VN_data_out(11359),
        VN2CN2_bit => VN_data_out(11360),
        VN2CN3_bit => VN_data_out(11361),
        VN2CN4_bit => VN_data_out(11362),
        VN2CN5_bit => VN_data_out(11363),
        VN2CN0_sign => VN_sign_out(11358),
        VN2CN1_sign => VN_sign_out(11359),
        VN2CN2_sign => VN_sign_out(11360),
        VN2CN3_sign => VN_sign_out(11361),
        VN2CN4_sign => VN_sign_out(11362),
        VN2CN5_sign => VN_sign_out(11363),
        codeword => codeword(1893),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1894 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11369 downto 11364),
        Din0 => VN1894_in0,
        Din1 => VN1894_in1,
        Din2 => VN1894_in2,
        Din3 => VN1894_in3,
        Din4 => VN1894_in4,
        Din5 => VN1894_in5,
        VN2CN0_bit => VN_data_out(11364),
        VN2CN1_bit => VN_data_out(11365),
        VN2CN2_bit => VN_data_out(11366),
        VN2CN3_bit => VN_data_out(11367),
        VN2CN4_bit => VN_data_out(11368),
        VN2CN5_bit => VN_data_out(11369),
        VN2CN0_sign => VN_sign_out(11364),
        VN2CN1_sign => VN_sign_out(11365),
        VN2CN2_sign => VN_sign_out(11366),
        VN2CN3_sign => VN_sign_out(11367),
        VN2CN4_sign => VN_sign_out(11368),
        VN2CN5_sign => VN_sign_out(11369),
        codeword => codeword(1894),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1895 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11375 downto 11370),
        Din0 => VN1895_in0,
        Din1 => VN1895_in1,
        Din2 => VN1895_in2,
        Din3 => VN1895_in3,
        Din4 => VN1895_in4,
        Din5 => VN1895_in5,
        VN2CN0_bit => VN_data_out(11370),
        VN2CN1_bit => VN_data_out(11371),
        VN2CN2_bit => VN_data_out(11372),
        VN2CN3_bit => VN_data_out(11373),
        VN2CN4_bit => VN_data_out(11374),
        VN2CN5_bit => VN_data_out(11375),
        VN2CN0_sign => VN_sign_out(11370),
        VN2CN1_sign => VN_sign_out(11371),
        VN2CN2_sign => VN_sign_out(11372),
        VN2CN3_sign => VN_sign_out(11373),
        VN2CN4_sign => VN_sign_out(11374),
        VN2CN5_sign => VN_sign_out(11375),
        codeword => codeword(1895),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1896 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11381 downto 11376),
        Din0 => VN1896_in0,
        Din1 => VN1896_in1,
        Din2 => VN1896_in2,
        Din3 => VN1896_in3,
        Din4 => VN1896_in4,
        Din5 => VN1896_in5,
        VN2CN0_bit => VN_data_out(11376),
        VN2CN1_bit => VN_data_out(11377),
        VN2CN2_bit => VN_data_out(11378),
        VN2CN3_bit => VN_data_out(11379),
        VN2CN4_bit => VN_data_out(11380),
        VN2CN5_bit => VN_data_out(11381),
        VN2CN0_sign => VN_sign_out(11376),
        VN2CN1_sign => VN_sign_out(11377),
        VN2CN2_sign => VN_sign_out(11378),
        VN2CN3_sign => VN_sign_out(11379),
        VN2CN4_sign => VN_sign_out(11380),
        VN2CN5_sign => VN_sign_out(11381),
        codeword => codeword(1896),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1897 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11387 downto 11382),
        Din0 => VN1897_in0,
        Din1 => VN1897_in1,
        Din2 => VN1897_in2,
        Din3 => VN1897_in3,
        Din4 => VN1897_in4,
        Din5 => VN1897_in5,
        VN2CN0_bit => VN_data_out(11382),
        VN2CN1_bit => VN_data_out(11383),
        VN2CN2_bit => VN_data_out(11384),
        VN2CN3_bit => VN_data_out(11385),
        VN2CN4_bit => VN_data_out(11386),
        VN2CN5_bit => VN_data_out(11387),
        VN2CN0_sign => VN_sign_out(11382),
        VN2CN1_sign => VN_sign_out(11383),
        VN2CN2_sign => VN_sign_out(11384),
        VN2CN3_sign => VN_sign_out(11385),
        VN2CN4_sign => VN_sign_out(11386),
        VN2CN5_sign => VN_sign_out(11387),
        codeword => codeword(1897),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1898 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11393 downto 11388),
        Din0 => VN1898_in0,
        Din1 => VN1898_in1,
        Din2 => VN1898_in2,
        Din3 => VN1898_in3,
        Din4 => VN1898_in4,
        Din5 => VN1898_in5,
        VN2CN0_bit => VN_data_out(11388),
        VN2CN1_bit => VN_data_out(11389),
        VN2CN2_bit => VN_data_out(11390),
        VN2CN3_bit => VN_data_out(11391),
        VN2CN4_bit => VN_data_out(11392),
        VN2CN5_bit => VN_data_out(11393),
        VN2CN0_sign => VN_sign_out(11388),
        VN2CN1_sign => VN_sign_out(11389),
        VN2CN2_sign => VN_sign_out(11390),
        VN2CN3_sign => VN_sign_out(11391),
        VN2CN4_sign => VN_sign_out(11392),
        VN2CN5_sign => VN_sign_out(11393),
        codeword => codeword(1898),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1899 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11399 downto 11394),
        Din0 => VN1899_in0,
        Din1 => VN1899_in1,
        Din2 => VN1899_in2,
        Din3 => VN1899_in3,
        Din4 => VN1899_in4,
        Din5 => VN1899_in5,
        VN2CN0_bit => VN_data_out(11394),
        VN2CN1_bit => VN_data_out(11395),
        VN2CN2_bit => VN_data_out(11396),
        VN2CN3_bit => VN_data_out(11397),
        VN2CN4_bit => VN_data_out(11398),
        VN2CN5_bit => VN_data_out(11399),
        VN2CN0_sign => VN_sign_out(11394),
        VN2CN1_sign => VN_sign_out(11395),
        VN2CN2_sign => VN_sign_out(11396),
        VN2CN3_sign => VN_sign_out(11397),
        VN2CN4_sign => VN_sign_out(11398),
        VN2CN5_sign => VN_sign_out(11399),
        codeword => codeword(1899),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1900 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11405 downto 11400),
        Din0 => VN1900_in0,
        Din1 => VN1900_in1,
        Din2 => VN1900_in2,
        Din3 => VN1900_in3,
        Din4 => VN1900_in4,
        Din5 => VN1900_in5,
        VN2CN0_bit => VN_data_out(11400),
        VN2CN1_bit => VN_data_out(11401),
        VN2CN2_bit => VN_data_out(11402),
        VN2CN3_bit => VN_data_out(11403),
        VN2CN4_bit => VN_data_out(11404),
        VN2CN5_bit => VN_data_out(11405),
        VN2CN0_sign => VN_sign_out(11400),
        VN2CN1_sign => VN_sign_out(11401),
        VN2CN2_sign => VN_sign_out(11402),
        VN2CN3_sign => VN_sign_out(11403),
        VN2CN4_sign => VN_sign_out(11404),
        VN2CN5_sign => VN_sign_out(11405),
        codeword => codeword(1900),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1901 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11411 downto 11406),
        Din0 => VN1901_in0,
        Din1 => VN1901_in1,
        Din2 => VN1901_in2,
        Din3 => VN1901_in3,
        Din4 => VN1901_in4,
        Din5 => VN1901_in5,
        VN2CN0_bit => VN_data_out(11406),
        VN2CN1_bit => VN_data_out(11407),
        VN2CN2_bit => VN_data_out(11408),
        VN2CN3_bit => VN_data_out(11409),
        VN2CN4_bit => VN_data_out(11410),
        VN2CN5_bit => VN_data_out(11411),
        VN2CN0_sign => VN_sign_out(11406),
        VN2CN1_sign => VN_sign_out(11407),
        VN2CN2_sign => VN_sign_out(11408),
        VN2CN3_sign => VN_sign_out(11409),
        VN2CN4_sign => VN_sign_out(11410),
        VN2CN5_sign => VN_sign_out(11411),
        codeword => codeword(1901),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1902 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11417 downto 11412),
        Din0 => VN1902_in0,
        Din1 => VN1902_in1,
        Din2 => VN1902_in2,
        Din3 => VN1902_in3,
        Din4 => VN1902_in4,
        Din5 => VN1902_in5,
        VN2CN0_bit => VN_data_out(11412),
        VN2CN1_bit => VN_data_out(11413),
        VN2CN2_bit => VN_data_out(11414),
        VN2CN3_bit => VN_data_out(11415),
        VN2CN4_bit => VN_data_out(11416),
        VN2CN5_bit => VN_data_out(11417),
        VN2CN0_sign => VN_sign_out(11412),
        VN2CN1_sign => VN_sign_out(11413),
        VN2CN2_sign => VN_sign_out(11414),
        VN2CN3_sign => VN_sign_out(11415),
        VN2CN4_sign => VN_sign_out(11416),
        VN2CN5_sign => VN_sign_out(11417),
        codeword => codeword(1902),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1903 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11423 downto 11418),
        Din0 => VN1903_in0,
        Din1 => VN1903_in1,
        Din2 => VN1903_in2,
        Din3 => VN1903_in3,
        Din4 => VN1903_in4,
        Din5 => VN1903_in5,
        VN2CN0_bit => VN_data_out(11418),
        VN2CN1_bit => VN_data_out(11419),
        VN2CN2_bit => VN_data_out(11420),
        VN2CN3_bit => VN_data_out(11421),
        VN2CN4_bit => VN_data_out(11422),
        VN2CN5_bit => VN_data_out(11423),
        VN2CN0_sign => VN_sign_out(11418),
        VN2CN1_sign => VN_sign_out(11419),
        VN2CN2_sign => VN_sign_out(11420),
        VN2CN3_sign => VN_sign_out(11421),
        VN2CN4_sign => VN_sign_out(11422),
        VN2CN5_sign => VN_sign_out(11423),
        codeword => codeword(1903),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1904 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11429 downto 11424),
        Din0 => VN1904_in0,
        Din1 => VN1904_in1,
        Din2 => VN1904_in2,
        Din3 => VN1904_in3,
        Din4 => VN1904_in4,
        Din5 => VN1904_in5,
        VN2CN0_bit => VN_data_out(11424),
        VN2CN1_bit => VN_data_out(11425),
        VN2CN2_bit => VN_data_out(11426),
        VN2CN3_bit => VN_data_out(11427),
        VN2CN4_bit => VN_data_out(11428),
        VN2CN5_bit => VN_data_out(11429),
        VN2CN0_sign => VN_sign_out(11424),
        VN2CN1_sign => VN_sign_out(11425),
        VN2CN2_sign => VN_sign_out(11426),
        VN2CN3_sign => VN_sign_out(11427),
        VN2CN4_sign => VN_sign_out(11428),
        VN2CN5_sign => VN_sign_out(11429),
        codeword => codeword(1904),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1905 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11435 downto 11430),
        Din0 => VN1905_in0,
        Din1 => VN1905_in1,
        Din2 => VN1905_in2,
        Din3 => VN1905_in3,
        Din4 => VN1905_in4,
        Din5 => VN1905_in5,
        VN2CN0_bit => VN_data_out(11430),
        VN2CN1_bit => VN_data_out(11431),
        VN2CN2_bit => VN_data_out(11432),
        VN2CN3_bit => VN_data_out(11433),
        VN2CN4_bit => VN_data_out(11434),
        VN2CN5_bit => VN_data_out(11435),
        VN2CN0_sign => VN_sign_out(11430),
        VN2CN1_sign => VN_sign_out(11431),
        VN2CN2_sign => VN_sign_out(11432),
        VN2CN3_sign => VN_sign_out(11433),
        VN2CN4_sign => VN_sign_out(11434),
        VN2CN5_sign => VN_sign_out(11435),
        codeword => codeword(1905),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1906 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11441 downto 11436),
        Din0 => VN1906_in0,
        Din1 => VN1906_in1,
        Din2 => VN1906_in2,
        Din3 => VN1906_in3,
        Din4 => VN1906_in4,
        Din5 => VN1906_in5,
        VN2CN0_bit => VN_data_out(11436),
        VN2CN1_bit => VN_data_out(11437),
        VN2CN2_bit => VN_data_out(11438),
        VN2CN3_bit => VN_data_out(11439),
        VN2CN4_bit => VN_data_out(11440),
        VN2CN5_bit => VN_data_out(11441),
        VN2CN0_sign => VN_sign_out(11436),
        VN2CN1_sign => VN_sign_out(11437),
        VN2CN2_sign => VN_sign_out(11438),
        VN2CN3_sign => VN_sign_out(11439),
        VN2CN4_sign => VN_sign_out(11440),
        VN2CN5_sign => VN_sign_out(11441),
        codeword => codeword(1906),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1907 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11447 downto 11442),
        Din0 => VN1907_in0,
        Din1 => VN1907_in1,
        Din2 => VN1907_in2,
        Din3 => VN1907_in3,
        Din4 => VN1907_in4,
        Din5 => VN1907_in5,
        VN2CN0_bit => VN_data_out(11442),
        VN2CN1_bit => VN_data_out(11443),
        VN2CN2_bit => VN_data_out(11444),
        VN2CN3_bit => VN_data_out(11445),
        VN2CN4_bit => VN_data_out(11446),
        VN2CN5_bit => VN_data_out(11447),
        VN2CN0_sign => VN_sign_out(11442),
        VN2CN1_sign => VN_sign_out(11443),
        VN2CN2_sign => VN_sign_out(11444),
        VN2CN3_sign => VN_sign_out(11445),
        VN2CN4_sign => VN_sign_out(11446),
        VN2CN5_sign => VN_sign_out(11447),
        codeword => codeword(1907),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1908 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11453 downto 11448),
        Din0 => VN1908_in0,
        Din1 => VN1908_in1,
        Din2 => VN1908_in2,
        Din3 => VN1908_in3,
        Din4 => VN1908_in4,
        Din5 => VN1908_in5,
        VN2CN0_bit => VN_data_out(11448),
        VN2CN1_bit => VN_data_out(11449),
        VN2CN2_bit => VN_data_out(11450),
        VN2CN3_bit => VN_data_out(11451),
        VN2CN4_bit => VN_data_out(11452),
        VN2CN5_bit => VN_data_out(11453),
        VN2CN0_sign => VN_sign_out(11448),
        VN2CN1_sign => VN_sign_out(11449),
        VN2CN2_sign => VN_sign_out(11450),
        VN2CN3_sign => VN_sign_out(11451),
        VN2CN4_sign => VN_sign_out(11452),
        VN2CN5_sign => VN_sign_out(11453),
        codeword => codeword(1908),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1909 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11459 downto 11454),
        Din0 => VN1909_in0,
        Din1 => VN1909_in1,
        Din2 => VN1909_in2,
        Din3 => VN1909_in3,
        Din4 => VN1909_in4,
        Din5 => VN1909_in5,
        VN2CN0_bit => VN_data_out(11454),
        VN2CN1_bit => VN_data_out(11455),
        VN2CN2_bit => VN_data_out(11456),
        VN2CN3_bit => VN_data_out(11457),
        VN2CN4_bit => VN_data_out(11458),
        VN2CN5_bit => VN_data_out(11459),
        VN2CN0_sign => VN_sign_out(11454),
        VN2CN1_sign => VN_sign_out(11455),
        VN2CN2_sign => VN_sign_out(11456),
        VN2CN3_sign => VN_sign_out(11457),
        VN2CN4_sign => VN_sign_out(11458),
        VN2CN5_sign => VN_sign_out(11459),
        codeword => codeword(1909),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1910 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11465 downto 11460),
        Din0 => VN1910_in0,
        Din1 => VN1910_in1,
        Din2 => VN1910_in2,
        Din3 => VN1910_in3,
        Din4 => VN1910_in4,
        Din5 => VN1910_in5,
        VN2CN0_bit => VN_data_out(11460),
        VN2CN1_bit => VN_data_out(11461),
        VN2CN2_bit => VN_data_out(11462),
        VN2CN3_bit => VN_data_out(11463),
        VN2CN4_bit => VN_data_out(11464),
        VN2CN5_bit => VN_data_out(11465),
        VN2CN0_sign => VN_sign_out(11460),
        VN2CN1_sign => VN_sign_out(11461),
        VN2CN2_sign => VN_sign_out(11462),
        VN2CN3_sign => VN_sign_out(11463),
        VN2CN4_sign => VN_sign_out(11464),
        VN2CN5_sign => VN_sign_out(11465),
        codeword => codeword(1910),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1911 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11471 downto 11466),
        Din0 => VN1911_in0,
        Din1 => VN1911_in1,
        Din2 => VN1911_in2,
        Din3 => VN1911_in3,
        Din4 => VN1911_in4,
        Din5 => VN1911_in5,
        VN2CN0_bit => VN_data_out(11466),
        VN2CN1_bit => VN_data_out(11467),
        VN2CN2_bit => VN_data_out(11468),
        VN2CN3_bit => VN_data_out(11469),
        VN2CN4_bit => VN_data_out(11470),
        VN2CN5_bit => VN_data_out(11471),
        VN2CN0_sign => VN_sign_out(11466),
        VN2CN1_sign => VN_sign_out(11467),
        VN2CN2_sign => VN_sign_out(11468),
        VN2CN3_sign => VN_sign_out(11469),
        VN2CN4_sign => VN_sign_out(11470),
        VN2CN5_sign => VN_sign_out(11471),
        codeword => codeword(1911),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1912 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11477 downto 11472),
        Din0 => VN1912_in0,
        Din1 => VN1912_in1,
        Din2 => VN1912_in2,
        Din3 => VN1912_in3,
        Din4 => VN1912_in4,
        Din5 => VN1912_in5,
        VN2CN0_bit => VN_data_out(11472),
        VN2CN1_bit => VN_data_out(11473),
        VN2CN2_bit => VN_data_out(11474),
        VN2CN3_bit => VN_data_out(11475),
        VN2CN4_bit => VN_data_out(11476),
        VN2CN5_bit => VN_data_out(11477),
        VN2CN0_sign => VN_sign_out(11472),
        VN2CN1_sign => VN_sign_out(11473),
        VN2CN2_sign => VN_sign_out(11474),
        VN2CN3_sign => VN_sign_out(11475),
        VN2CN4_sign => VN_sign_out(11476),
        VN2CN5_sign => VN_sign_out(11477),
        codeword => codeword(1912),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1913 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11483 downto 11478),
        Din0 => VN1913_in0,
        Din1 => VN1913_in1,
        Din2 => VN1913_in2,
        Din3 => VN1913_in3,
        Din4 => VN1913_in4,
        Din5 => VN1913_in5,
        VN2CN0_bit => VN_data_out(11478),
        VN2CN1_bit => VN_data_out(11479),
        VN2CN2_bit => VN_data_out(11480),
        VN2CN3_bit => VN_data_out(11481),
        VN2CN4_bit => VN_data_out(11482),
        VN2CN5_bit => VN_data_out(11483),
        VN2CN0_sign => VN_sign_out(11478),
        VN2CN1_sign => VN_sign_out(11479),
        VN2CN2_sign => VN_sign_out(11480),
        VN2CN3_sign => VN_sign_out(11481),
        VN2CN4_sign => VN_sign_out(11482),
        VN2CN5_sign => VN_sign_out(11483),
        codeword => codeword(1913),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1914 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11489 downto 11484),
        Din0 => VN1914_in0,
        Din1 => VN1914_in1,
        Din2 => VN1914_in2,
        Din3 => VN1914_in3,
        Din4 => VN1914_in4,
        Din5 => VN1914_in5,
        VN2CN0_bit => VN_data_out(11484),
        VN2CN1_bit => VN_data_out(11485),
        VN2CN2_bit => VN_data_out(11486),
        VN2CN3_bit => VN_data_out(11487),
        VN2CN4_bit => VN_data_out(11488),
        VN2CN5_bit => VN_data_out(11489),
        VN2CN0_sign => VN_sign_out(11484),
        VN2CN1_sign => VN_sign_out(11485),
        VN2CN2_sign => VN_sign_out(11486),
        VN2CN3_sign => VN_sign_out(11487),
        VN2CN4_sign => VN_sign_out(11488),
        VN2CN5_sign => VN_sign_out(11489),
        codeword => codeword(1914),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1915 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11495 downto 11490),
        Din0 => VN1915_in0,
        Din1 => VN1915_in1,
        Din2 => VN1915_in2,
        Din3 => VN1915_in3,
        Din4 => VN1915_in4,
        Din5 => VN1915_in5,
        VN2CN0_bit => VN_data_out(11490),
        VN2CN1_bit => VN_data_out(11491),
        VN2CN2_bit => VN_data_out(11492),
        VN2CN3_bit => VN_data_out(11493),
        VN2CN4_bit => VN_data_out(11494),
        VN2CN5_bit => VN_data_out(11495),
        VN2CN0_sign => VN_sign_out(11490),
        VN2CN1_sign => VN_sign_out(11491),
        VN2CN2_sign => VN_sign_out(11492),
        VN2CN3_sign => VN_sign_out(11493),
        VN2CN4_sign => VN_sign_out(11494),
        VN2CN5_sign => VN_sign_out(11495),
        codeword => codeword(1915),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1916 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11501 downto 11496),
        Din0 => VN1916_in0,
        Din1 => VN1916_in1,
        Din2 => VN1916_in2,
        Din3 => VN1916_in3,
        Din4 => VN1916_in4,
        Din5 => VN1916_in5,
        VN2CN0_bit => VN_data_out(11496),
        VN2CN1_bit => VN_data_out(11497),
        VN2CN2_bit => VN_data_out(11498),
        VN2CN3_bit => VN_data_out(11499),
        VN2CN4_bit => VN_data_out(11500),
        VN2CN5_bit => VN_data_out(11501),
        VN2CN0_sign => VN_sign_out(11496),
        VN2CN1_sign => VN_sign_out(11497),
        VN2CN2_sign => VN_sign_out(11498),
        VN2CN3_sign => VN_sign_out(11499),
        VN2CN4_sign => VN_sign_out(11500),
        VN2CN5_sign => VN_sign_out(11501),
        codeword => codeword(1916),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1917 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11507 downto 11502),
        Din0 => VN1917_in0,
        Din1 => VN1917_in1,
        Din2 => VN1917_in2,
        Din3 => VN1917_in3,
        Din4 => VN1917_in4,
        Din5 => VN1917_in5,
        VN2CN0_bit => VN_data_out(11502),
        VN2CN1_bit => VN_data_out(11503),
        VN2CN2_bit => VN_data_out(11504),
        VN2CN3_bit => VN_data_out(11505),
        VN2CN4_bit => VN_data_out(11506),
        VN2CN5_bit => VN_data_out(11507),
        VN2CN0_sign => VN_sign_out(11502),
        VN2CN1_sign => VN_sign_out(11503),
        VN2CN2_sign => VN_sign_out(11504),
        VN2CN3_sign => VN_sign_out(11505),
        VN2CN4_sign => VN_sign_out(11506),
        VN2CN5_sign => VN_sign_out(11507),
        codeword => codeword(1917),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1918 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11513 downto 11508),
        Din0 => VN1918_in0,
        Din1 => VN1918_in1,
        Din2 => VN1918_in2,
        Din3 => VN1918_in3,
        Din4 => VN1918_in4,
        Din5 => VN1918_in5,
        VN2CN0_bit => VN_data_out(11508),
        VN2CN1_bit => VN_data_out(11509),
        VN2CN2_bit => VN_data_out(11510),
        VN2CN3_bit => VN_data_out(11511),
        VN2CN4_bit => VN_data_out(11512),
        VN2CN5_bit => VN_data_out(11513),
        VN2CN0_sign => VN_sign_out(11508),
        VN2CN1_sign => VN_sign_out(11509),
        VN2CN2_sign => VN_sign_out(11510),
        VN2CN3_sign => VN_sign_out(11511),
        VN2CN4_sign => VN_sign_out(11512),
        VN2CN5_sign => VN_sign_out(11513),
        codeword => codeword(1918),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1919 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11519 downto 11514),
        Din0 => VN1919_in0,
        Din1 => VN1919_in1,
        Din2 => VN1919_in2,
        Din3 => VN1919_in3,
        Din4 => VN1919_in4,
        Din5 => VN1919_in5,
        VN2CN0_bit => VN_data_out(11514),
        VN2CN1_bit => VN_data_out(11515),
        VN2CN2_bit => VN_data_out(11516),
        VN2CN3_bit => VN_data_out(11517),
        VN2CN4_bit => VN_data_out(11518),
        VN2CN5_bit => VN_data_out(11519),
        VN2CN0_sign => VN_sign_out(11514),
        VN2CN1_sign => VN_sign_out(11515),
        VN2CN2_sign => VN_sign_out(11516),
        VN2CN3_sign => VN_sign_out(11517),
        VN2CN4_sign => VN_sign_out(11518),
        VN2CN5_sign => VN_sign_out(11519),
        codeword => codeword(1919),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1920 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11525 downto 11520),
        Din0 => VN1920_in0,
        Din1 => VN1920_in1,
        Din2 => VN1920_in2,
        Din3 => VN1920_in3,
        Din4 => VN1920_in4,
        Din5 => VN1920_in5,
        VN2CN0_bit => VN_data_out(11520),
        VN2CN1_bit => VN_data_out(11521),
        VN2CN2_bit => VN_data_out(11522),
        VN2CN3_bit => VN_data_out(11523),
        VN2CN4_bit => VN_data_out(11524),
        VN2CN5_bit => VN_data_out(11525),
        VN2CN0_sign => VN_sign_out(11520),
        VN2CN1_sign => VN_sign_out(11521),
        VN2CN2_sign => VN_sign_out(11522),
        VN2CN3_sign => VN_sign_out(11523),
        VN2CN4_sign => VN_sign_out(11524),
        VN2CN5_sign => VN_sign_out(11525),
        codeword => codeword(1920),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1921 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11531 downto 11526),
        Din0 => VN1921_in0,
        Din1 => VN1921_in1,
        Din2 => VN1921_in2,
        Din3 => VN1921_in3,
        Din4 => VN1921_in4,
        Din5 => VN1921_in5,
        VN2CN0_bit => VN_data_out(11526),
        VN2CN1_bit => VN_data_out(11527),
        VN2CN2_bit => VN_data_out(11528),
        VN2CN3_bit => VN_data_out(11529),
        VN2CN4_bit => VN_data_out(11530),
        VN2CN5_bit => VN_data_out(11531),
        VN2CN0_sign => VN_sign_out(11526),
        VN2CN1_sign => VN_sign_out(11527),
        VN2CN2_sign => VN_sign_out(11528),
        VN2CN3_sign => VN_sign_out(11529),
        VN2CN4_sign => VN_sign_out(11530),
        VN2CN5_sign => VN_sign_out(11531),
        codeword => codeword(1921),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1922 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11537 downto 11532),
        Din0 => VN1922_in0,
        Din1 => VN1922_in1,
        Din2 => VN1922_in2,
        Din3 => VN1922_in3,
        Din4 => VN1922_in4,
        Din5 => VN1922_in5,
        VN2CN0_bit => VN_data_out(11532),
        VN2CN1_bit => VN_data_out(11533),
        VN2CN2_bit => VN_data_out(11534),
        VN2CN3_bit => VN_data_out(11535),
        VN2CN4_bit => VN_data_out(11536),
        VN2CN5_bit => VN_data_out(11537),
        VN2CN0_sign => VN_sign_out(11532),
        VN2CN1_sign => VN_sign_out(11533),
        VN2CN2_sign => VN_sign_out(11534),
        VN2CN3_sign => VN_sign_out(11535),
        VN2CN4_sign => VN_sign_out(11536),
        VN2CN5_sign => VN_sign_out(11537),
        codeword => codeword(1922),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1923 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11543 downto 11538),
        Din0 => VN1923_in0,
        Din1 => VN1923_in1,
        Din2 => VN1923_in2,
        Din3 => VN1923_in3,
        Din4 => VN1923_in4,
        Din5 => VN1923_in5,
        VN2CN0_bit => VN_data_out(11538),
        VN2CN1_bit => VN_data_out(11539),
        VN2CN2_bit => VN_data_out(11540),
        VN2CN3_bit => VN_data_out(11541),
        VN2CN4_bit => VN_data_out(11542),
        VN2CN5_bit => VN_data_out(11543),
        VN2CN0_sign => VN_sign_out(11538),
        VN2CN1_sign => VN_sign_out(11539),
        VN2CN2_sign => VN_sign_out(11540),
        VN2CN3_sign => VN_sign_out(11541),
        VN2CN4_sign => VN_sign_out(11542),
        VN2CN5_sign => VN_sign_out(11543),
        codeword => codeword(1923),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1924 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11549 downto 11544),
        Din0 => VN1924_in0,
        Din1 => VN1924_in1,
        Din2 => VN1924_in2,
        Din3 => VN1924_in3,
        Din4 => VN1924_in4,
        Din5 => VN1924_in5,
        VN2CN0_bit => VN_data_out(11544),
        VN2CN1_bit => VN_data_out(11545),
        VN2CN2_bit => VN_data_out(11546),
        VN2CN3_bit => VN_data_out(11547),
        VN2CN4_bit => VN_data_out(11548),
        VN2CN5_bit => VN_data_out(11549),
        VN2CN0_sign => VN_sign_out(11544),
        VN2CN1_sign => VN_sign_out(11545),
        VN2CN2_sign => VN_sign_out(11546),
        VN2CN3_sign => VN_sign_out(11547),
        VN2CN4_sign => VN_sign_out(11548),
        VN2CN5_sign => VN_sign_out(11549),
        codeword => codeword(1924),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1925 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11555 downto 11550),
        Din0 => VN1925_in0,
        Din1 => VN1925_in1,
        Din2 => VN1925_in2,
        Din3 => VN1925_in3,
        Din4 => VN1925_in4,
        Din5 => VN1925_in5,
        VN2CN0_bit => VN_data_out(11550),
        VN2CN1_bit => VN_data_out(11551),
        VN2CN2_bit => VN_data_out(11552),
        VN2CN3_bit => VN_data_out(11553),
        VN2CN4_bit => VN_data_out(11554),
        VN2CN5_bit => VN_data_out(11555),
        VN2CN0_sign => VN_sign_out(11550),
        VN2CN1_sign => VN_sign_out(11551),
        VN2CN2_sign => VN_sign_out(11552),
        VN2CN3_sign => VN_sign_out(11553),
        VN2CN4_sign => VN_sign_out(11554),
        VN2CN5_sign => VN_sign_out(11555),
        codeword => codeword(1925),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1926 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11561 downto 11556),
        Din0 => VN1926_in0,
        Din1 => VN1926_in1,
        Din2 => VN1926_in2,
        Din3 => VN1926_in3,
        Din4 => VN1926_in4,
        Din5 => VN1926_in5,
        VN2CN0_bit => VN_data_out(11556),
        VN2CN1_bit => VN_data_out(11557),
        VN2CN2_bit => VN_data_out(11558),
        VN2CN3_bit => VN_data_out(11559),
        VN2CN4_bit => VN_data_out(11560),
        VN2CN5_bit => VN_data_out(11561),
        VN2CN0_sign => VN_sign_out(11556),
        VN2CN1_sign => VN_sign_out(11557),
        VN2CN2_sign => VN_sign_out(11558),
        VN2CN3_sign => VN_sign_out(11559),
        VN2CN4_sign => VN_sign_out(11560),
        VN2CN5_sign => VN_sign_out(11561),
        codeword => codeword(1926),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1927 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11567 downto 11562),
        Din0 => VN1927_in0,
        Din1 => VN1927_in1,
        Din2 => VN1927_in2,
        Din3 => VN1927_in3,
        Din4 => VN1927_in4,
        Din5 => VN1927_in5,
        VN2CN0_bit => VN_data_out(11562),
        VN2CN1_bit => VN_data_out(11563),
        VN2CN2_bit => VN_data_out(11564),
        VN2CN3_bit => VN_data_out(11565),
        VN2CN4_bit => VN_data_out(11566),
        VN2CN5_bit => VN_data_out(11567),
        VN2CN0_sign => VN_sign_out(11562),
        VN2CN1_sign => VN_sign_out(11563),
        VN2CN2_sign => VN_sign_out(11564),
        VN2CN3_sign => VN_sign_out(11565),
        VN2CN4_sign => VN_sign_out(11566),
        VN2CN5_sign => VN_sign_out(11567),
        codeword => codeword(1927),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1928 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11573 downto 11568),
        Din0 => VN1928_in0,
        Din1 => VN1928_in1,
        Din2 => VN1928_in2,
        Din3 => VN1928_in3,
        Din4 => VN1928_in4,
        Din5 => VN1928_in5,
        VN2CN0_bit => VN_data_out(11568),
        VN2CN1_bit => VN_data_out(11569),
        VN2CN2_bit => VN_data_out(11570),
        VN2CN3_bit => VN_data_out(11571),
        VN2CN4_bit => VN_data_out(11572),
        VN2CN5_bit => VN_data_out(11573),
        VN2CN0_sign => VN_sign_out(11568),
        VN2CN1_sign => VN_sign_out(11569),
        VN2CN2_sign => VN_sign_out(11570),
        VN2CN3_sign => VN_sign_out(11571),
        VN2CN4_sign => VN_sign_out(11572),
        VN2CN5_sign => VN_sign_out(11573),
        codeword => codeword(1928),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1929 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11579 downto 11574),
        Din0 => VN1929_in0,
        Din1 => VN1929_in1,
        Din2 => VN1929_in2,
        Din3 => VN1929_in3,
        Din4 => VN1929_in4,
        Din5 => VN1929_in5,
        VN2CN0_bit => VN_data_out(11574),
        VN2CN1_bit => VN_data_out(11575),
        VN2CN2_bit => VN_data_out(11576),
        VN2CN3_bit => VN_data_out(11577),
        VN2CN4_bit => VN_data_out(11578),
        VN2CN5_bit => VN_data_out(11579),
        VN2CN0_sign => VN_sign_out(11574),
        VN2CN1_sign => VN_sign_out(11575),
        VN2CN2_sign => VN_sign_out(11576),
        VN2CN3_sign => VN_sign_out(11577),
        VN2CN4_sign => VN_sign_out(11578),
        VN2CN5_sign => VN_sign_out(11579),
        codeword => codeword(1929),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1930 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11585 downto 11580),
        Din0 => VN1930_in0,
        Din1 => VN1930_in1,
        Din2 => VN1930_in2,
        Din3 => VN1930_in3,
        Din4 => VN1930_in4,
        Din5 => VN1930_in5,
        VN2CN0_bit => VN_data_out(11580),
        VN2CN1_bit => VN_data_out(11581),
        VN2CN2_bit => VN_data_out(11582),
        VN2CN3_bit => VN_data_out(11583),
        VN2CN4_bit => VN_data_out(11584),
        VN2CN5_bit => VN_data_out(11585),
        VN2CN0_sign => VN_sign_out(11580),
        VN2CN1_sign => VN_sign_out(11581),
        VN2CN2_sign => VN_sign_out(11582),
        VN2CN3_sign => VN_sign_out(11583),
        VN2CN4_sign => VN_sign_out(11584),
        VN2CN5_sign => VN_sign_out(11585),
        codeword => codeword(1930),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1931 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11591 downto 11586),
        Din0 => VN1931_in0,
        Din1 => VN1931_in1,
        Din2 => VN1931_in2,
        Din3 => VN1931_in3,
        Din4 => VN1931_in4,
        Din5 => VN1931_in5,
        VN2CN0_bit => VN_data_out(11586),
        VN2CN1_bit => VN_data_out(11587),
        VN2CN2_bit => VN_data_out(11588),
        VN2CN3_bit => VN_data_out(11589),
        VN2CN4_bit => VN_data_out(11590),
        VN2CN5_bit => VN_data_out(11591),
        VN2CN0_sign => VN_sign_out(11586),
        VN2CN1_sign => VN_sign_out(11587),
        VN2CN2_sign => VN_sign_out(11588),
        VN2CN3_sign => VN_sign_out(11589),
        VN2CN4_sign => VN_sign_out(11590),
        VN2CN5_sign => VN_sign_out(11591),
        codeword => codeword(1931),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1932 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11597 downto 11592),
        Din0 => VN1932_in0,
        Din1 => VN1932_in1,
        Din2 => VN1932_in2,
        Din3 => VN1932_in3,
        Din4 => VN1932_in4,
        Din5 => VN1932_in5,
        VN2CN0_bit => VN_data_out(11592),
        VN2CN1_bit => VN_data_out(11593),
        VN2CN2_bit => VN_data_out(11594),
        VN2CN3_bit => VN_data_out(11595),
        VN2CN4_bit => VN_data_out(11596),
        VN2CN5_bit => VN_data_out(11597),
        VN2CN0_sign => VN_sign_out(11592),
        VN2CN1_sign => VN_sign_out(11593),
        VN2CN2_sign => VN_sign_out(11594),
        VN2CN3_sign => VN_sign_out(11595),
        VN2CN4_sign => VN_sign_out(11596),
        VN2CN5_sign => VN_sign_out(11597),
        codeword => codeword(1932),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1933 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11603 downto 11598),
        Din0 => VN1933_in0,
        Din1 => VN1933_in1,
        Din2 => VN1933_in2,
        Din3 => VN1933_in3,
        Din4 => VN1933_in4,
        Din5 => VN1933_in5,
        VN2CN0_bit => VN_data_out(11598),
        VN2CN1_bit => VN_data_out(11599),
        VN2CN2_bit => VN_data_out(11600),
        VN2CN3_bit => VN_data_out(11601),
        VN2CN4_bit => VN_data_out(11602),
        VN2CN5_bit => VN_data_out(11603),
        VN2CN0_sign => VN_sign_out(11598),
        VN2CN1_sign => VN_sign_out(11599),
        VN2CN2_sign => VN_sign_out(11600),
        VN2CN3_sign => VN_sign_out(11601),
        VN2CN4_sign => VN_sign_out(11602),
        VN2CN5_sign => VN_sign_out(11603),
        codeword => codeword(1933),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1934 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11609 downto 11604),
        Din0 => VN1934_in0,
        Din1 => VN1934_in1,
        Din2 => VN1934_in2,
        Din3 => VN1934_in3,
        Din4 => VN1934_in4,
        Din5 => VN1934_in5,
        VN2CN0_bit => VN_data_out(11604),
        VN2CN1_bit => VN_data_out(11605),
        VN2CN2_bit => VN_data_out(11606),
        VN2CN3_bit => VN_data_out(11607),
        VN2CN4_bit => VN_data_out(11608),
        VN2CN5_bit => VN_data_out(11609),
        VN2CN0_sign => VN_sign_out(11604),
        VN2CN1_sign => VN_sign_out(11605),
        VN2CN2_sign => VN_sign_out(11606),
        VN2CN3_sign => VN_sign_out(11607),
        VN2CN4_sign => VN_sign_out(11608),
        VN2CN5_sign => VN_sign_out(11609),
        codeword => codeword(1934),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1935 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11615 downto 11610),
        Din0 => VN1935_in0,
        Din1 => VN1935_in1,
        Din2 => VN1935_in2,
        Din3 => VN1935_in3,
        Din4 => VN1935_in4,
        Din5 => VN1935_in5,
        VN2CN0_bit => VN_data_out(11610),
        VN2CN1_bit => VN_data_out(11611),
        VN2CN2_bit => VN_data_out(11612),
        VN2CN3_bit => VN_data_out(11613),
        VN2CN4_bit => VN_data_out(11614),
        VN2CN5_bit => VN_data_out(11615),
        VN2CN0_sign => VN_sign_out(11610),
        VN2CN1_sign => VN_sign_out(11611),
        VN2CN2_sign => VN_sign_out(11612),
        VN2CN3_sign => VN_sign_out(11613),
        VN2CN4_sign => VN_sign_out(11614),
        VN2CN5_sign => VN_sign_out(11615),
        codeword => codeword(1935),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1936 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11621 downto 11616),
        Din0 => VN1936_in0,
        Din1 => VN1936_in1,
        Din2 => VN1936_in2,
        Din3 => VN1936_in3,
        Din4 => VN1936_in4,
        Din5 => VN1936_in5,
        VN2CN0_bit => VN_data_out(11616),
        VN2CN1_bit => VN_data_out(11617),
        VN2CN2_bit => VN_data_out(11618),
        VN2CN3_bit => VN_data_out(11619),
        VN2CN4_bit => VN_data_out(11620),
        VN2CN5_bit => VN_data_out(11621),
        VN2CN0_sign => VN_sign_out(11616),
        VN2CN1_sign => VN_sign_out(11617),
        VN2CN2_sign => VN_sign_out(11618),
        VN2CN3_sign => VN_sign_out(11619),
        VN2CN4_sign => VN_sign_out(11620),
        VN2CN5_sign => VN_sign_out(11621),
        codeword => codeword(1936),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1937 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11627 downto 11622),
        Din0 => VN1937_in0,
        Din1 => VN1937_in1,
        Din2 => VN1937_in2,
        Din3 => VN1937_in3,
        Din4 => VN1937_in4,
        Din5 => VN1937_in5,
        VN2CN0_bit => VN_data_out(11622),
        VN2CN1_bit => VN_data_out(11623),
        VN2CN2_bit => VN_data_out(11624),
        VN2CN3_bit => VN_data_out(11625),
        VN2CN4_bit => VN_data_out(11626),
        VN2CN5_bit => VN_data_out(11627),
        VN2CN0_sign => VN_sign_out(11622),
        VN2CN1_sign => VN_sign_out(11623),
        VN2CN2_sign => VN_sign_out(11624),
        VN2CN3_sign => VN_sign_out(11625),
        VN2CN4_sign => VN_sign_out(11626),
        VN2CN5_sign => VN_sign_out(11627),
        codeword => codeword(1937),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1938 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11633 downto 11628),
        Din0 => VN1938_in0,
        Din1 => VN1938_in1,
        Din2 => VN1938_in2,
        Din3 => VN1938_in3,
        Din4 => VN1938_in4,
        Din5 => VN1938_in5,
        VN2CN0_bit => VN_data_out(11628),
        VN2CN1_bit => VN_data_out(11629),
        VN2CN2_bit => VN_data_out(11630),
        VN2CN3_bit => VN_data_out(11631),
        VN2CN4_bit => VN_data_out(11632),
        VN2CN5_bit => VN_data_out(11633),
        VN2CN0_sign => VN_sign_out(11628),
        VN2CN1_sign => VN_sign_out(11629),
        VN2CN2_sign => VN_sign_out(11630),
        VN2CN3_sign => VN_sign_out(11631),
        VN2CN4_sign => VN_sign_out(11632),
        VN2CN5_sign => VN_sign_out(11633),
        codeword => codeword(1938),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1939 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11639 downto 11634),
        Din0 => VN1939_in0,
        Din1 => VN1939_in1,
        Din2 => VN1939_in2,
        Din3 => VN1939_in3,
        Din4 => VN1939_in4,
        Din5 => VN1939_in5,
        VN2CN0_bit => VN_data_out(11634),
        VN2CN1_bit => VN_data_out(11635),
        VN2CN2_bit => VN_data_out(11636),
        VN2CN3_bit => VN_data_out(11637),
        VN2CN4_bit => VN_data_out(11638),
        VN2CN5_bit => VN_data_out(11639),
        VN2CN0_sign => VN_sign_out(11634),
        VN2CN1_sign => VN_sign_out(11635),
        VN2CN2_sign => VN_sign_out(11636),
        VN2CN3_sign => VN_sign_out(11637),
        VN2CN4_sign => VN_sign_out(11638),
        VN2CN5_sign => VN_sign_out(11639),
        codeword => codeword(1939),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1940 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11645 downto 11640),
        Din0 => VN1940_in0,
        Din1 => VN1940_in1,
        Din2 => VN1940_in2,
        Din3 => VN1940_in3,
        Din4 => VN1940_in4,
        Din5 => VN1940_in5,
        VN2CN0_bit => VN_data_out(11640),
        VN2CN1_bit => VN_data_out(11641),
        VN2CN2_bit => VN_data_out(11642),
        VN2CN3_bit => VN_data_out(11643),
        VN2CN4_bit => VN_data_out(11644),
        VN2CN5_bit => VN_data_out(11645),
        VN2CN0_sign => VN_sign_out(11640),
        VN2CN1_sign => VN_sign_out(11641),
        VN2CN2_sign => VN_sign_out(11642),
        VN2CN3_sign => VN_sign_out(11643),
        VN2CN4_sign => VN_sign_out(11644),
        VN2CN5_sign => VN_sign_out(11645),
        codeword => codeword(1940),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1941 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11651 downto 11646),
        Din0 => VN1941_in0,
        Din1 => VN1941_in1,
        Din2 => VN1941_in2,
        Din3 => VN1941_in3,
        Din4 => VN1941_in4,
        Din5 => VN1941_in5,
        VN2CN0_bit => VN_data_out(11646),
        VN2CN1_bit => VN_data_out(11647),
        VN2CN2_bit => VN_data_out(11648),
        VN2CN3_bit => VN_data_out(11649),
        VN2CN4_bit => VN_data_out(11650),
        VN2CN5_bit => VN_data_out(11651),
        VN2CN0_sign => VN_sign_out(11646),
        VN2CN1_sign => VN_sign_out(11647),
        VN2CN2_sign => VN_sign_out(11648),
        VN2CN3_sign => VN_sign_out(11649),
        VN2CN4_sign => VN_sign_out(11650),
        VN2CN5_sign => VN_sign_out(11651),
        codeword => codeword(1941),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1942 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11657 downto 11652),
        Din0 => VN1942_in0,
        Din1 => VN1942_in1,
        Din2 => VN1942_in2,
        Din3 => VN1942_in3,
        Din4 => VN1942_in4,
        Din5 => VN1942_in5,
        VN2CN0_bit => VN_data_out(11652),
        VN2CN1_bit => VN_data_out(11653),
        VN2CN2_bit => VN_data_out(11654),
        VN2CN3_bit => VN_data_out(11655),
        VN2CN4_bit => VN_data_out(11656),
        VN2CN5_bit => VN_data_out(11657),
        VN2CN0_sign => VN_sign_out(11652),
        VN2CN1_sign => VN_sign_out(11653),
        VN2CN2_sign => VN_sign_out(11654),
        VN2CN3_sign => VN_sign_out(11655),
        VN2CN4_sign => VN_sign_out(11656),
        VN2CN5_sign => VN_sign_out(11657),
        codeword => codeword(1942),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1943 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11663 downto 11658),
        Din0 => VN1943_in0,
        Din1 => VN1943_in1,
        Din2 => VN1943_in2,
        Din3 => VN1943_in3,
        Din4 => VN1943_in4,
        Din5 => VN1943_in5,
        VN2CN0_bit => VN_data_out(11658),
        VN2CN1_bit => VN_data_out(11659),
        VN2CN2_bit => VN_data_out(11660),
        VN2CN3_bit => VN_data_out(11661),
        VN2CN4_bit => VN_data_out(11662),
        VN2CN5_bit => VN_data_out(11663),
        VN2CN0_sign => VN_sign_out(11658),
        VN2CN1_sign => VN_sign_out(11659),
        VN2CN2_sign => VN_sign_out(11660),
        VN2CN3_sign => VN_sign_out(11661),
        VN2CN4_sign => VN_sign_out(11662),
        VN2CN5_sign => VN_sign_out(11663),
        codeword => codeword(1943),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1944 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11669 downto 11664),
        Din0 => VN1944_in0,
        Din1 => VN1944_in1,
        Din2 => VN1944_in2,
        Din3 => VN1944_in3,
        Din4 => VN1944_in4,
        Din5 => VN1944_in5,
        VN2CN0_bit => VN_data_out(11664),
        VN2CN1_bit => VN_data_out(11665),
        VN2CN2_bit => VN_data_out(11666),
        VN2CN3_bit => VN_data_out(11667),
        VN2CN4_bit => VN_data_out(11668),
        VN2CN5_bit => VN_data_out(11669),
        VN2CN0_sign => VN_sign_out(11664),
        VN2CN1_sign => VN_sign_out(11665),
        VN2CN2_sign => VN_sign_out(11666),
        VN2CN3_sign => VN_sign_out(11667),
        VN2CN4_sign => VN_sign_out(11668),
        VN2CN5_sign => VN_sign_out(11669),
        codeword => codeword(1944),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1945 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11675 downto 11670),
        Din0 => VN1945_in0,
        Din1 => VN1945_in1,
        Din2 => VN1945_in2,
        Din3 => VN1945_in3,
        Din4 => VN1945_in4,
        Din5 => VN1945_in5,
        VN2CN0_bit => VN_data_out(11670),
        VN2CN1_bit => VN_data_out(11671),
        VN2CN2_bit => VN_data_out(11672),
        VN2CN3_bit => VN_data_out(11673),
        VN2CN4_bit => VN_data_out(11674),
        VN2CN5_bit => VN_data_out(11675),
        VN2CN0_sign => VN_sign_out(11670),
        VN2CN1_sign => VN_sign_out(11671),
        VN2CN2_sign => VN_sign_out(11672),
        VN2CN3_sign => VN_sign_out(11673),
        VN2CN4_sign => VN_sign_out(11674),
        VN2CN5_sign => VN_sign_out(11675),
        codeword => codeword(1945),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1946 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11681 downto 11676),
        Din0 => VN1946_in0,
        Din1 => VN1946_in1,
        Din2 => VN1946_in2,
        Din3 => VN1946_in3,
        Din4 => VN1946_in4,
        Din5 => VN1946_in5,
        VN2CN0_bit => VN_data_out(11676),
        VN2CN1_bit => VN_data_out(11677),
        VN2CN2_bit => VN_data_out(11678),
        VN2CN3_bit => VN_data_out(11679),
        VN2CN4_bit => VN_data_out(11680),
        VN2CN5_bit => VN_data_out(11681),
        VN2CN0_sign => VN_sign_out(11676),
        VN2CN1_sign => VN_sign_out(11677),
        VN2CN2_sign => VN_sign_out(11678),
        VN2CN3_sign => VN_sign_out(11679),
        VN2CN4_sign => VN_sign_out(11680),
        VN2CN5_sign => VN_sign_out(11681),
        codeword => codeword(1946),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1947 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11687 downto 11682),
        Din0 => VN1947_in0,
        Din1 => VN1947_in1,
        Din2 => VN1947_in2,
        Din3 => VN1947_in3,
        Din4 => VN1947_in4,
        Din5 => VN1947_in5,
        VN2CN0_bit => VN_data_out(11682),
        VN2CN1_bit => VN_data_out(11683),
        VN2CN2_bit => VN_data_out(11684),
        VN2CN3_bit => VN_data_out(11685),
        VN2CN4_bit => VN_data_out(11686),
        VN2CN5_bit => VN_data_out(11687),
        VN2CN0_sign => VN_sign_out(11682),
        VN2CN1_sign => VN_sign_out(11683),
        VN2CN2_sign => VN_sign_out(11684),
        VN2CN3_sign => VN_sign_out(11685),
        VN2CN4_sign => VN_sign_out(11686),
        VN2CN5_sign => VN_sign_out(11687),
        codeword => codeword(1947),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1948 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11693 downto 11688),
        Din0 => VN1948_in0,
        Din1 => VN1948_in1,
        Din2 => VN1948_in2,
        Din3 => VN1948_in3,
        Din4 => VN1948_in4,
        Din5 => VN1948_in5,
        VN2CN0_bit => VN_data_out(11688),
        VN2CN1_bit => VN_data_out(11689),
        VN2CN2_bit => VN_data_out(11690),
        VN2CN3_bit => VN_data_out(11691),
        VN2CN4_bit => VN_data_out(11692),
        VN2CN5_bit => VN_data_out(11693),
        VN2CN0_sign => VN_sign_out(11688),
        VN2CN1_sign => VN_sign_out(11689),
        VN2CN2_sign => VN_sign_out(11690),
        VN2CN3_sign => VN_sign_out(11691),
        VN2CN4_sign => VN_sign_out(11692),
        VN2CN5_sign => VN_sign_out(11693),
        codeword => codeword(1948),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1949 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11699 downto 11694),
        Din0 => VN1949_in0,
        Din1 => VN1949_in1,
        Din2 => VN1949_in2,
        Din3 => VN1949_in3,
        Din4 => VN1949_in4,
        Din5 => VN1949_in5,
        VN2CN0_bit => VN_data_out(11694),
        VN2CN1_bit => VN_data_out(11695),
        VN2CN2_bit => VN_data_out(11696),
        VN2CN3_bit => VN_data_out(11697),
        VN2CN4_bit => VN_data_out(11698),
        VN2CN5_bit => VN_data_out(11699),
        VN2CN0_sign => VN_sign_out(11694),
        VN2CN1_sign => VN_sign_out(11695),
        VN2CN2_sign => VN_sign_out(11696),
        VN2CN3_sign => VN_sign_out(11697),
        VN2CN4_sign => VN_sign_out(11698),
        VN2CN5_sign => VN_sign_out(11699),
        codeword => codeword(1949),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1950 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11705 downto 11700),
        Din0 => VN1950_in0,
        Din1 => VN1950_in1,
        Din2 => VN1950_in2,
        Din3 => VN1950_in3,
        Din4 => VN1950_in4,
        Din5 => VN1950_in5,
        VN2CN0_bit => VN_data_out(11700),
        VN2CN1_bit => VN_data_out(11701),
        VN2CN2_bit => VN_data_out(11702),
        VN2CN3_bit => VN_data_out(11703),
        VN2CN4_bit => VN_data_out(11704),
        VN2CN5_bit => VN_data_out(11705),
        VN2CN0_sign => VN_sign_out(11700),
        VN2CN1_sign => VN_sign_out(11701),
        VN2CN2_sign => VN_sign_out(11702),
        VN2CN3_sign => VN_sign_out(11703),
        VN2CN4_sign => VN_sign_out(11704),
        VN2CN5_sign => VN_sign_out(11705),
        codeword => codeword(1950),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1951 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11711 downto 11706),
        Din0 => VN1951_in0,
        Din1 => VN1951_in1,
        Din2 => VN1951_in2,
        Din3 => VN1951_in3,
        Din4 => VN1951_in4,
        Din5 => VN1951_in5,
        VN2CN0_bit => VN_data_out(11706),
        VN2CN1_bit => VN_data_out(11707),
        VN2CN2_bit => VN_data_out(11708),
        VN2CN3_bit => VN_data_out(11709),
        VN2CN4_bit => VN_data_out(11710),
        VN2CN5_bit => VN_data_out(11711),
        VN2CN0_sign => VN_sign_out(11706),
        VN2CN1_sign => VN_sign_out(11707),
        VN2CN2_sign => VN_sign_out(11708),
        VN2CN3_sign => VN_sign_out(11709),
        VN2CN4_sign => VN_sign_out(11710),
        VN2CN5_sign => VN_sign_out(11711),
        codeword => codeword(1951),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1952 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11717 downto 11712),
        Din0 => VN1952_in0,
        Din1 => VN1952_in1,
        Din2 => VN1952_in2,
        Din3 => VN1952_in3,
        Din4 => VN1952_in4,
        Din5 => VN1952_in5,
        VN2CN0_bit => VN_data_out(11712),
        VN2CN1_bit => VN_data_out(11713),
        VN2CN2_bit => VN_data_out(11714),
        VN2CN3_bit => VN_data_out(11715),
        VN2CN4_bit => VN_data_out(11716),
        VN2CN5_bit => VN_data_out(11717),
        VN2CN0_sign => VN_sign_out(11712),
        VN2CN1_sign => VN_sign_out(11713),
        VN2CN2_sign => VN_sign_out(11714),
        VN2CN3_sign => VN_sign_out(11715),
        VN2CN4_sign => VN_sign_out(11716),
        VN2CN5_sign => VN_sign_out(11717),
        codeword => codeword(1952),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1953 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11723 downto 11718),
        Din0 => VN1953_in0,
        Din1 => VN1953_in1,
        Din2 => VN1953_in2,
        Din3 => VN1953_in3,
        Din4 => VN1953_in4,
        Din5 => VN1953_in5,
        VN2CN0_bit => VN_data_out(11718),
        VN2CN1_bit => VN_data_out(11719),
        VN2CN2_bit => VN_data_out(11720),
        VN2CN3_bit => VN_data_out(11721),
        VN2CN4_bit => VN_data_out(11722),
        VN2CN5_bit => VN_data_out(11723),
        VN2CN0_sign => VN_sign_out(11718),
        VN2CN1_sign => VN_sign_out(11719),
        VN2CN2_sign => VN_sign_out(11720),
        VN2CN3_sign => VN_sign_out(11721),
        VN2CN4_sign => VN_sign_out(11722),
        VN2CN5_sign => VN_sign_out(11723),
        codeword => codeword(1953),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1954 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11729 downto 11724),
        Din0 => VN1954_in0,
        Din1 => VN1954_in1,
        Din2 => VN1954_in2,
        Din3 => VN1954_in3,
        Din4 => VN1954_in4,
        Din5 => VN1954_in5,
        VN2CN0_bit => VN_data_out(11724),
        VN2CN1_bit => VN_data_out(11725),
        VN2CN2_bit => VN_data_out(11726),
        VN2CN3_bit => VN_data_out(11727),
        VN2CN4_bit => VN_data_out(11728),
        VN2CN5_bit => VN_data_out(11729),
        VN2CN0_sign => VN_sign_out(11724),
        VN2CN1_sign => VN_sign_out(11725),
        VN2CN2_sign => VN_sign_out(11726),
        VN2CN3_sign => VN_sign_out(11727),
        VN2CN4_sign => VN_sign_out(11728),
        VN2CN5_sign => VN_sign_out(11729),
        codeword => codeword(1954),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1955 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11735 downto 11730),
        Din0 => VN1955_in0,
        Din1 => VN1955_in1,
        Din2 => VN1955_in2,
        Din3 => VN1955_in3,
        Din4 => VN1955_in4,
        Din5 => VN1955_in5,
        VN2CN0_bit => VN_data_out(11730),
        VN2CN1_bit => VN_data_out(11731),
        VN2CN2_bit => VN_data_out(11732),
        VN2CN3_bit => VN_data_out(11733),
        VN2CN4_bit => VN_data_out(11734),
        VN2CN5_bit => VN_data_out(11735),
        VN2CN0_sign => VN_sign_out(11730),
        VN2CN1_sign => VN_sign_out(11731),
        VN2CN2_sign => VN_sign_out(11732),
        VN2CN3_sign => VN_sign_out(11733),
        VN2CN4_sign => VN_sign_out(11734),
        VN2CN5_sign => VN_sign_out(11735),
        codeword => codeword(1955),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1956 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11741 downto 11736),
        Din0 => VN1956_in0,
        Din1 => VN1956_in1,
        Din2 => VN1956_in2,
        Din3 => VN1956_in3,
        Din4 => VN1956_in4,
        Din5 => VN1956_in5,
        VN2CN0_bit => VN_data_out(11736),
        VN2CN1_bit => VN_data_out(11737),
        VN2CN2_bit => VN_data_out(11738),
        VN2CN3_bit => VN_data_out(11739),
        VN2CN4_bit => VN_data_out(11740),
        VN2CN5_bit => VN_data_out(11741),
        VN2CN0_sign => VN_sign_out(11736),
        VN2CN1_sign => VN_sign_out(11737),
        VN2CN2_sign => VN_sign_out(11738),
        VN2CN3_sign => VN_sign_out(11739),
        VN2CN4_sign => VN_sign_out(11740),
        VN2CN5_sign => VN_sign_out(11741),
        codeword => codeword(1956),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1957 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11747 downto 11742),
        Din0 => VN1957_in0,
        Din1 => VN1957_in1,
        Din2 => VN1957_in2,
        Din3 => VN1957_in3,
        Din4 => VN1957_in4,
        Din5 => VN1957_in5,
        VN2CN0_bit => VN_data_out(11742),
        VN2CN1_bit => VN_data_out(11743),
        VN2CN2_bit => VN_data_out(11744),
        VN2CN3_bit => VN_data_out(11745),
        VN2CN4_bit => VN_data_out(11746),
        VN2CN5_bit => VN_data_out(11747),
        VN2CN0_sign => VN_sign_out(11742),
        VN2CN1_sign => VN_sign_out(11743),
        VN2CN2_sign => VN_sign_out(11744),
        VN2CN3_sign => VN_sign_out(11745),
        VN2CN4_sign => VN_sign_out(11746),
        VN2CN5_sign => VN_sign_out(11747),
        codeword => codeword(1957),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1958 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11753 downto 11748),
        Din0 => VN1958_in0,
        Din1 => VN1958_in1,
        Din2 => VN1958_in2,
        Din3 => VN1958_in3,
        Din4 => VN1958_in4,
        Din5 => VN1958_in5,
        VN2CN0_bit => VN_data_out(11748),
        VN2CN1_bit => VN_data_out(11749),
        VN2CN2_bit => VN_data_out(11750),
        VN2CN3_bit => VN_data_out(11751),
        VN2CN4_bit => VN_data_out(11752),
        VN2CN5_bit => VN_data_out(11753),
        VN2CN0_sign => VN_sign_out(11748),
        VN2CN1_sign => VN_sign_out(11749),
        VN2CN2_sign => VN_sign_out(11750),
        VN2CN3_sign => VN_sign_out(11751),
        VN2CN4_sign => VN_sign_out(11752),
        VN2CN5_sign => VN_sign_out(11753),
        codeword => codeword(1958),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1959 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11759 downto 11754),
        Din0 => VN1959_in0,
        Din1 => VN1959_in1,
        Din2 => VN1959_in2,
        Din3 => VN1959_in3,
        Din4 => VN1959_in4,
        Din5 => VN1959_in5,
        VN2CN0_bit => VN_data_out(11754),
        VN2CN1_bit => VN_data_out(11755),
        VN2CN2_bit => VN_data_out(11756),
        VN2CN3_bit => VN_data_out(11757),
        VN2CN4_bit => VN_data_out(11758),
        VN2CN5_bit => VN_data_out(11759),
        VN2CN0_sign => VN_sign_out(11754),
        VN2CN1_sign => VN_sign_out(11755),
        VN2CN2_sign => VN_sign_out(11756),
        VN2CN3_sign => VN_sign_out(11757),
        VN2CN4_sign => VN_sign_out(11758),
        VN2CN5_sign => VN_sign_out(11759),
        codeword => codeword(1959),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1960 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11765 downto 11760),
        Din0 => VN1960_in0,
        Din1 => VN1960_in1,
        Din2 => VN1960_in2,
        Din3 => VN1960_in3,
        Din4 => VN1960_in4,
        Din5 => VN1960_in5,
        VN2CN0_bit => VN_data_out(11760),
        VN2CN1_bit => VN_data_out(11761),
        VN2CN2_bit => VN_data_out(11762),
        VN2CN3_bit => VN_data_out(11763),
        VN2CN4_bit => VN_data_out(11764),
        VN2CN5_bit => VN_data_out(11765),
        VN2CN0_sign => VN_sign_out(11760),
        VN2CN1_sign => VN_sign_out(11761),
        VN2CN2_sign => VN_sign_out(11762),
        VN2CN3_sign => VN_sign_out(11763),
        VN2CN4_sign => VN_sign_out(11764),
        VN2CN5_sign => VN_sign_out(11765),
        codeword => codeword(1960),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1961 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11771 downto 11766),
        Din0 => VN1961_in0,
        Din1 => VN1961_in1,
        Din2 => VN1961_in2,
        Din3 => VN1961_in3,
        Din4 => VN1961_in4,
        Din5 => VN1961_in5,
        VN2CN0_bit => VN_data_out(11766),
        VN2CN1_bit => VN_data_out(11767),
        VN2CN2_bit => VN_data_out(11768),
        VN2CN3_bit => VN_data_out(11769),
        VN2CN4_bit => VN_data_out(11770),
        VN2CN5_bit => VN_data_out(11771),
        VN2CN0_sign => VN_sign_out(11766),
        VN2CN1_sign => VN_sign_out(11767),
        VN2CN2_sign => VN_sign_out(11768),
        VN2CN3_sign => VN_sign_out(11769),
        VN2CN4_sign => VN_sign_out(11770),
        VN2CN5_sign => VN_sign_out(11771),
        codeword => codeword(1961),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1962 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11777 downto 11772),
        Din0 => VN1962_in0,
        Din1 => VN1962_in1,
        Din2 => VN1962_in2,
        Din3 => VN1962_in3,
        Din4 => VN1962_in4,
        Din5 => VN1962_in5,
        VN2CN0_bit => VN_data_out(11772),
        VN2CN1_bit => VN_data_out(11773),
        VN2CN2_bit => VN_data_out(11774),
        VN2CN3_bit => VN_data_out(11775),
        VN2CN4_bit => VN_data_out(11776),
        VN2CN5_bit => VN_data_out(11777),
        VN2CN0_sign => VN_sign_out(11772),
        VN2CN1_sign => VN_sign_out(11773),
        VN2CN2_sign => VN_sign_out(11774),
        VN2CN3_sign => VN_sign_out(11775),
        VN2CN4_sign => VN_sign_out(11776),
        VN2CN5_sign => VN_sign_out(11777),
        codeword => codeword(1962),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1963 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11783 downto 11778),
        Din0 => VN1963_in0,
        Din1 => VN1963_in1,
        Din2 => VN1963_in2,
        Din3 => VN1963_in3,
        Din4 => VN1963_in4,
        Din5 => VN1963_in5,
        VN2CN0_bit => VN_data_out(11778),
        VN2CN1_bit => VN_data_out(11779),
        VN2CN2_bit => VN_data_out(11780),
        VN2CN3_bit => VN_data_out(11781),
        VN2CN4_bit => VN_data_out(11782),
        VN2CN5_bit => VN_data_out(11783),
        VN2CN0_sign => VN_sign_out(11778),
        VN2CN1_sign => VN_sign_out(11779),
        VN2CN2_sign => VN_sign_out(11780),
        VN2CN3_sign => VN_sign_out(11781),
        VN2CN4_sign => VN_sign_out(11782),
        VN2CN5_sign => VN_sign_out(11783),
        codeword => codeword(1963),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1964 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11789 downto 11784),
        Din0 => VN1964_in0,
        Din1 => VN1964_in1,
        Din2 => VN1964_in2,
        Din3 => VN1964_in3,
        Din4 => VN1964_in4,
        Din5 => VN1964_in5,
        VN2CN0_bit => VN_data_out(11784),
        VN2CN1_bit => VN_data_out(11785),
        VN2CN2_bit => VN_data_out(11786),
        VN2CN3_bit => VN_data_out(11787),
        VN2CN4_bit => VN_data_out(11788),
        VN2CN5_bit => VN_data_out(11789),
        VN2CN0_sign => VN_sign_out(11784),
        VN2CN1_sign => VN_sign_out(11785),
        VN2CN2_sign => VN_sign_out(11786),
        VN2CN3_sign => VN_sign_out(11787),
        VN2CN4_sign => VN_sign_out(11788),
        VN2CN5_sign => VN_sign_out(11789),
        codeword => codeword(1964),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1965 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11795 downto 11790),
        Din0 => VN1965_in0,
        Din1 => VN1965_in1,
        Din2 => VN1965_in2,
        Din3 => VN1965_in3,
        Din4 => VN1965_in4,
        Din5 => VN1965_in5,
        VN2CN0_bit => VN_data_out(11790),
        VN2CN1_bit => VN_data_out(11791),
        VN2CN2_bit => VN_data_out(11792),
        VN2CN3_bit => VN_data_out(11793),
        VN2CN4_bit => VN_data_out(11794),
        VN2CN5_bit => VN_data_out(11795),
        VN2CN0_sign => VN_sign_out(11790),
        VN2CN1_sign => VN_sign_out(11791),
        VN2CN2_sign => VN_sign_out(11792),
        VN2CN3_sign => VN_sign_out(11793),
        VN2CN4_sign => VN_sign_out(11794),
        VN2CN5_sign => VN_sign_out(11795),
        codeword => codeword(1965),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1966 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11801 downto 11796),
        Din0 => VN1966_in0,
        Din1 => VN1966_in1,
        Din2 => VN1966_in2,
        Din3 => VN1966_in3,
        Din4 => VN1966_in4,
        Din5 => VN1966_in5,
        VN2CN0_bit => VN_data_out(11796),
        VN2CN1_bit => VN_data_out(11797),
        VN2CN2_bit => VN_data_out(11798),
        VN2CN3_bit => VN_data_out(11799),
        VN2CN4_bit => VN_data_out(11800),
        VN2CN5_bit => VN_data_out(11801),
        VN2CN0_sign => VN_sign_out(11796),
        VN2CN1_sign => VN_sign_out(11797),
        VN2CN2_sign => VN_sign_out(11798),
        VN2CN3_sign => VN_sign_out(11799),
        VN2CN4_sign => VN_sign_out(11800),
        VN2CN5_sign => VN_sign_out(11801),
        codeword => codeword(1966),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1967 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11807 downto 11802),
        Din0 => VN1967_in0,
        Din1 => VN1967_in1,
        Din2 => VN1967_in2,
        Din3 => VN1967_in3,
        Din4 => VN1967_in4,
        Din5 => VN1967_in5,
        VN2CN0_bit => VN_data_out(11802),
        VN2CN1_bit => VN_data_out(11803),
        VN2CN2_bit => VN_data_out(11804),
        VN2CN3_bit => VN_data_out(11805),
        VN2CN4_bit => VN_data_out(11806),
        VN2CN5_bit => VN_data_out(11807),
        VN2CN0_sign => VN_sign_out(11802),
        VN2CN1_sign => VN_sign_out(11803),
        VN2CN2_sign => VN_sign_out(11804),
        VN2CN3_sign => VN_sign_out(11805),
        VN2CN4_sign => VN_sign_out(11806),
        VN2CN5_sign => VN_sign_out(11807),
        codeword => codeword(1967),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1968 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11813 downto 11808),
        Din0 => VN1968_in0,
        Din1 => VN1968_in1,
        Din2 => VN1968_in2,
        Din3 => VN1968_in3,
        Din4 => VN1968_in4,
        Din5 => VN1968_in5,
        VN2CN0_bit => VN_data_out(11808),
        VN2CN1_bit => VN_data_out(11809),
        VN2CN2_bit => VN_data_out(11810),
        VN2CN3_bit => VN_data_out(11811),
        VN2CN4_bit => VN_data_out(11812),
        VN2CN5_bit => VN_data_out(11813),
        VN2CN0_sign => VN_sign_out(11808),
        VN2CN1_sign => VN_sign_out(11809),
        VN2CN2_sign => VN_sign_out(11810),
        VN2CN3_sign => VN_sign_out(11811),
        VN2CN4_sign => VN_sign_out(11812),
        VN2CN5_sign => VN_sign_out(11813),
        codeword => codeword(1968),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1969 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11819 downto 11814),
        Din0 => VN1969_in0,
        Din1 => VN1969_in1,
        Din2 => VN1969_in2,
        Din3 => VN1969_in3,
        Din4 => VN1969_in4,
        Din5 => VN1969_in5,
        VN2CN0_bit => VN_data_out(11814),
        VN2CN1_bit => VN_data_out(11815),
        VN2CN2_bit => VN_data_out(11816),
        VN2CN3_bit => VN_data_out(11817),
        VN2CN4_bit => VN_data_out(11818),
        VN2CN5_bit => VN_data_out(11819),
        VN2CN0_sign => VN_sign_out(11814),
        VN2CN1_sign => VN_sign_out(11815),
        VN2CN2_sign => VN_sign_out(11816),
        VN2CN3_sign => VN_sign_out(11817),
        VN2CN4_sign => VN_sign_out(11818),
        VN2CN5_sign => VN_sign_out(11819),
        codeword => codeword(1969),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1970 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11825 downto 11820),
        Din0 => VN1970_in0,
        Din1 => VN1970_in1,
        Din2 => VN1970_in2,
        Din3 => VN1970_in3,
        Din4 => VN1970_in4,
        Din5 => VN1970_in5,
        VN2CN0_bit => VN_data_out(11820),
        VN2CN1_bit => VN_data_out(11821),
        VN2CN2_bit => VN_data_out(11822),
        VN2CN3_bit => VN_data_out(11823),
        VN2CN4_bit => VN_data_out(11824),
        VN2CN5_bit => VN_data_out(11825),
        VN2CN0_sign => VN_sign_out(11820),
        VN2CN1_sign => VN_sign_out(11821),
        VN2CN2_sign => VN_sign_out(11822),
        VN2CN3_sign => VN_sign_out(11823),
        VN2CN4_sign => VN_sign_out(11824),
        VN2CN5_sign => VN_sign_out(11825),
        codeword => codeword(1970),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1971 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11831 downto 11826),
        Din0 => VN1971_in0,
        Din1 => VN1971_in1,
        Din2 => VN1971_in2,
        Din3 => VN1971_in3,
        Din4 => VN1971_in4,
        Din5 => VN1971_in5,
        VN2CN0_bit => VN_data_out(11826),
        VN2CN1_bit => VN_data_out(11827),
        VN2CN2_bit => VN_data_out(11828),
        VN2CN3_bit => VN_data_out(11829),
        VN2CN4_bit => VN_data_out(11830),
        VN2CN5_bit => VN_data_out(11831),
        VN2CN0_sign => VN_sign_out(11826),
        VN2CN1_sign => VN_sign_out(11827),
        VN2CN2_sign => VN_sign_out(11828),
        VN2CN3_sign => VN_sign_out(11829),
        VN2CN4_sign => VN_sign_out(11830),
        VN2CN5_sign => VN_sign_out(11831),
        codeword => codeword(1971),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1972 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11837 downto 11832),
        Din0 => VN1972_in0,
        Din1 => VN1972_in1,
        Din2 => VN1972_in2,
        Din3 => VN1972_in3,
        Din4 => VN1972_in4,
        Din5 => VN1972_in5,
        VN2CN0_bit => VN_data_out(11832),
        VN2CN1_bit => VN_data_out(11833),
        VN2CN2_bit => VN_data_out(11834),
        VN2CN3_bit => VN_data_out(11835),
        VN2CN4_bit => VN_data_out(11836),
        VN2CN5_bit => VN_data_out(11837),
        VN2CN0_sign => VN_sign_out(11832),
        VN2CN1_sign => VN_sign_out(11833),
        VN2CN2_sign => VN_sign_out(11834),
        VN2CN3_sign => VN_sign_out(11835),
        VN2CN4_sign => VN_sign_out(11836),
        VN2CN5_sign => VN_sign_out(11837),
        codeword => codeword(1972),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1973 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11843 downto 11838),
        Din0 => VN1973_in0,
        Din1 => VN1973_in1,
        Din2 => VN1973_in2,
        Din3 => VN1973_in3,
        Din4 => VN1973_in4,
        Din5 => VN1973_in5,
        VN2CN0_bit => VN_data_out(11838),
        VN2CN1_bit => VN_data_out(11839),
        VN2CN2_bit => VN_data_out(11840),
        VN2CN3_bit => VN_data_out(11841),
        VN2CN4_bit => VN_data_out(11842),
        VN2CN5_bit => VN_data_out(11843),
        VN2CN0_sign => VN_sign_out(11838),
        VN2CN1_sign => VN_sign_out(11839),
        VN2CN2_sign => VN_sign_out(11840),
        VN2CN3_sign => VN_sign_out(11841),
        VN2CN4_sign => VN_sign_out(11842),
        VN2CN5_sign => VN_sign_out(11843),
        codeword => codeword(1973),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1974 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11849 downto 11844),
        Din0 => VN1974_in0,
        Din1 => VN1974_in1,
        Din2 => VN1974_in2,
        Din3 => VN1974_in3,
        Din4 => VN1974_in4,
        Din5 => VN1974_in5,
        VN2CN0_bit => VN_data_out(11844),
        VN2CN1_bit => VN_data_out(11845),
        VN2CN2_bit => VN_data_out(11846),
        VN2CN3_bit => VN_data_out(11847),
        VN2CN4_bit => VN_data_out(11848),
        VN2CN5_bit => VN_data_out(11849),
        VN2CN0_sign => VN_sign_out(11844),
        VN2CN1_sign => VN_sign_out(11845),
        VN2CN2_sign => VN_sign_out(11846),
        VN2CN3_sign => VN_sign_out(11847),
        VN2CN4_sign => VN_sign_out(11848),
        VN2CN5_sign => VN_sign_out(11849),
        codeword => codeword(1974),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1975 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11855 downto 11850),
        Din0 => VN1975_in0,
        Din1 => VN1975_in1,
        Din2 => VN1975_in2,
        Din3 => VN1975_in3,
        Din4 => VN1975_in4,
        Din5 => VN1975_in5,
        VN2CN0_bit => VN_data_out(11850),
        VN2CN1_bit => VN_data_out(11851),
        VN2CN2_bit => VN_data_out(11852),
        VN2CN3_bit => VN_data_out(11853),
        VN2CN4_bit => VN_data_out(11854),
        VN2CN5_bit => VN_data_out(11855),
        VN2CN0_sign => VN_sign_out(11850),
        VN2CN1_sign => VN_sign_out(11851),
        VN2CN2_sign => VN_sign_out(11852),
        VN2CN3_sign => VN_sign_out(11853),
        VN2CN4_sign => VN_sign_out(11854),
        VN2CN5_sign => VN_sign_out(11855),
        codeword => codeword(1975),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1976 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11861 downto 11856),
        Din0 => VN1976_in0,
        Din1 => VN1976_in1,
        Din2 => VN1976_in2,
        Din3 => VN1976_in3,
        Din4 => VN1976_in4,
        Din5 => VN1976_in5,
        VN2CN0_bit => VN_data_out(11856),
        VN2CN1_bit => VN_data_out(11857),
        VN2CN2_bit => VN_data_out(11858),
        VN2CN3_bit => VN_data_out(11859),
        VN2CN4_bit => VN_data_out(11860),
        VN2CN5_bit => VN_data_out(11861),
        VN2CN0_sign => VN_sign_out(11856),
        VN2CN1_sign => VN_sign_out(11857),
        VN2CN2_sign => VN_sign_out(11858),
        VN2CN3_sign => VN_sign_out(11859),
        VN2CN4_sign => VN_sign_out(11860),
        VN2CN5_sign => VN_sign_out(11861),
        codeword => codeword(1976),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1977 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11867 downto 11862),
        Din0 => VN1977_in0,
        Din1 => VN1977_in1,
        Din2 => VN1977_in2,
        Din3 => VN1977_in3,
        Din4 => VN1977_in4,
        Din5 => VN1977_in5,
        VN2CN0_bit => VN_data_out(11862),
        VN2CN1_bit => VN_data_out(11863),
        VN2CN2_bit => VN_data_out(11864),
        VN2CN3_bit => VN_data_out(11865),
        VN2CN4_bit => VN_data_out(11866),
        VN2CN5_bit => VN_data_out(11867),
        VN2CN0_sign => VN_sign_out(11862),
        VN2CN1_sign => VN_sign_out(11863),
        VN2CN2_sign => VN_sign_out(11864),
        VN2CN3_sign => VN_sign_out(11865),
        VN2CN4_sign => VN_sign_out(11866),
        VN2CN5_sign => VN_sign_out(11867),
        codeword => codeword(1977),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1978 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11873 downto 11868),
        Din0 => VN1978_in0,
        Din1 => VN1978_in1,
        Din2 => VN1978_in2,
        Din3 => VN1978_in3,
        Din4 => VN1978_in4,
        Din5 => VN1978_in5,
        VN2CN0_bit => VN_data_out(11868),
        VN2CN1_bit => VN_data_out(11869),
        VN2CN2_bit => VN_data_out(11870),
        VN2CN3_bit => VN_data_out(11871),
        VN2CN4_bit => VN_data_out(11872),
        VN2CN5_bit => VN_data_out(11873),
        VN2CN0_sign => VN_sign_out(11868),
        VN2CN1_sign => VN_sign_out(11869),
        VN2CN2_sign => VN_sign_out(11870),
        VN2CN3_sign => VN_sign_out(11871),
        VN2CN4_sign => VN_sign_out(11872),
        VN2CN5_sign => VN_sign_out(11873),
        codeword => codeword(1978),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1979 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11879 downto 11874),
        Din0 => VN1979_in0,
        Din1 => VN1979_in1,
        Din2 => VN1979_in2,
        Din3 => VN1979_in3,
        Din4 => VN1979_in4,
        Din5 => VN1979_in5,
        VN2CN0_bit => VN_data_out(11874),
        VN2CN1_bit => VN_data_out(11875),
        VN2CN2_bit => VN_data_out(11876),
        VN2CN3_bit => VN_data_out(11877),
        VN2CN4_bit => VN_data_out(11878),
        VN2CN5_bit => VN_data_out(11879),
        VN2CN0_sign => VN_sign_out(11874),
        VN2CN1_sign => VN_sign_out(11875),
        VN2CN2_sign => VN_sign_out(11876),
        VN2CN3_sign => VN_sign_out(11877),
        VN2CN4_sign => VN_sign_out(11878),
        VN2CN5_sign => VN_sign_out(11879),
        codeword => codeword(1979),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1980 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11885 downto 11880),
        Din0 => VN1980_in0,
        Din1 => VN1980_in1,
        Din2 => VN1980_in2,
        Din3 => VN1980_in3,
        Din4 => VN1980_in4,
        Din5 => VN1980_in5,
        VN2CN0_bit => VN_data_out(11880),
        VN2CN1_bit => VN_data_out(11881),
        VN2CN2_bit => VN_data_out(11882),
        VN2CN3_bit => VN_data_out(11883),
        VN2CN4_bit => VN_data_out(11884),
        VN2CN5_bit => VN_data_out(11885),
        VN2CN0_sign => VN_sign_out(11880),
        VN2CN1_sign => VN_sign_out(11881),
        VN2CN2_sign => VN_sign_out(11882),
        VN2CN3_sign => VN_sign_out(11883),
        VN2CN4_sign => VN_sign_out(11884),
        VN2CN5_sign => VN_sign_out(11885),
        codeword => codeword(1980),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1981 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11891 downto 11886),
        Din0 => VN1981_in0,
        Din1 => VN1981_in1,
        Din2 => VN1981_in2,
        Din3 => VN1981_in3,
        Din4 => VN1981_in4,
        Din5 => VN1981_in5,
        VN2CN0_bit => VN_data_out(11886),
        VN2CN1_bit => VN_data_out(11887),
        VN2CN2_bit => VN_data_out(11888),
        VN2CN3_bit => VN_data_out(11889),
        VN2CN4_bit => VN_data_out(11890),
        VN2CN5_bit => VN_data_out(11891),
        VN2CN0_sign => VN_sign_out(11886),
        VN2CN1_sign => VN_sign_out(11887),
        VN2CN2_sign => VN_sign_out(11888),
        VN2CN3_sign => VN_sign_out(11889),
        VN2CN4_sign => VN_sign_out(11890),
        VN2CN5_sign => VN_sign_out(11891),
        codeword => codeword(1981),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1982 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11897 downto 11892),
        Din0 => VN1982_in0,
        Din1 => VN1982_in1,
        Din2 => VN1982_in2,
        Din3 => VN1982_in3,
        Din4 => VN1982_in4,
        Din5 => VN1982_in5,
        VN2CN0_bit => VN_data_out(11892),
        VN2CN1_bit => VN_data_out(11893),
        VN2CN2_bit => VN_data_out(11894),
        VN2CN3_bit => VN_data_out(11895),
        VN2CN4_bit => VN_data_out(11896),
        VN2CN5_bit => VN_data_out(11897),
        VN2CN0_sign => VN_sign_out(11892),
        VN2CN1_sign => VN_sign_out(11893),
        VN2CN2_sign => VN_sign_out(11894),
        VN2CN3_sign => VN_sign_out(11895),
        VN2CN4_sign => VN_sign_out(11896),
        VN2CN5_sign => VN_sign_out(11897),
        codeword => codeword(1982),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1983 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11903 downto 11898),
        Din0 => VN1983_in0,
        Din1 => VN1983_in1,
        Din2 => VN1983_in2,
        Din3 => VN1983_in3,
        Din4 => VN1983_in4,
        Din5 => VN1983_in5,
        VN2CN0_bit => VN_data_out(11898),
        VN2CN1_bit => VN_data_out(11899),
        VN2CN2_bit => VN_data_out(11900),
        VN2CN3_bit => VN_data_out(11901),
        VN2CN4_bit => VN_data_out(11902),
        VN2CN5_bit => VN_data_out(11903),
        VN2CN0_sign => VN_sign_out(11898),
        VN2CN1_sign => VN_sign_out(11899),
        VN2CN2_sign => VN_sign_out(11900),
        VN2CN3_sign => VN_sign_out(11901),
        VN2CN4_sign => VN_sign_out(11902),
        VN2CN5_sign => VN_sign_out(11903),
        codeword => codeword(1983),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1984 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11909 downto 11904),
        Din0 => VN1984_in0,
        Din1 => VN1984_in1,
        Din2 => VN1984_in2,
        Din3 => VN1984_in3,
        Din4 => VN1984_in4,
        Din5 => VN1984_in5,
        VN2CN0_bit => VN_data_out(11904),
        VN2CN1_bit => VN_data_out(11905),
        VN2CN2_bit => VN_data_out(11906),
        VN2CN3_bit => VN_data_out(11907),
        VN2CN4_bit => VN_data_out(11908),
        VN2CN5_bit => VN_data_out(11909),
        VN2CN0_sign => VN_sign_out(11904),
        VN2CN1_sign => VN_sign_out(11905),
        VN2CN2_sign => VN_sign_out(11906),
        VN2CN3_sign => VN_sign_out(11907),
        VN2CN4_sign => VN_sign_out(11908),
        VN2CN5_sign => VN_sign_out(11909),
        codeword => codeword(1984),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1985 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11915 downto 11910),
        Din0 => VN1985_in0,
        Din1 => VN1985_in1,
        Din2 => VN1985_in2,
        Din3 => VN1985_in3,
        Din4 => VN1985_in4,
        Din5 => VN1985_in5,
        VN2CN0_bit => VN_data_out(11910),
        VN2CN1_bit => VN_data_out(11911),
        VN2CN2_bit => VN_data_out(11912),
        VN2CN3_bit => VN_data_out(11913),
        VN2CN4_bit => VN_data_out(11914),
        VN2CN5_bit => VN_data_out(11915),
        VN2CN0_sign => VN_sign_out(11910),
        VN2CN1_sign => VN_sign_out(11911),
        VN2CN2_sign => VN_sign_out(11912),
        VN2CN3_sign => VN_sign_out(11913),
        VN2CN4_sign => VN_sign_out(11914),
        VN2CN5_sign => VN_sign_out(11915),
        codeword => codeword(1985),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1986 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11921 downto 11916),
        Din0 => VN1986_in0,
        Din1 => VN1986_in1,
        Din2 => VN1986_in2,
        Din3 => VN1986_in3,
        Din4 => VN1986_in4,
        Din5 => VN1986_in5,
        VN2CN0_bit => VN_data_out(11916),
        VN2CN1_bit => VN_data_out(11917),
        VN2CN2_bit => VN_data_out(11918),
        VN2CN3_bit => VN_data_out(11919),
        VN2CN4_bit => VN_data_out(11920),
        VN2CN5_bit => VN_data_out(11921),
        VN2CN0_sign => VN_sign_out(11916),
        VN2CN1_sign => VN_sign_out(11917),
        VN2CN2_sign => VN_sign_out(11918),
        VN2CN3_sign => VN_sign_out(11919),
        VN2CN4_sign => VN_sign_out(11920),
        VN2CN5_sign => VN_sign_out(11921),
        codeword => codeword(1986),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1987 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11927 downto 11922),
        Din0 => VN1987_in0,
        Din1 => VN1987_in1,
        Din2 => VN1987_in2,
        Din3 => VN1987_in3,
        Din4 => VN1987_in4,
        Din5 => VN1987_in5,
        VN2CN0_bit => VN_data_out(11922),
        VN2CN1_bit => VN_data_out(11923),
        VN2CN2_bit => VN_data_out(11924),
        VN2CN3_bit => VN_data_out(11925),
        VN2CN4_bit => VN_data_out(11926),
        VN2CN5_bit => VN_data_out(11927),
        VN2CN0_sign => VN_sign_out(11922),
        VN2CN1_sign => VN_sign_out(11923),
        VN2CN2_sign => VN_sign_out(11924),
        VN2CN3_sign => VN_sign_out(11925),
        VN2CN4_sign => VN_sign_out(11926),
        VN2CN5_sign => VN_sign_out(11927),
        codeword => codeword(1987),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1988 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11933 downto 11928),
        Din0 => VN1988_in0,
        Din1 => VN1988_in1,
        Din2 => VN1988_in2,
        Din3 => VN1988_in3,
        Din4 => VN1988_in4,
        Din5 => VN1988_in5,
        VN2CN0_bit => VN_data_out(11928),
        VN2CN1_bit => VN_data_out(11929),
        VN2CN2_bit => VN_data_out(11930),
        VN2CN3_bit => VN_data_out(11931),
        VN2CN4_bit => VN_data_out(11932),
        VN2CN5_bit => VN_data_out(11933),
        VN2CN0_sign => VN_sign_out(11928),
        VN2CN1_sign => VN_sign_out(11929),
        VN2CN2_sign => VN_sign_out(11930),
        VN2CN3_sign => VN_sign_out(11931),
        VN2CN4_sign => VN_sign_out(11932),
        VN2CN5_sign => VN_sign_out(11933),
        codeword => codeword(1988),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1989 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11939 downto 11934),
        Din0 => VN1989_in0,
        Din1 => VN1989_in1,
        Din2 => VN1989_in2,
        Din3 => VN1989_in3,
        Din4 => VN1989_in4,
        Din5 => VN1989_in5,
        VN2CN0_bit => VN_data_out(11934),
        VN2CN1_bit => VN_data_out(11935),
        VN2CN2_bit => VN_data_out(11936),
        VN2CN3_bit => VN_data_out(11937),
        VN2CN4_bit => VN_data_out(11938),
        VN2CN5_bit => VN_data_out(11939),
        VN2CN0_sign => VN_sign_out(11934),
        VN2CN1_sign => VN_sign_out(11935),
        VN2CN2_sign => VN_sign_out(11936),
        VN2CN3_sign => VN_sign_out(11937),
        VN2CN4_sign => VN_sign_out(11938),
        VN2CN5_sign => VN_sign_out(11939),
        codeword => codeword(1989),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1990 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11945 downto 11940),
        Din0 => VN1990_in0,
        Din1 => VN1990_in1,
        Din2 => VN1990_in2,
        Din3 => VN1990_in3,
        Din4 => VN1990_in4,
        Din5 => VN1990_in5,
        VN2CN0_bit => VN_data_out(11940),
        VN2CN1_bit => VN_data_out(11941),
        VN2CN2_bit => VN_data_out(11942),
        VN2CN3_bit => VN_data_out(11943),
        VN2CN4_bit => VN_data_out(11944),
        VN2CN5_bit => VN_data_out(11945),
        VN2CN0_sign => VN_sign_out(11940),
        VN2CN1_sign => VN_sign_out(11941),
        VN2CN2_sign => VN_sign_out(11942),
        VN2CN3_sign => VN_sign_out(11943),
        VN2CN4_sign => VN_sign_out(11944),
        VN2CN5_sign => VN_sign_out(11945),
        codeword => codeword(1990),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1991 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11951 downto 11946),
        Din0 => VN1991_in0,
        Din1 => VN1991_in1,
        Din2 => VN1991_in2,
        Din3 => VN1991_in3,
        Din4 => VN1991_in4,
        Din5 => VN1991_in5,
        VN2CN0_bit => VN_data_out(11946),
        VN2CN1_bit => VN_data_out(11947),
        VN2CN2_bit => VN_data_out(11948),
        VN2CN3_bit => VN_data_out(11949),
        VN2CN4_bit => VN_data_out(11950),
        VN2CN5_bit => VN_data_out(11951),
        VN2CN0_sign => VN_sign_out(11946),
        VN2CN1_sign => VN_sign_out(11947),
        VN2CN2_sign => VN_sign_out(11948),
        VN2CN3_sign => VN_sign_out(11949),
        VN2CN4_sign => VN_sign_out(11950),
        VN2CN5_sign => VN_sign_out(11951),
        codeword => codeword(1991),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1992 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11957 downto 11952),
        Din0 => VN1992_in0,
        Din1 => VN1992_in1,
        Din2 => VN1992_in2,
        Din3 => VN1992_in3,
        Din4 => VN1992_in4,
        Din5 => VN1992_in5,
        VN2CN0_bit => VN_data_out(11952),
        VN2CN1_bit => VN_data_out(11953),
        VN2CN2_bit => VN_data_out(11954),
        VN2CN3_bit => VN_data_out(11955),
        VN2CN4_bit => VN_data_out(11956),
        VN2CN5_bit => VN_data_out(11957),
        VN2CN0_sign => VN_sign_out(11952),
        VN2CN1_sign => VN_sign_out(11953),
        VN2CN2_sign => VN_sign_out(11954),
        VN2CN3_sign => VN_sign_out(11955),
        VN2CN4_sign => VN_sign_out(11956),
        VN2CN5_sign => VN_sign_out(11957),
        codeword => codeword(1992),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1993 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11963 downto 11958),
        Din0 => VN1993_in0,
        Din1 => VN1993_in1,
        Din2 => VN1993_in2,
        Din3 => VN1993_in3,
        Din4 => VN1993_in4,
        Din5 => VN1993_in5,
        VN2CN0_bit => VN_data_out(11958),
        VN2CN1_bit => VN_data_out(11959),
        VN2CN2_bit => VN_data_out(11960),
        VN2CN3_bit => VN_data_out(11961),
        VN2CN4_bit => VN_data_out(11962),
        VN2CN5_bit => VN_data_out(11963),
        VN2CN0_sign => VN_sign_out(11958),
        VN2CN1_sign => VN_sign_out(11959),
        VN2CN2_sign => VN_sign_out(11960),
        VN2CN3_sign => VN_sign_out(11961),
        VN2CN4_sign => VN_sign_out(11962),
        VN2CN5_sign => VN_sign_out(11963),
        codeword => codeword(1993),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1994 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11969 downto 11964),
        Din0 => VN1994_in0,
        Din1 => VN1994_in1,
        Din2 => VN1994_in2,
        Din3 => VN1994_in3,
        Din4 => VN1994_in4,
        Din5 => VN1994_in5,
        VN2CN0_bit => VN_data_out(11964),
        VN2CN1_bit => VN_data_out(11965),
        VN2CN2_bit => VN_data_out(11966),
        VN2CN3_bit => VN_data_out(11967),
        VN2CN4_bit => VN_data_out(11968),
        VN2CN5_bit => VN_data_out(11969),
        VN2CN0_sign => VN_sign_out(11964),
        VN2CN1_sign => VN_sign_out(11965),
        VN2CN2_sign => VN_sign_out(11966),
        VN2CN3_sign => VN_sign_out(11967),
        VN2CN4_sign => VN_sign_out(11968),
        VN2CN5_sign => VN_sign_out(11969),
        codeword => codeword(1994),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1995 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11975 downto 11970),
        Din0 => VN1995_in0,
        Din1 => VN1995_in1,
        Din2 => VN1995_in2,
        Din3 => VN1995_in3,
        Din4 => VN1995_in4,
        Din5 => VN1995_in5,
        VN2CN0_bit => VN_data_out(11970),
        VN2CN1_bit => VN_data_out(11971),
        VN2CN2_bit => VN_data_out(11972),
        VN2CN3_bit => VN_data_out(11973),
        VN2CN4_bit => VN_data_out(11974),
        VN2CN5_bit => VN_data_out(11975),
        VN2CN0_sign => VN_sign_out(11970),
        VN2CN1_sign => VN_sign_out(11971),
        VN2CN2_sign => VN_sign_out(11972),
        VN2CN3_sign => VN_sign_out(11973),
        VN2CN4_sign => VN_sign_out(11974),
        VN2CN5_sign => VN_sign_out(11975),
        codeword => codeword(1995),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1996 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11981 downto 11976),
        Din0 => VN1996_in0,
        Din1 => VN1996_in1,
        Din2 => VN1996_in2,
        Din3 => VN1996_in3,
        Din4 => VN1996_in4,
        Din5 => VN1996_in5,
        VN2CN0_bit => VN_data_out(11976),
        VN2CN1_bit => VN_data_out(11977),
        VN2CN2_bit => VN_data_out(11978),
        VN2CN3_bit => VN_data_out(11979),
        VN2CN4_bit => VN_data_out(11980),
        VN2CN5_bit => VN_data_out(11981),
        VN2CN0_sign => VN_sign_out(11976),
        VN2CN1_sign => VN_sign_out(11977),
        VN2CN2_sign => VN_sign_out(11978),
        VN2CN3_sign => VN_sign_out(11979),
        VN2CN4_sign => VN_sign_out(11980),
        VN2CN5_sign => VN_sign_out(11981),
        codeword => codeword(1996),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1997 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11987 downto 11982),
        Din0 => VN1997_in0,
        Din1 => VN1997_in1,
        Din2 => VN1997_in2,
        Din3 => VN1997_in3,
        Din4 => VN1997_in4,
        Din5 => VN1997_in5,
        VN2CN0_bit => VN_data_out(11982),
        VN2CN1_bit => VN_data_out(11983),
        VN2CN2_bit => VN_data_out(11984),
        VN2CN3_bit => VN_data_out(11985),
        VN2CN4_bit => VN_data_out(11986),
        VN2CN5_bit => VN_data_out(11987),
        VN2CN0_sign => VN_sign_out(11982),
        VN2CN1_sign => VN_sign_out(11983),
        VN2CN2_sign => VN_sign_out(11984),
        VN2CN3_sign => VN_sign_out(11985),
        VN2CN4_sign => VN_sign_out(11986),
        VN2CN5_sign => VN_sign_out(11987),
        codeword => codeword(1997),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1998 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11993 downto 11988),
        Din0 => VN1998_in0,
        Din1 => VN1998_in1,
        Din2 => VN1998_in2,
        Din3 => VN1998_in3,
        Din4 => VN1998_in4,
        Din5 => VN1998_in5,
        VN2CN0_bit => VN_data_out(11988),
        VN2CN1_bit => VN_data_out(11989),
        VN2CN2_bit => VN_data_out(11990),
        VN2CN3_bit => VN_data_out(11991),
        VN2CN4_bit => VN_data_out(11992),
        VN2CN5_bit => VN_data_out(11993),
        VN2CN0_sign => VN_sign_out(11988),
        VN2CN1_sign => VN_sign_out(11989),
        VN2CN2_sign => VN_sign_out(11990),
        VN2CN3_sign => VN_sign_out(11991),
        VN2CN4_sign => VN_sign_out(11992),
        VN2CN5_sign => VN_sign_out(11993),
        codeword => codeword(1998),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN1999 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(11999 downto 11994),
        Din0 => VN1999_in0,
        Din1 => VN1999_in1,
        Din2 => VN1999_in2,
        Din3 => VN1999_in3,
        Din4 => VN1999_in4,
        Din5 => VN1999_in5,
        VN2CN0_bit => VN_data_out(11994),
        VN2CN1_bit => VN_data_out(11995),
        VN2CN2_bit => VN_data_out(11996),
        VN2CN3_bit => VN_data_out(11997),
        VN2CN4_bit => VN_data_out(11998),
        VN2CN5_bit => VN_data_out(11999),
        VN2CN0_sign => VN_sign_out(11994),
        VN2CN1_sign => VN_sign_out(11995),
        VN2CN2_sign => VN_sign_out(11996),
        VN2CN3_sign => VN_sign_out(11997),
        VN2CN4_sign => VN_sign_out(11998),
        VN2CN5_sign => VN_sign_out(11999),
        codeword => codeword(1999),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2000 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12005 downto 12000),
        Din0 => VN2000_in0,
        Din1 => VN2000_in1,
        Din2 => VN2000_in2,
        Din3 => VN2000_in3,
        Din4 => VN2000_in4,
        Din5 => VN2000_in5,
        VN2CN0_bit => VN_data_out(12000),
        VN2CN1_bit => VN_data_out(12001),
        VN2CN2_bit => VN_data_out(12002),
        VN2CN3_bit => VN_data_out(12003),
        VN2CN4_bit => VN_data_out(12004),
        VN2CN5_bit => VN_data_out(12005),
        VN2CN0_sign => VN_sign_out(12000),
        VN2CN1_sign => VN_sign_out(12001),
        VN2CN2_sign => VN_sign_out(12002),
        VN2CN3_sign => VN_sign_out(12003),
        VN2CN4_sign => VN_sign_out(12004),
        VN2CN5_sign => VN_sign_out(12005),
        codeword => codeword(2000),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2001 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12011 downto 12006),
        Din0 => VN2001_in0,
        Din1 => VN2001_in1,
        Din2 => VN2001_in2,
        Din3 => VN2001_in3,
        Din4 => VN2001_in4,
        Din5 => VN2001_in5,
        VN2CN0_bit => VN_data_out(12006),
        VN2CN1_bit => VN_data_out(12007),
        VN2CN2_bit => VN_data_out(12008),
        VN2CN3_bit => VN_data_out(12009),
        VN2CN4_bit => VN_data_out(12010),
        VN2CN5_bit => VN_data_out(12011),
        VN2CN0_sign => VN_sign_out(12006),
        VN2CN1_sign => VN_sign_out(12007),
        VN2CN2_sign => VN_sign_out(12008),
        VN2CN3_sign => VN_sign_out(12009),
        VN2CN4_sign => VN_sign_out(12010),
        VN2CN5_sign => VN_sign_out(12011),
        codeword => codeword(2001),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2002 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12017 downto 12012),
        Din0 => VN2002_in0,
        Din1 => VN2002_in1,
        Din2 => VN2002_in2,
        Din3 => VN2002_in3,
        Din4 => VN2002_in4,
        Din5 => VN2002_in5,
        VN2CN0_bit => VN_data_out(12012),
        VN2CN1_bit => VN_data_out(12013),
        VN2CN2_bit => VN_data_out(12014),
        VN2CN3_bit => VN_data_out(12015),
        VN2CN4_bit => VN_data_out(12016),
        VN2CN5_bit => VN_data_out(12017),
        VN2CN0_sign => VN_sign_out(12012),
        VN2CN1_sign => VN_sign_out(12013),
        VN2CN2_sign => VN_sign_out(12014),
        VN2CN3_sign => VN_sign_out(12015),
        VN2CN4_sign => VN_sign_out(12016),
        VN2CN5_sign => VN_sign_out(12017),
        codeword => codeword(2002),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2003 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12023 downto 12018),
        Din0 => VN2003_in0,
        Din1 => VN2003_in1,
        Din2 => VN2003_in2,
        Din3 => VN2003_in3,
        Din4 => VN2003_in4,
        Din5 => VN2003_in5,
        VN2CN0_bit => VN_data_out(12018),
        VN2CN1_bit => VN_data_out(12019),
        VN2CN2_bit => VN_data_out(12020),
        VN2CN3_bit => VN_data_out(12021),
        VN2CN4_bit => VN_data_out(12022),
        VN2CN5_bit => VN_data_out(12023),
        VN2CN0_sign => VN_sign_out(12018),
        VN2CN1_sign => VN_sign_out(12019),
        VN2CN2_sign => VN_sign_out(12020),
        VN2CN3_sign => VN_sign_out(12021),
        VN2CN4_sign => VN_sign_out(12022),
        VN2CN5_sign => VN_sign_out(12023),
        codeword => codeword(2003),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2004 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12029 downto 12024),
        Din0 => VN2004_in0,
        Din1 => VN2004_in1,
        Din2 => VN2004_in2,
        Din3 => VN2004_in3,
        Din4 => VN2004_in4,
        Din5 => VN2004_in5,
        VN2CN0_bit => VN_data_out(12024),
        VN2CN1_bit => VN_data_out(12025),
        VN2CN2_bit => VN_data_out(12026),
        VN2CN3_bit => VN_data_out(12027),
        VN2CN4_bit => VN_data_out(12028),
        VN2CN5_bit => VN_data_out(12029),
        VN2CN0_sign => VN_sign_out(12024),
        VN2CN1_sign => VN_sign_out(12025),
        VN2CN2_sign => VN_sign_out(12026),
        VN2CN3_sign => VN_sign_out(12027),
        VN2CN4_sign => VN_sign_out(12028),
        VN2CN5_sign => VN_sign_out(12029),
        codeword => codeword(2004),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2005 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12035 downto 12030),
        Din0 => VN2005_in0,
        Din1 => VN2005_in1,
        Din2 => VN2005_in2,
        Din3 => VN2005_in3,
        Din4 => VN2005_in4,
        Din5 => VN2005_in5,
        VN2CN0_bit => VN_data_out(12030),
        VN2CN1_bit => VN_data_out(12031),
        VN2CN2_bit => VN_data_out(12032),
        VN2CN3_bit => VN_data_out(12033),
        VN2CN4_bit => VN_data_out(12034),
        VN2CN5_bit => VN_data_out(12035),
        VN2CN0_sign => VN_sign_out(12030),
        VN2CN1_sign => VN_sign_out(12031),
        VN2CN2_sign => VN_sign_out(12032),
        VN2CN3_sign => VN_sign_out(12033),
        VN2CN4_sign => VN_sign_out(12034),
        VN2CN5_sign => VN_sign_out(12035),
        codeword => codeword(2005),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2006 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12041 downto 12036),
        Din0 => VN2006_in0,
        Din1 => VN2006_in1,
        Din2 => VN2006_in2,
        Din3 => VN2006_in3,
        Din4 => VN2006_in4,
        Din5 => VN2006_in5,
        VN2CN0_bit => VN_data_out(12036),
        VN2CN1_bit => VN_data_out(12037),
        VN2CN2_bit => VN_data_out(12038),
        VN2CN3_bit => VN_data_out(12039),
        VN2CN4_bit => VN_data_out(12040),
        VN2CN5_bit => VN_data_out(12041),
        VN2CN0_sign => VN_sign_out(12036),
        VN2CN1_sign => VN_sign_out(12037),
        VN2CN2_sign => VN_sign_out(12038),
        VN2CN3_sign => VN_sign_out(12039),
        VN2CN4_sign => VN_sign_out(12040),
        VN2CN5_sign => VN_sign_out(12041),
        codeword => codeword(2006),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2007 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12047 downto 12042),
        Din0 => VN2007_in0,
        Din1 => VN2007_in1,
        Din2 => VN2007_in2,
        Din3 => VN2007_in3,
        Din4 => VN2007_in4,
        Din5 => VN2007_in5,
        VN2CN0_bit => VN_data_out(12042),
        VN2CN1_bit => VN_data_out(12043),
        VN2CN2_bit => VN_data_out(12044),
        VN2CN3_bit => VN_data_out(12045),
        VN2CN4_bit => VN_data_out(12046),
        VN2CN5_bit => VN_data_out(12047),
        VN2CN0_sign => VN_sign_out(12042),
        VN2CN1_sign => VN_sign_out(12043),
        VN2CN2_sign => VN_sign_out(12044),
        VN2CN3_sign => VN_sign_out(12045),
        VN2CN4_sign => VN_sign_out(12046),
        VN2CN5_sign => VN_sign_out(12047),
        codeword => codeword(2007),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2008 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12053 downto 12048),
        Din0 => VN2008_in0,
        Din1 => VN2008_in1,
        Din2 => VN2008_in2,
        Din3 => VN2008_in3,
        Din4 => VN2008_in4,
        Din5 => VN2008_in5,
        VN2CN0_bit => VN_data_out(12048),
        VN2CN1_bit => VN_data_out(12049),
        VN2CN2_bit => VN_data_out(12050),
        VN2CN3_bit => VN_data_out(12051),
        VN2CN4_bit => VN_data_out(12052),
        VN2CN5_bit => VN_data_out(12053),
        VN2CN0_sign => VN_sign_out(12048),
        VN2CN1_sign => VN_sign_out(12049),
        VN2CN2_sign => VN_sign_out(12050),
        VN2CN3_sign => VN_sign_out(12051),
        VN2CN4_sign => VN_sign_out(12052),
        VN2CN5_sign => VN_sign_out(12053),
        codeword => codeword(2008),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2009 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12059 downto 12054),
        Din0 => VN2009_in0,
        Din1 => VN2009_in1,
        Din2 => VN2009_in2,
        Din3 => VN2009_in3,
        Din4 => VN2009_in4,
        Din5 => VN2009_in5,
        VN2CN0_bit => VN_data_out(12054),
        VN2CN1_bit => VN_data_out(12055),
        VN2CN2_bit => VN_data_out(12056),
        VN2CN3_bit => VN_data_out(12057),
        VN2CN4_bit => VN_data_out(12058),
        VN2CN5_bit => VN_data_out(12059),
        VN2CN0_sign => VN_sign_out(12054),
        VN2CN1_sign => VN_sign_out(12055),
        VN2CN2_sign => VN_sign_out(12056),
        VN2CN3_sign => VN_sign_out(12057),
        VN2CN4_sign => VN_sign_out(12058),
        VN2CN5_sign => VN_sign_out(12059),
        codeword => codeword(2009),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2010 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12065 downto 12060),
        Din0 => VN2010_in0,
        Din1 => VN2010_in1,
        Din2 => VN2010_in2,
        Din3 => VN2010_in3,
        Din4 => VN2010_in4,
        Din5 => VN2010_in5,
        VN2CN0_bit => VN_data_out(12060),
        VN2CN1_bit => VN_data_out(12061),
        VN2CN2_bit => VN_data_out(12062),
        VN2CN3_bit => VN_data_out(12063),
        VN2CN4_bit => VN_data_out(12064),
        VN2CN5_bit => VN_data_out(12065),
        VN2CN0_sign => VN_sign_out(12060),
        VN2CN1_sign => VN_sign_out(12061),
        VN2CN2_sign => VN_sign_out(12062),
        VN2CN3_sign => VN_sign_out(12063),
        VN2CN4_sign => VN_sign_out(12064),
        VN2CN5_sign => VN_sign_out(12065),
        codeword => codeword(2010),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2011 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12071 downto 12066),
        Din0 => VN2011_in0,
        Din1 => VN2011_in1,
        Din2 => VN2011_in2,
        Din3 => VN2011_in3,
        Din4 => VN2011_in4,
        Din5 => VN2011_in5,
        VN2CN0_bit => VN_data_out(12066),
        VN2CN1_bit => VN_data_out(12067),
        VN2CN2_bit => VN_data_out(12068),
        VN2CN3_bit => VN_data_out(12069),
        VN2CN4_bit => VN_data_out(12070),
        VN2CN5_bit => VN_data_out(12071),
        VN2CN0_sign => VN_sign_out(12066),
        VN2CN1_sign => VN_sign_out(12067),
        VN2CN2_sign => VN_sign_out(12068),
        VN2CN3_sign => VN_sign_out(12069),
        VN2CN4_sign => VN_sign_out(12070),
        VN2CN5_sign => VN_sign_out(12071),
        codeword => codeword(2011),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2012 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12077 downto 12072),
        Din0 => VN2012_in0,
        Din1 => VN2012_in1,
        Din2 => VN2012_in2,
        Din3 => VN2012_in3,
        Din4 => VN2012_in4,
        Din5 => VN2012_in5,
        VN2CN0_bit => VN_data_out(12072),
        VN2CN1_bit => VN_data_out(12073),
        VN2CN2_bit => VN_data_out(12074),
        VN2CN3_bit => VN_data_out(12075),
        VN2CN4_bit => VN_data_out(12076),
        VN2CN5_bit => VN_data_out(12077),
        VN2CN0_sign => VN_sign_out(12072),
        VN2CN1_sign => VN_sign_out(12073),
        VN2CN2_sign => VN_sign_out(12074),
        VN2CN3_sign => VN_sign_out(12075),
        VN2CN4_sign => VN_sign_out(12076),
        VN2CN5_sign => VN_sign_out(12077),
        codeword => codeword(2012),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2013 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12083 downto 12078),
        Din0 => VN2013_in0,
        Din1 => VN2013_in1,
        Din2 => VN2013_in2,
        Din3 => VN2013_in3,
        Din4 => VN2013_in4,
        Din5 => VN2013_in5,
        VN2CN0_bit => VN_data_out(12078),
        VN2CN1_bit => VN_data_out(12079),
        VN2CN2_bit => VN_data_out(12080),
        VN2CN3_bit => VN_data_out(12081),
        VN2CN4_bit => VN_data_out(12082),
        VN2CN5_bit => VN_data_out(12083),
        VN2CN0_sign => VN_sign_out(12078),
        VN2CN1_sign => VN_sign_out(12079),
        VN2CN2_sign => VN_sign_out(12080),
        VN2CN3_sign => VN_sign_out(12081),
        VN2CN4_sign => VN_sign_out(12082),
        VN2CN5_sign => VN_sign_out(12083),
        codeword => codeword(2013),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2014 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12089 downto 12084),
        Din0 => VN2014_in0,
        Din1 => VN2014_in1,
        Din2 => VN2014_in2,
        Din3 => VN2014_in3,
        Din4 => VN2014_in4,
        Din5 => VN2014_in5,
        VN2CN0_bit => VN_data_out(12084),
        VN2CN1_bit => VN_data_out(12085),
        VN2CN2_bit => VN_data_out(12086),
        VN2CN3_bit => VN_data_out(12087),
        VN2CN4_bit => VN_data_out(12088),
        VN2CN5_bit => VN_data_out(12089),
        VN2CN0_sign => VN_sign_out(12084),
        VN2CN1_sign => VN_sign_out(12085),
        VN2CN2_sign => VN_sign_out(12086),
        VN2CN3_sign => VN_sign_out(12087),
        VN2CN4_sign => VN_sign_out(12088),
        VN2CN5_sign => VN_sign_out(12089),
        codeword => codeword(2014),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2015 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12095 downto 12090),
        Din0 => VN2015_in0,
        Din1 => VN2015_in1,
        Din2 => VN2015_in2,
        Din3 => VN2015_in3,
        Din4 => VN2015_in4,
        Din5 => VN2015_in5,
        VN2CN0_bit => VN_data_out(12090),
        VN2CN1_bit => VN_data_out(12091),
        VN2CN2_bit => VN_data_out(12092),
        VN2CN3_bit => VN_data_out(12093),
        VN2CN4_bit => VN_data_out(12094),
        VN2CN5_bit => VN_data_out(12095),
        VN2CN0_sign => VN_sign_out(12090),
        VN2CN1_sign => VN_sign_out(12091),
        VN2CN2_sign => VN_sign_out(12092),
        VN2CN3_sign => VN_sign_out(12093),
        VN2CN4_sign => VN_sign_out(12094),
        VN2CN5_sign => VN_sign_out(12095),
        codeword => codeword(2015),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2016 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12101 downto 12096),
        Din0 => VN2016_in0,
        Din1 => VN2016_in1,
        Din2 => VN2016_in2,
        Din3 => VN2016_in3,
        Din4 => VN2016_in4,
        Din5 => VN2016_in5,
        VN2CN0_bit => VN_data_out(12096),
        VN2CN1_bit => VN_data_out(12097),
        VN2CN2_bit => VN_data_out(12098),
        VN2CN3_bit => VN_data_out(12099),
        VN2CN4_bit => VN_data_out(12100),
        VN2CN5_bit => VN_data_out(12101),
        VN2CN0_sign => VN_sign_out(12096),
        VN2CN1_sign => VN_sign_out(12097),
        VN2CN2_sign => VN_sign_out(12098),
        VN2CN3_sign => VN_sign_out(12099),
        VN2CN4_sign => VN_sign_out(12100),
        VN2CN5_sign => VN_sign_out(12101),
        codeword => codeword(2016),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2017 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12107 downto 12102),
        Din0 => VN2017_in0,
        Din1 => VN2017_in1,
        Din2 => VN2017_in2,
        Din3 => VN2017_in3,
        Din4 => VN2017_in4,
        Din5 => VN2017_in5,
        VN2CN0_bit => VN_data_out(12102),
        VN2CN1_bit => VN_data_out(12103),
        VN2CN2_bit => VN_data_out(12104),
        VN2CN3_bit => VN_data_out(12105),
        VN2CN4_bit => VN_data_out(12106),
        VN2CN5_bit => VN_data_out(12107),
        VN2CN0_sign => VN_sign_out(12102),
        VN2CN1_sign => VN_sign_out(12103),
        VN2CN2_sign => VN_sign_out(12104),
        VN2CN3_sign => VN_sign_out(12105),
        VN2CN4_sign => VN_sign_out(12106),
        VN2CN5_sign => VN_sign_out(12107),
        codeword => codeword(2017),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2018 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12113 downto 12108),
        Din0 => VN2018_in0,
        Din1 => VN2018_in1,
        Din2 => VN2018_in2,
        Din3 => VN2018_in3,
        Din4 => VN2018_in4,
        Din5 => VN2018_in5,
        VN2CN0_bit => VN_data_out(12108),
        VN2CN1_bit => VN_data_out(12109),
        VN2CN2_bit => VN_data_out(12110),
        VN2CN3_bit => VN_data_out(12111),
        VN2CN4_bit => VN_data_out(12112),
        VN2CN5_bit => VN_data_out(12113),
        VN2CN0_sign => VN_sign_out(12108),
        VN2CN1_sign => VN_sign_out(12109),
        VN2CN2_sign => VN_sign_out(12110),
        VN2CN3_sign => VN_sign_out(12111),
        VN2CN4_sign => VN_sign_out(12112),
        VN2CN5_sign => VN_sign_out(12113),
        codeword => codeword(2018),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2019 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12119 downto 12114),
        Din0 => VN2019_in0,
        Din1 => VN2019_in1,
        Din2 => VN2019_in2,
        Din3 => VN2019_in3,
        Din4 => VN2019_in4,
        Din5 => VN2019_in5,
        VN2CN0_bit => VN_data_out(12114),
        VN2CN1_bit => VN_data_out(12115),
        VN2CN2_bit => VN_data_out(12116),
        VN2CN3_bit => VN_data_out(12117),
        VN2CN4_bit => VN_data_out(12118),
        VN2CN5_bit => VN_data_out(12119),
        VN2CN0_sign => VN_sign_out(12114),
        VN2CN1_sign => VN_sign_out(12115),
        VN2CN2_sign => VN_sign_out(12116),
        VN2CN3_sign => VN_sign_out(12117),
        VN2CN4_sign => VN_sign_out(12118),
        VN2CN5_sign => VN_sign_out(12119),
        codeword => codeword(2019),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2020 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12125 downto 12120),
        Din0 => VN2020_in0,
        Din1 => VN2020_in1,
        Din2 => VN2020_in2,
        Din3 => VN2020_in3,
        Din4 => VN2020_in4,
        Din5 => VN2020_in5,
        VN2CN0_bit => VN_data_out(12120),
        VN2CN1_bit => VN_data_out(12121),
        VN2CN2_bit => VN_data_out(12122),
        VN2CN3_bit => VN_data_out(12123),
        VN2CN4_bit => VN_data_out(12124),
        VN2CN5_bit => VN_data_out(12125),
        VN2CN0_sign => VN_sign_out(12120),
        VN2CN1_sign => VN_sign_out(12121),
        VN2CN2_sign => VN_sign_out(12122),
        VN2CN3_sign => VN_sign_out(12123),
        VN2CN4_sign => VN_sign_out(12124),
        VN2CN5_sign => VN_sign_out(12125),
        codeword => codeword(2020),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2021 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12131 downto 12126),
        Din0 => VN2021_in0,
        Din1 => VN2021_in1,
        Din2 => VN2021_in2,
        Din3 => VN2021_in3,
        Din4 => VN2021_in4,
        Din5 => VN2021_in5,
        VN2CN0_bit => VN_data_out(12126),
        VN2CN1_bit => VN_data_out(12127),
        VN2CN2_bit => VN_data_out(12128),
        VN2CN3_bit => VN_data_out(12129),
        VN2CN4_bit => VN_data_out(12130),
        VN2CN5_bit => VN_data_out(12131),
        VN2CN0_sign => VN_sign_out(12126),
        VN2CN1_sign => VN_sign_out(12127),
        VN2CN2_sign => VN_sign_out(12128),
        VN2CN3_sign => VN_sign_out(12129),
        VN2CN4_sign => VN_sign_out(12130),
        VN2CN5_sign => VN_sign_out(12131),
        codeword => codeword(2021),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2022 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12137 downto 12132),
        Din0 => VN2022_in0,
        Din1 => VN2022_in1,
        Din2 => VN2022_in2,
        Din3 => VN2022_in3,
        Din4 => VN2022_in4,
        Din5 => VN2022_in5,
        VN2CN0_bit => VN_data_out(12132),
        VN2CN1_bit => VN_data_out(12133),
        VN2CN2_bit => VN_data_out(12134),
        VN2CN3_bit => VN_data_out(12135),
        VN2CN4_bit => VN_data_out(12136),
        VN2CN5_bit => VN_data_out(12137),
        VN2CN0_sign => VN_sign_out(12132),
        VN2CN1_sign => VN_sign_out(12133),
        VN2CN2_sign => VN_sign_out(12134),
        VN2CN3_sign => VN_sign_out(12135),
        VN2CN4_sign => VN_sign_out(12136),
        VN2CN5_sign => VN_sign_out(12137),
        codeword => codeword(2022),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2023 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12143 downto 12138),
        Din0 => VN2023_in0,
        Din1 => VN2023_in1,
        Din2 => VN2023_in2,
        Din3 => VN2023_in3,
        Din4 => VN2023_in4,
        Din5 => VN2023_in5,
        VN2CN0_bit => VN_data_out(12138),
        VN2CN1_bit => VN_data_out(12139),
        VN2CN2_bit => VN_data_out(12140),
        VN2CN3_bit => VN_data_out(12141),
        VN2CN4_bit => VN_data_out(12142),
        VN2CN5_bit => VN_data_out(12143),
        VN2CN0_sign => VN_sign_out(12138),
        VN2CN1_sign => VN_sign_out(12139),
        VN2CN2_sign => VN_sign_out(12140),
        VN2CN3_sign => VN_sign_out(12141),
        VN2CN4_sign => VN_sign_out(12142),
        VN2CN5_sign => VN_sign_out(12143),
        codeword => codeword(2023),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2024 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12149 downto 12144),
        Din0 => VN2024_in0,
        Din1 => VN2024_in1,
        Din2 => VN2024_in2,
        Din3 => VN2024_in3,
        Din4 => VN2024_in4,
        Din5 => VN2024_in5,
        VN2CN0_bit => VN_data_out(12144),
        VN2CN1_bit => VN_data_out(12145),
        VN2CN2_bit => VN_data_out(12146),
        VN2CN3_bit => VN_data_out(12147),
        VN2CN4_bit => VN_data_out(12148),
        VN2CN5_bit => VN_data_out(12149),
        VN2CN0_sign => VN_sign_out(12144),
        VN2CN1_sign => VN_sign_out(12145),
        VN2CN2_sign => VN_sign_out(12146),
        VN2CN3_sign => VN_sign_out(12147),
        VN2CN4_sign => VN_sign_out(12148),
        VN2CN5_sign => VN_sign_out(12149),
        codeword => codeword(2024),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2025 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12155 downto 12150),
        Din0 => VN2025_in0,
        Din1 => VN2025_in1,
        Din2 => VN2025_in2,
        Din3 => VN2025_in3,
        Din4 => VN2025_in4,
        Din5 => VN2025_in5,
        VN2CN0_bit => VN_data_out(12150),
        VN2CN1_bit => VN_data_out(12151),
        VN2CN2_bit => VN_data_out(12152),
        VN2CN3_bit => VN_data_out(12153),
        VN2CN4_bit => VN_data_out(12154),
        VN2CN5_bit => VN_data_out(12155),
        VN2CN0_sign => VN_sign_out(12150),
        VN2CN1_sign => VN_sign_out(12151),
        VN2CN2_sign => VN_sign_out(12152),
        VN2CN3_sign => VN_sign_out(12153),
        VN2CN4_sign => VN_sign_out(12154),
        VN2CN5_sign => VN_sign_out(12155),
        codeword => codeword(2025),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2026 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12161 downto 12156),
        Din0 => VN2026_in0,
        Din1 => VN2026_in1,
        Din2 => VN2026_in2,
        Din3 => VN2026_in3,
        Din4 => VN2026_in4,
        Din5 => VN2026_in5,
        VN2CN0_bit => VN_data_out(12156),
        VN2CN1_bit => VN_data_out(12157),
        VN2CN2_bit => VN_data_out(12158),
        VN2CN3_bit => VN_data_out(12159),
        VN2CN4_bit => VN_data_out(12160),
        VN2CN5_bit => VN_data_out(12161),
        VN2CN0_sign => VN_sign_out(12156),
        VN2CN1_sign => VN_sign_out(12157),
        VN2CN2_sign => VN_sign_out(12158),
        VN2CN3_sign => VN_sign_out(12159),
        VN2CN4_sign => VN_sign_out(12160),
        VN2CN5_sign => VN_sign_out(12161),
        codeword => codeword(2026),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2027 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12167 downto 12162),
        Din0 => VN2027_in0,
        Din1 => VN2027_in1,
        Din2 => VN2027_in2,
        Din3 => VN2027_in3,
        Din4 => VN2027_in4,
        Din5 => VN2027_in5,
        VN2CN0_bit => VN_data_out(12162),
        VN2CN1_bit => VN_data_out(12163),
        VN2CN2_bit => VN_data_out(12164),
        VN2CN3_bit => VN_data_out(12165),
        VN2CN4_bit => VN_data_out(12166),
        VN2CN5_bit => VN_data_out(12167),
        VN2CN0_sign => VN_sign_out(12162),
        VN2CN1_sign => VN_sign_out(12163),
        VN2CN2_sign => VN_sign_out(12164),
        VN2CN3_sign => VN_sign_out(12165),
        VN2CN4_sign => VN_sign_out(12166),
        VN2CN5_sign => VN_sign_out(12167),
        codeword => codeword(2027),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2028 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12173 downto 12168),
        Din0 => VN2028_in0,
        Din1 => VN2028_in1,
        Din2 => VN2028_in2,
        Din3 => VN2028_in3,
        Din4 => VN2028_in4,
        Din5 => VN2028_in5,
        VN2CN0_bit => VN_data_out(12168),
        VN2CN1_bit => VN_data_out(12169),
        VN2CN2_bit => VN_data_out(12170),
        VN2CN3_bit => VN_data_out(12171),
        VN2CN4_bit => VN_data_out(12172),
        VN2CN5_bit => VN_data_out(12173),
        VN2CN0_sign => VN_sign_out(12168),
        VN2CN1_sign => VN_sign_out(12169),
        VN2CN2_sign => VN_sign_out(12170),
        VN2CN3_sign => VN_sign_out(12171),
        VN2CN4_sign => VN_sign_out(12172),
        VN2CN5_sign => VN_sign_out(12173),
        codeword => codeword(2028),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2029 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12179 downto 12174),
        Din0 => VN2029_in0,
        Din1 => VN2029_in1,
        Din2 => VN2029_in2,
        Din3 => VN2029_in3,
        Din4 => VN2029_in4,
        Din5 => VN2029_in5,
        VN2CN0_bit => VN_data_out(12174),
        VN2CN1_bit => VN_data_out(12175),
        VN2CN2_bit => VN_data_out(12176),
        VN2CN3_bit => VN_data_out(12177),
        VN2CN4_bit => VN_data_out(12178),
        VN2CN5_bit => VN_data_out(12179),
        VN2CN0_sign => VN_sign_out(12174),
        VN2CN1_sign => VN_sign_out(12175),
        VN2CN2_sign => VN_sign_out(12176),
        VN2CN3_sign => VN_sign_out(12177),
        VN2CN4_sign => VN_sign_out(12178),
        VN2CN5_sign => VN_sign_out(12179),
        codeword => codeword(2029),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2030 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12185 downto 12180),
        Din0 => VN2030_in0,
        Din1 => VN2030_in1,
        Din2 => VN2030_in2,
        Din3 => VN2030_in3,
        Din4 => VN2030_in4,
        Din5 => VN2030_in5,
        VN2CN0_bit => VN_data_out(12180),
        VN2CN1_bit => VN_data_out(12181),
        VN2CN2_bit => VN_data_out(12182),
        VN2CN3_bit => VN_data_out(12183),
        VN2CN4_bit => VN_data_out(12184),
        VN2CN5_bit => VN_data_out(12185),
        VN2CN0_sign => VN_sign_out(12180),
        VN2CN1_sign => VN_sign_out(12181),
        VN2CN2_sign => VN_sign_out(12182),
        VN2CN3_sign => VN_sign_out(12183),
        VN2CN4_sign => VN_sign_out(12184),
        VN2CN5_sign => VN_sign_out(12185),
        codeword => codeword(2030),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2031 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12191 downto 12186),
        Din0 => VN2031_in0,
        Din1 => VN2031_in1,
        Din2 => VN2031_in2,
        Din3 => VN2031_in3,
        Din4 => VN2031_in4,
        Din5 => VN2031_in5,
        VN2CN0_bit => VN_data_out(12186),
        VN2CN1_bit => VN_data_out(12187),
        VN2CN2_bit => VN_data_out(12188),
        VN2CN3_bit => VN_data_out(12189),
        VN2CN4_bit => VN_data_out(12190),
        VN2CN5_bit => VN_data_out(12191),
        VN2CN0_sign => VN_sign_out(12186),
        VN2CN1_sign => VN_sign_out(12187),
        VN2CN2_sign => VN_sign_out(12188),
        VN2CN3_sign => VN_sign_out(12189),
        VN2CN4_sign => VN_sign_out(12190),
        VN2CN5_sign => VN_sign_out(12191),
        codeword => codeword(2031),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2032 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12197 downto 12192),
        Din0 => VN2032_in0,
        Din1 => VN2032_in1,
        Din2 => VN2032_in2,
        Din3 => VN2032_in3,
        Din4 => VN2032_in4,
        Din5 => VN2032_in5,
        VN2CN0_bit => VN_data_out(12192),
        VN2CN1_bit => VN_data_out(12193),
        VN2CN2_bit => VN_data_out(12194),
        VN2CN3_bit => VN_data_out(12195),
        VN2CN4_bit => VN_data_out(12196),
        VN2CN5_bit => VN_data_out(12197),
        VN2CN0_sign => VN_sign_out(12192),
        VN2CN1_sign => VN_sign_out(12193),
        VN2CN2_sign => VN_sign_out(12194),
        VN2CN3_sign => VN_sign_out(12195),
        VN2CN4_sign => VN_sign_out(12196),
        VN2CN5_sign => VN_sign_out(12197),
        codeword => codeword(2032),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2033 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12203 downto 12198),
        Din0 => VN2033_in0,
        Din1 => VN2033_in1,
        Din2 => VN2033_in2,
        Din3 => VN2033_in3,
        Din4 => VN2033_in4,
        Din5 => VN2033_in5,
        VN2CN0_bit => VN_data_out(12198),
        VN2CN1_bit => VN_data_out(12199),
        VN2CN2_bit => VN_data_out(12200),
        VN2CN3_bit => VN_data_out(12201),
        VN2CN4_bit => VN_data_out(12202),
        VN2CN5_bit => VN_data_out(12203),
        VN2CN0_sign => VN_sign_out(12198),
        VN2CN1_sign => VN_sign_out(12199),
        VN2CN2_sign => VN_sign_out(12200),
        VN2CN3_sign => VN_sign_out(12201),
        VN2CN4_sign => VN_sign_out(12202),
        VN2CN5_sign => VN_sign_out(12203),
        codeword => codeword(2033),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2034 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12209 downto 12204),
        Din0 => VN2034_in0,
        Din1 => VN2034_in1,
        Din2 => VN2034_in2,
        Din3 => VN2034_in3,
        Din4 => VN2034_in4,
        Din5 => VN2034_in5,
        VN2CN0_bit => VN_data_out(12204),
        VN2CN1_bit => VN_data_out(12205),
        VN2CN2_bit => VN_data_out(12206),
        VN2CN3_bit => VN_data_out(12207),
        VN2CN4_bit => VN_data_out(12208),
        VN2CN5_bit => VN_data_out(12209),
        VN2CN0_sign => VN_sign_out(12204),
        VN2CN1_sign => VN_sign_out(12205),
        VN2CN2_sign => VN_sign_out(12206),
        VN2CN3_sign => VN_sign_out(12207),
        VN2CN4_sign => VN_sign_out(12208),
        VN2CN5_sign => VN_sign_out(12209),
        codeword => codeword(2034),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2035 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12215 downto 12210),
        Din0 => VN2035_in0,
        Din1 => VN2035_in1,
        Din2 => VN2035_in2,
        Din3 => VN2035_in3,
        Din4 => VN2035_in4,
        Din5 => VN2035_in5,
        VN2CN0_bit => VN_data_out(12210),
        VN2CN1_bit => VN_data_out(12211),
        VN2CN2_bit => VN_data_out(12212),
        VN2CN3_bit => VN_data_out(12213),
        VN2CN4_bit => VN_data_out(12214),
        VN2CN5_bit => VN_data_out(12215),
        VN2CN0_sign => VN_sign_out(12210),
        VN2CN1_sign => VN_sign_out(12211),
        VN2CN2_sign => VN_sign_out(12212),
        VN2CN3_sign => VN_sign_out(12213),
        VN2CN4_sign => VN_sign_out(12214),
        VN2CN5_sign => VN_sign_out(12215),
        codeword => codeword(2035),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2036 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12221 downto 12216),
        Din0 => VN2036_in0,
        Din1 => VN2036_in1,
        Din2 => VN2036_in2,
        Din3 => VN2036_in3,
        Din4 => VN2036_in4,
        Din5 => VN2036_in5,
        VN2CN0_bit => VN_data_out(12216),
        VN2CN1_bit => VN_data_out(12217),
        VN2CN2_bit => VN_data_out(12218),
        VN2CN3_bit => VN_data_out(12219),
        VN2CN4_bit => VN_data_out(12220),
        VN2CN5_bit => VN_data_out(12221),
        VN2CN0_sign => VN_sign_out(12216),
        VN2CN1_sign => VN_sign_out(12217),
        VN2CN2_sign => VN_sign_out(12218),
        VN2CN3_sign => VN_sign_out(12219),
        VN2CN4_sign => VN_sign_out(12220),
        VN2CN5_sign => VN_sign_out(12221),
        codeword => codeword(2036),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2037 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12227 downto 12222),
        Din0 => VN2037_in0,
        Din1 => VN2037_in1,
        Din2 => VN2037_in2,
        Din3 => VN2037_in3,
        Din4 => VN2037_in4,
        Din5 => VN2037_in5,
        VN2CN0_bit => VN_data_out(12222),
        VN2CN1_bit => VN_data_out(12223),
        VN2CN2_bit => VN_data_out(12224),
        VN2CN3_bit => VN_data_out(12225),
        VN2CN4_bit => VN_data_out(12226),
        VN2CN5_bit => VN_data_out(12227),
        VN2CN0_sign => VN_sign_out(12222),
        VN2CN1_sign => VN_sign_out(12223),
        VN2CN2_sign => VN_sign_out(12224),
        VN2CN3_sign => VN_sign_out(12225),
        VN2CN4_sign => VN_sign_out(12226),
        VN2CN5_sign => VN_sign_out(12227),
        codeword => codeword(2037),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2038 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12233 downto 12228),
        Din0 => VN2038_in0,
        Din1 => VN2038_in1,
        Din2 => VN2038_in2,
        Din3 => VN2038_in3,
        Din4 => VN2038_in4,
        Din5 => VN2038_in5,
        VN2CN0_bit => VN_data_out(12228),
        VN2CN1_bit => VN_data_out(12229),
        VN2CN2_bit => VN_data_out(12230),
        VN2CN3_bit => VN_data_out(12231),
        VN2CN4_bit => VN_data_out(12232),
        VN2CN5_bit => VN_data_out(12233),
        VN2CN0_sign => VN_sign_out(12228),
        VN2CN1_sign => VN_sign_out(12229),
        VN2CN2_sign => VN_sign_out(12230),
        VN2CN3_sign => VN_sign_out(12231),
        VN2CN4_sign => VN_sign_out(12232),
        VN2CN5_sign => VN_sign_out(12233),
        codeword => codeword(2038),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2039 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12239 downto 12234),
        Din0 => VN2039_in0,
        Din1 => VN2039_in1,
        Din2 => VN2039_in2,
        Din3 => VN2039_in3,
        Din4 => VN2039_in4,
        Din5 => VN2039_in5,
        VN2CN0_bit => VN_data_out(12234),
        VN2CN1_bit => VN_data_out(12235),
        VN2CN2_bit => VN_data_out(12236),
        VN2CN3_bit => VN_data_out(12237),
        VN2CN4_bit => VN_data_out(12238),
        VN2CN5_bit => VN_data_out(12239),
        VN2CN0_sign => VN_sign_out(12234),
        VN2CN1_sign => VN_sign_out(12235),
        VN2CN2_sign => VN_sign_out(12236),
        VN2CN3_sign => VN_sign_out(12237),
        VN2CN4_sign => VN_sign_out(12238),
        VN2CN5_sign => VN_sign_out(12239),
        codeword => codeword(2039),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2040 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12245 downto 12240),
        Din0 => VN2040_in0,
        Din1 => VN2040_in1,
        Din2 => VN2040_in2,
        Din3 => VN2040_in3,
        Din4 => VN2040_in4,
        Din5 => VN2040_in5,
        VN2CN0_bit => VN_data_out(12240),
        VN2CN1_bit => VN_data_out(12241),
        VN2CN2_bit => VN_data_out(12242),
        VN2CN3_bit => VN_data_out(12243),
        VN2CN4_bit => VN_data_out(12244),
        VN2CN5_bit => VN_data_out(12245),
        VN2CN0_sign => VN_sign_out(12240),
        VN2CN1_sign => VN_sign_out(12241),
        VN2CN2_sign => VN_sign_out(12242),
        VN2CN3_sign => VN_sign_out(12243),
        VN2CN4_sign => VN_sign_out(12244),
        VN2CN5_sign => VN_sign_out(12245),
        codeword => codeword(2040),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2041 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12251 downto 12246),
        Din0 => VN2041_in0,
        Din1 => VN2041_in1,
        Din2 => VN2041_in2,
        Din3 => VN2041_in3,
        Din4 => VN2041_in4,
        Din5 => VN2041_in5,
        VN2CN0_bit => VN_data_out(12246),
        VN2CN1_bit => VN_data_out(12247),
        VN2CN2_bit => VN_data_out(12248),
        VN2CN3_bit => VN_data_out(12249),
        VN2CN4_bit => VN_data_out(12250),
        VN2CN5_bit => VN_data_out(12251),
        VN2CN0_sign => VN_sign_out(12246),
        VN2CN1_sign => VN_sign_out(12247),
        VN2CN2_sign => VN_sign_out(12248),
        VN2CN3_sign => VN_sign_out(12249),
        VN2CN4_sign => VN_sign_out(12250),
        VN2CN5_sign => VN_sign_out(12251),
        codeword => codeword(2041),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2042 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12257 downto 12252),
        Din0 => VN2042_in0,
        Din1 => VN2042_in1,
        Din2 => VN2042_in2,
        Din3 => VN2042_in3,
        Din4 => VN2042_in4,
        Din5 => VN2042_in5,
        VN2CN0_bit => VN_data_out(12252),
        VN2CN1_bit => VN_data_out(12253),
        VN2CN2_bit => VN_data_out(12254),
        VN2CN3_bit => VN_data_out(12255),
        VN2CN4_bit => VN_data_out(12256),
        VN2CN5_bit => VN_data_out(12257),
        VN2CN0_sign => VN_sign_out(12252),
        VN2CN1_sign => VN_sign_out(12253),
        VN2CN2_sign => VN_sign_out(12254),
        VN2CN3_sign => VN_sign_out(12255),
        VN2CN4_sign => VN_sign_out(12256),
        VN2CN5_sign => VN_sign_out(12257),
        codeword => codeword(2042),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2043 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12263 downto 12258),
        Din0 => VN2043_in0,
        Din1 => VN2043_in1,
        Din2 => VN2043_in2,
        Din3 => VN2043_in3,
        Din4 => VN2043_in4,
        Din5 => VN2043_in5,
        VN2CN0_bit => VN_data_out(12258),
        VN2CN1_bit => VN_data_out(12259),
        VN2CN2_bit => VN_data_out(12260),
        VN2CN3_bit => VN_data_out(12261),
        VN2CN4_bit => VN_data_out(12262),
        VN2CN5_bit => VN_data_out(12263),
        VN2CN0_sign => VN_sign_out(12258),
        VN2CN1_sign => VN_sign_out(12259),
        VN2CN2_sign => VN_sign_out(12260),
        VN2CN3_sign => VN_sign_out(12261),
        VN2CN4_sign => VN_sign_out(12262),
        VN2CN5_sign => VN_sign_out(12263),
        codeword => codeword(2043),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2044 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12269 downto 12264),
        Din0 => VN2044_in0,
        Din1 => VN2044_in1,
        Din2 => VN2044_in2,
        Din3 => VN2044_in3,
        Din4 => VN2044_in4,
        Din5 => VN2044_in5,
        VN2CN0_bit => VN_data_out(12264),
        VN2CN1_bit => VN_data_out(12265),
        VN2CN2_bit => VN_data_out(12266),
        VN2CN3_bit => VN_data_out(12267),
        VN2CN4_bit => VN_data_out(12268),
        VN2CN5_bit => VN_data_out(12269),
        VN2CN0_sign => VN_sign_out(12264),
        VN2CN1_sign => VN_sign_out(12265),
        VN2CN2_sign => VN_sign_out(12266),
        VN2CN3_sign => VN_sign_out(12267),
        VN2CN4_sign => VN_sign_out(12268),
        VN2CN5_sign => VN_sign_out(12269),
        codeword => codeword(2044),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2045 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12275 downto 12270),
        Din0 => VN2045_in0,
        Din1 => VN2045_in1,
        Din2 => VN2045_in2,
        Din3 => VN2045_in3,
        Din4 => VN2045_in4,
        Din5 => VN2045_in5,
        VN2CN0_bit => VN_data_out(12270),
        VN2CN1_bit => VN_data_out(12271),
        VN2CN2_bit => VN_data_out(12272),
        VN2CN3_bit => VN_data_out(12273),
        VN2CN4_bit => VN_data_out(12274),
        VN2CN5_bit => VN_data_out(12275),
        VN2CN0_sign => VN_sign_out(12270),
        VN2CN1_sign => VN_sign_out(12271),
        VN2CN2_sign => VN_sign_out(12272),
        VN2CN3_sign => VN_sign_out(12273),
        VN2CN4_sign => VN_sign_out(12274),
        VN2CN5_sign => VN_sign_out(12275),
        codeword => codeword(2045),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2046 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12281 downto 12276),
        Din0 => VN2046_in0,
        Din1 => VN2046_in1,
        Din2 => VN2046_in2,
        Din3 => VN2046_in3,
        Din4 => VN2046_in4,
        Din5 => VN2046_in5,
        VN2CN0_bit => VN_data_out(12276),
        VN2CN1_bit => VN_data_out(12277),
        VN2CN2_bit => VN_data_out(12278),
        VN2CN3_bit => VN_data_out(12279),
        VN2CN4_bit => VN_data_out(12280),
        VN2CN5_bit => VN_data_out(12281),
        VN2CN0_sign => VN_sign_out(12276),
        VN2CN1_sign => VN_sign_out(12277),
        VN2CN2_sign => VN_sign_out(12278),
        VN2CN3_sign => VN_sign_out(12279),
        VN2CN4_sign => VN_sign_out(12280),
        VN2CN5_sign => VN_sign_out(12281),
        codeword => codeword(2046),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );
    VN2047 : VN_Dv6 port map(
        clk =>clk,
        rst_n => rst_n,
        New_LLR => New_LLR,
        DecoderOver => DecoderOver,
        RandomNum => RandomNum,
        LLR => LLR(12287 downto 12282),
        Din0 => VN2047_in0,
        Din1 => VN2047_in1,
        Din2 => VN2047_in2,
        Din3 => VN2047_in3,
        Din4 => VN2047_in4,
        Din5 => VN2047_in5,
        VN2CN0_bit => VN_data_out(12282),
        VN2CN1_bit => VN_data_out(12283),
        VN2CN2_bit => VN_data_out(12284),
        VN2CN3_bit => VN_data_out(12285),
        VN2CN4_bit => VN_data_out(12286),
        VN2CN5_bit => VN_data_out(12287),
        VN2CN0_sign => VN_sign_out(12282),
        VN2CN1_sign => VN_sign_out(12283),
        VN2CN2_sign => VN_sign_out(12284),
        VN2CN3_sign => VN_sign_out(12285),
        VN2CN4_sign => VN_sign_out(12286),
        VN2CN5_sign => VN_sign_out(12287),
        codeword => codeword(2047),
        Iterations => open,
        DV_out => open,
        DecodeState => open
    );

end architecture; --arch  

